// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bx+9j49KajS4xJK1DcBIKk/IoMpJehgb5H04UVoj0/50TdQ59FICT/7OG189AwCz
J31RBpRiHnfShdZgxOhmNFTIBm2SCekxIKY/h1/YlTi9c90p29YEo+v8ZWb+BaPn
6Oc8i1+J4ztARSkTKu/0bFDj2tVQsr7CUH+V74AEPGA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3344)
rABlU3qNIcsZhICAX+Lyxnx6jHxZnduPfiNCue/l+7GdFEA70JPFJyPGRhNWF46M
91BwL1aLguBKlc9iBRs+J0IDcV6geetMIMSNPHa6QEFooanHZSJs4bRDAm85C9U6
JCPAy2wp9vogXxiWyN2Bnst+d176M8xtFzTrXiou1KevUdfjujwXBG/ILgDW7RNu
8vUpTF98AHzHwiLALqpeijEVUbsPkPy8xV7ka8s9AbEzQklTXJdYu5tkb8u06zwQ
V1AW0tkVzlln+PvNZyBXFcocNdW6rt6xJ96UR/Lvt3gFID+FThTQsOwnMbrM3U3w
hVkFZ63oij+0tu9AiOOTX+B5w/J+xQvYg9RVHNxqDqzMCqVUav6oTpa0+TpmseQr
fNrUe0yTjL+PztBZ4Gdy8KTH7HT8YqspkxdffxzNe2Uk1rOGjC9outxaoIuonJ5f
H9tnWGiJL3jtdTBL9vpMCSSU64hU1ry6oAqEoV0qcioY+/xR5yGkVmITut7IFs07
h1PSbMIk/+yQ+uxZmDfnyjhiDNI775o3CtOxydVe+CKWEazh/Tu/fT7xye38akDY
TosMyDFQ+YsEJBm3R9ISyd3BrflEDaH0NLc/lg+q+7YvtjtGLJIJjNt51ltJHIIu
5guSqDP0nfqwQd2fTABAilfdQjPrFbx6zkuOhXmBzzBp2ZS44l1qkWbqj2hBC29p
EZ89ggxKclr6ugoXMz3YRGnxK95sywrXhLTcyqsPA4z3jSE7/tuXz3k9WcxpHHVr
qI/jJ6/QXXSl3nQylYiE/IsK5uvvcJKj4/I58eFHAagLs5iMbz23nWpEKObX6B3Q
dWcgrzR207hh1q5L85QEPNfIfRAvD4Sd8nbp2bGr/X0+HJc6LqpzP6dlW27YPxRW
S7TGF/1xdfNC3O5sqN8KQwqGpUvom7/ijaOuySYLHG2vX67xWLfEYXw/hdLU57xe
9OWDCvB+65if15ehd5zD1T4kmNs8yX4ZQ4itrbv7YSyqJdvYrS3Bd9rER0Wj5V2X
YggRjnkTn1VsWDKth0wDd0mJRUymrtB4uCdz7q/Wkcg7K3o9+ppkSVpWEFlGO3mG
j3wUOEVzH1uZ293n0GrMJJNHjydWfQU11j3v1G5gmF9vbwgWAPtzsqzgT2CSapbG
RN0j3v376+sl3pEcE7poHoAZgnF640/IHJ10yGhreHcT0jb63LLDoIof9dm7H55V
ieGJ24pduA07aXlQXWJm5iudiCgmsZSVjqbdfqO93OxxOhhw0J1CAEk9k4tgoeoD
KlEFBdJqHGrGEMfFtejrtFNNE7zqwgMRkpEZ23DaDa+beqr+Lgf9c/8tyOkKi6A/
t8Fn79f+XWmxTKC/tKy8oHpFJnlGd/sUKj7ubJsIFk1Wnl4YrSAnn5ujNmM4DVuV
8/pStNOgy1m9sGzy9JFts2E9WwKcqiJS0WiehuiI1Zw/QSeQgGc6jG7HKfGE0pFI
IoFkK/WjuJ1lAxR5p9oUKLC+1ReAk9T1Q7Wj3C6fDOCHdcrIwcSh6JzT+ZB0J4/1
MLhxOl/bIAWm0bwCJb0SMG5IrAXUE5+T82ZQf45pzMAzxRZ69xJ7++VyJp2VhBho
OpftcEk5fQ+L4ib5LXDl40oBnpYlP+kltdFVIDbrygS8WTLPSt/t/HnvEtcYI+UN
e2NirQe3rXrBJeglkO3cjT+0QrUWHCNpOVAmo1Zj80hy0sFU3KB7Wtf44+/YQ3JJ
mY9AhGhYmsmzgRDI2k/zQY55XRPAkJFX4Xuh9tr966NymVoWavZE8nV8L5l/ubJq
KdiRJYspD2aGNZ9DNwkY8ZWR3Mx574KshQJItUyg2fcJqEFEnCrBSkY7kkOprPfW
zNjTHqv49Ukdt3KQGVj6F0QeVtPMVPNb6Pj7TzIgwmawo/MLBNw6b1IB5Pa5Ms+A
yjPGrxKFR2A+vgTWruCxnV63Ux+nBy+7V0US3UUsh+abOCv2091a1HBgEPmzI6EF
krsDY/US1MUUxdjWWAfwOZ7YzEKqbb0Di/LuGkUXwTmBoV8fh8s3uDvKqeftjaAb
hm/k2lMB4BngOyziFhKbiMM4SdHZZgi/2LER+aev73FfHZ5T55bimSCNe2M0pSX6
iQRoYrVdXWv7XR7BlrlRZRZhIkLYykv3UruBp2BqQg2NRO53v9FN7wQRN0+61Va3
gobGdcJTfoDH01BH6EuHrz+0DSCOTn2MpjvTRfT9emlYqfWKtizTiaEkb72pGqTM
gSWvrO8xdUmQL8PHEfvFxoFbML9XUNNrgz9yGdKIDRiWBI/XYDcjct8XSol0va2N
YWoW28hH0nocnjYpDgLQN6CMmYoFVwpLsGoeU8sQQX+UOPtxuxgMc0Dkoj+LyWrV
CGgcVORJW7LY61DtQzPOjqmDjkh86NR3GFsfw5IdzpEdApxqHiVHhOtAo5Tbmx7e
SW2r0E7uNlLTIuk7r8x5+ij3heNH/FIsrcomOhUBfoufBQTmV3qaRsavswZ1tfQw
rroLboveYO+Rrvn75uaAONPGoLY8Ucn9bJG6V0trd6yIL1ej1JIu4u3vfrK66cNB
e+kUADKwuC5BvqTkSJlqP+wMETT0sblufQfnnWozcL74diPd7Zqm+ulUgzfmVIFK
PXGxNcYzOWDh1wawnNH3UG3B8opm5iAPYo7DFUaKHxDJRSbWlzkIv1vQFk1XQiSD
lRx8Pa/6Imk7RCu3etbfsKGoLeO/e1Z82QQR2p6jKi95sVQmE/JHZi5qtsJXjTvU
JZWgMKqj10WDsji6UmGUsEsgu+8oHdxfNccHM8Yu5mv5SwGOhIDYYuKWV1ai4sy4
RXQ15oteQmpONiZJNR0bCfszXMFsiIxkdFiQ72rbap/8gcQhIUDUXxa+kCxNPkIZ
a4iHBUmwdxG2DrkXJ5F0olewcLB109vre7oYYbC8y5ahiyM1mb2i9hOhJ9erYvmE
DqSh+WIHGQqSlsSqoHH9m1rOKLsHdgN8PHIE6qloUf5YWFbCvw5IJ7L+b/2c0P6t
LWDxFBHti/nj/3upi2R3b7USo07KSSr7gWxh+A5d4xLE0DB39Kfu4EX8ULORZasu
iHFM/eUoLtF5y70rGeOQq+T31lwerJ3+aSP6a/NXNuSpiYf6M3sddCx9Rf/Mqc4W
0tyHE5hOxmGLWgA2XBMRubySA4qvg5aZTX/Hi0cqQNUvKA4pqu0PxXJ0IX3X9fgA
OnJiaatmniK/uKRrSKgGuF3YelVTJi2bmLAG9eY3uSHaq4mQO2RCiVGQRjtPpWK2
KqmIXOk3r6yz4wSIiPym+9LcQcB/b+NkhCo5TAAOFF73PUf0PHjDu/L7NfBhaTJT
I+z+U3Lu4nvnDKNf1lXN/2OHubIGoM+REVo2XRAc0SmxXuuglEGYKNDCkQQF2bBm
Ir89sfNncYU/1Yu1tHcd8td8OhGTGd9efVryi6WK19ymWOw+CVv2pRgbGAdaISn6
hVMw3iC0hiCBrmpg6ShuRlNsECLkFQ6tSEdlVQ1vLj61gs1EToNkkK7ZRV4YKl5U
pvcMiXVZuYGTDFSiAKguelj9uKra/AU8kt9ryTagyKhiARl0Qqj3BEjac3b9GZ36
zshC6/NNKmI2C0xH+s5GI0IExjbu8gVCPAG9JZAnfSrCCw+Hpw2Ba6FDvMXjq9fP
0IZzOuGmCh0lLHO9lYEYlLPyZ4MedSJxcuIPnxFwsGtCFTBxR8HzpBOfBY4Ulyw5
gSSVvMkqTvJaK9BJ2KuiKaJQ1vgBaIfSxsVePYYJB4S8cY1RMUbx6QZjjxGLwe+Y
2QMgyPM5YghVXix9gsA8rdIm1TuScVDfIPf+fevbTbBHp6PJGZx5jEh9kT1UkEqB
2+iR9yfuQ/N1BY2+J3XJcfT3TaHLV7qlOsYVCYmN8aYD7oXLlK1XX96MeP/5pJh/
9HwciRYxVx5nZjiKli+Zb+/jqF59yBYhb/GnP+hnOz+OlnkBadTm7V0GvFOdJHaa
ZYRGHal3Ro3ekLY96U9GztEowBZXIUFoyjqM/GkxGHd1thptS1sRH5+fN/RIGXf8
HubcqaIfTQsPRWln/QBM+bfW1WGXx2MmCZNLiXq3zG+dkKiV/bK/FCeULWCghv+7
r0I55cRvhsv5oHUKS73d76eIF7MQTW3rkk6S4666ibx5QouzemAKmIvIZkBq38x0
v9Gz2rcUV5S2T4O1/kgOK5UUy2vkGalEWrZNttMvdF/aDVHz/5tWTW/N3ag2IcVQ
rEelX2EBzcS8hFxVrEJrUOr41dWdAf8BMHUqd6w72wQ33aNzIlEClFvv5sgZeOfT
4piy/3+3GTU0im6XaD1jyr1d1iyxz6w63+CLkl4P2vSfDVGC7WsXt8bo7ypH97+V
cV0mtbnl1L4nSwrKFOjYF6aE7vm6Inz6R+7OVhPXFM6ZZDyo4ez6pfm8KMN0aWPP
K9CMbF27AqN6tcZ3ky/aOXJ/QbGz1aOTzDGN4mdgzFE=
`pragma protect end_protected
