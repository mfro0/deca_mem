// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:45:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
or4mHdZAca7RfyRG4uyeE/NI4Mjz5maC1Bhj1ZMxC3DJ/pngXe/UTDb1TEDQ1joV
wfwmM6aA50CJsL9EOJmtMLjcusXa6lY6CIT2JHQOGgawuCzfu0ceQORJSPxOX8ad
XWOOHQuzIUV2TqSnV8VueBv0uuab9V03AST/zVKgViE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
sL2axmGMcqqR/yKzAiTqToOJWC9WgQ0PfndUpU/O4HpOo5j/zYx7egiMzRplUpXE
UFrPpS6zAMSbTCO624nMG7NgsQmig+6OjxRUTtmChkw91mjy76vK7SL5mZ0yXWcY
LPcTQwgMBguKtD8xMwrzsgjOfpoIFjnUsxJTywazmQWsjTiwt1X+ulkvkD0DgGxL
A8rheq0hfk6+ievxkRxIDMbeFUAMmroYVHvuI2vrRufbM1q2jwpDesNElv9b8G/Y
fxPT/PQr6PVmLCCiSF8YBqPdc/kPY990YEi0npC6oXY73uZhPKMykWgBHB7ANRE3
DkFJvJby+De+XKTqB83ZLTuPQnLdtNBzhYM1MHlucst32dSjxeFzaT1xt20EmlVt
Dr3WAhie4TienUPnnbIkwJvGVfvGgLTEod5pra+XOFbEo2+iU2PXTDRjWrX8En7i
lUQho/zhzrUID8jtGvNEVq0Ji3iUIqsbtJ29bPz3rQSrb2MFDLtUrieH3mCF3eXI
C1m5b0X7zICz+yCTH2fvcTLnhHmZ9mGHeueNq26MuZCgMgsf4PDYbC5vpNAAabPi
HfCy/xKN8TvRbX/m0o0KqR9vHkOff8XS89bLrEGNEhESSg3N6lfw3hk3WEt1vADh
2hFbfWOcrkIpsq8IDfw/fXIJbmMb1GBhtNXw10akWBACArajp5XpTOCktdBgeJnh
E2YN9L/eF1Z3A3xGqdKHgmRPOm3YiTidvZYJvGIEfFoOlFwkFT+BHpzBT0WGrhXs
l03hkK+Q/rgk8VoZWnvKXRAqnriQcEszFMKNadh5gu//5WWW7oSD4eKa6PKtpdIU
lUnjEQfOio6ZJavHhPI0BxmefWc8ZnM1UaKOwlnb2wNWv7hxmVlNSFFJKaF1QJNh
bOuExJCRIuhHIKhjM1RYpGggz9eEGeP6/V2BNxs8ELSStVYI4yA+hHltDwF1kh35
TReozdZYz52idqp2EdJ5VfpbaAzygrLUnakdbsE2bxbOxDIvtAyprAcQkUuV4XWp
lq3nS0Eq7XgflH2TE6LgKGTwCB6hKKBkRfFV6tiwnK7YQtblEhwYcDjhFxC6+pz0
40jiTCj3WopKGLOdLV889TNhVIjmIVRBhWz6bJ4bFs+8R1EIfPM+XhOljZ3EIMiO
I5dqOjOnUvyJs3c8bMMbrU24B81FiduCtlGhHKyf9u+5eo7YzLqlTnm0eWtCT9gx
2SGkrU1uRWBijAybknq0kBbxfILPJIrQNnCM3M237tanxelonKBbOpVFnj0ieQwb
61qiS0U/tC8/ls/pVWnfadQHs2TbjGD63t/9q4B3U/x5RywpjNh9MkA6+0renoiJ
Eln8fXRO/I/8NlhNcPEl7fgXqmzQjean9UEeAm+0fm1FX39m4gugBKInbV1J54BF
9UvRt9DXrjgdkqR7eO11uS0ugTZglHZqD0uR36QcgusnG1CSOKTQf94nVsRif3Uw
ecylS7cpWZ74jUAN6CyxJE9ZtKgC/7GlXuXkhs04tSO84A30fq22uSDK4z917omw
eG9PkWn97WusDSmqTB4iMz3mt3n/W8zghe0Dkc2GUrJSlYGaNjxFxBEhkajxNGpB
pz0JZE/QnRGySYARYDQWQZ2wTqRaIXF89OmbFjgw/uM271lBvNXtejcLgTdE9qRn
6cgUxI+OTx1MAePXENG0Lst2OMg+ybg+eEekItk/tK8Ez9/2xivJF74x1vzet9V6
BBGQVOxIPwWuHzcpVbNezZBuLRWFPLJcgKqcV9alXIVdbeimCEJJi9UFToPFbore
fRamhpi0MorBoWob4+6cBDYJaeawsZCGvzWLQnofjWtFZuGgSwfUiNMbwhtYtKMr
z49AWeHCN46ztJAbQqMVIKWLu53AwPeUuwjt6SEUVbwYJxZsrE+H0/ZVSQGZGNyJ
Rc9n8O/sMiBWG+60bjS/AFM/D+Jme2qk85sD1Mtf3w1MgP2s0c4+nZOPAtZmQNDP
cZC34O5uqgLRyzr0sJL8QWxNDfce0dqB+5JV+KrGmnSDuSMkh0Umx7nRMVrgxjoq
uTAIqDmZqVzSzUydEtjVHLSkyQ2q7gmljC1BUD6HDbL+HqHUukkpMdC9NkZllL0a
x3oHDh+62N6WyRGtdQsEVHf01C5uOKbqdRkgGaNhvMzF2q3MwPfxRZV+kIt4fTym
rE+B/5KvuP+JUw3LimATg+L8UKo3XwmFP07UBlMrU9cGhAnQMXg88BQf8gy672fZ
5dCwFgKFRBtfQnMn7/uW11z6zY89UH23CW18bOOtlLJX6k6DpYQqnyoOGHUtFc2f
CqEu3x5YQFroBgrU3X/UeWd4ef9oMAft0ecwwJRwkn0145TyWhcuCn2WgzrZNmct
vAMoV43WT4bnGX1oDd3aVDVnEWWFPEBOYTIYc3BxFFFe4+2eW/Q1jnGeaZwfQCTh
QlSi48T8MbCxlWlWKb7oC/EtkAf1gWbpM/o03/1Pp886XJZJjm3VLovVH27lriZA
eCHa74ff6RYCnMGvpQfJXVQxA1lxb77Oh7qXVr+Y4nprWZyVH/hHPb4mAJbdm5DV
QzD7tE93QIiouhMcnWhAwUi1DXeO82mQ9vY60qcfu+t49GiYX1dAaqrpVPfHmIzp
0/NWrDsFL17YJ50OnQr/v0A4D94p7QZoZGiY8ZRcSwsv7uG2TsQGlEQIztaHw1NS
LaN0tm5LTpj4KBIDQnUIeW1JyPOiQcZHWyiyVzyz7X/ZEKuuJcErihO7uq4AnBq4
gnc+MVuivbf1lIfTQYDUTU/ypomK3Pvq5NYcpU3cQB1Zz29whvNbrYI/0xW90MYM
EvjZlNS9nUggLeOpvKisKbPPpD9xKCPYyGW7bDHilwJvZrK6Tp31NqimEHjU8GPJ
FjthMBGcxDIcN1rYvyZmhLXIcr1tYX30BTKbv/kcGWn0kPTeojPJn6J9xQCSSlsp
g2A9DmwYWfNGHpJvv72MMnasQc9eu7R0KM6vZ+RO+NUbOLKjl36PssWVLLGBpMK0
W+vC4pqZYe4J0yqkkRWTwX949HnW44Xv4cMwIFE1lU897lumZuzX3lUP9sDTlVrv
eDcoP11xfN/Gcrnm7xa8RLH3z71MQLp7bheIEF7wM5c+uoFoGnvvR/lS2fqCq1Yj
H6XXyRFr+5bajV0+Be6uWu6dJEpf3NGY1i0oCuM+P6yWiE7OCRD5YF6zLMD60vGS
Zr2LV+e/G9UojtcSAk/wplJG7mwgzqgKfpbYf66TPI3yasJEBptRpWU1kH1/HPcL
wut+PZZoz5q61sbuF48Vep6smJaxoKmXlZs/0J1/mHjYfne501JR38Wx/B98yhjc
zpEnwC3yex7sYFU/w3PS7LuMB3aSwIYE6BFI8RKgYWI88laIu4Z34LjRdTPM0JsP
1Djbs5EanS+PxgAvGTDFK/wnhvqv3r3ePKGtU7HssIHQpjk3sXMiKk6pJZ4RKNAT
Ax24jq7KOgBeQlSwqqO853uAY4ocbkcjHpCPnZh0ZhpaFaQAvPaNNXI2IeXwuOGZ
nZR6SWgqmp3d6vvEhDJbGCA+LgTAWzuTYbj0qiMdrjzaPB54LHdPPUwjp67vKJhd
0lX93+7WZx7J9+IKnVPfWcvCsGrnO9ThIsbbCz1XVPf1SBCO42IWBAuU1Lnu6FS6
eS/gbLCIOavsR5eXrdrMBvr0WJ34O4bAgiZhF1gMxjckTplkCzvcxxlGfNvfjq3q
D2TIdoZAjjUTruqVurGwb7Ti14UtcNakFAyg6p8no/pfUycWoZUhsb7YgBXxW+DN
Uvw8M9WOZ0WyQu67FoZrpNQNgl1ozQYNYkCkVJA0f/MldyFO13sFp8TFnzJiR2qL
TkT1t3hRHf+6FPgGhPEJJn/KjYnvhr32C4MQ8pjyGRD+/p5mkF03NTTsfDJiHtha
eAuCRVFe6CpRcdGq92MfLzMCCzB6cRQxE7chCy2S0pYHYVxTZXkaS7wkllWjz1Zi
fvAAqaflvxvC2XyBpdUds8FbhAfGAzfhWZKVIATO32Yq4qPB017Pn5ta0dZZ2u/n
6cqIy8gTn7mq4CtITOXzVxpL5XAi/5BjQd//0AmnswXdYy8hqXKQdEvvHNUk0TOB
/foZ909JPzn0hOIa0ZRe1Z9nJnK9CckMQqr5XJY524+d+EaicH+4NI6olv4zb1KX
PnwDClcilIWdDD3FL64Fmhf6+l5YuQEJliF7G8RLrP043MbsjQYBQje8F6HbZbg5
1cfgjFF7tus3JduFwEBne4XkOSlmz9rKnDyDVhn61XWqbfyIsEbVnUwCVislZ2QS
r9ZxD1iRplmjvaQdOkSU4a0ih7g0/W36kl0mCSRjULh4uAiEWDXmBfH9HeOzMaO8
N7dIrQCaIQTZ7b8ZrVppy/jc+rjTw4OFFG8V27NI43pX7lZKlf+QapZmbnDHxcbW
XsnayFMdYaPMTMDsAy4s53HNavLF3bajIbm4TyGdwq+Rqce6m0s0f855nBMuUQ5Q
690y0RNe/UUp7byLZFGO8+K8PNqr1QR8fMitHqq0RWTQtuPVfPN0ySSK6a300WHe
4l691GsYxD/ftUy4Y9RzcgB/Z9lAnzBbsNxgKJxRFmOMpGTYnuz7soNswoMYvZF7
QrTfyiz/6XFH85GPx0m/qnVUwsYgfpM0oBSNYWnPbasFLdtqidzSRndrnXdgpHgL
uWM6xBZVjJBx+Z1ETkofYrN8voRT79yeaPHtAVo4R2I0qmo9i7svxhFBiQUL1Apr
iDSOhqfxhi4BP/eq5lInLM6254vmwq3QXVXEb5swANS1UinuUqrhnKyHnqtlih4W
Asv6eh+0NPrmINDE7wJtSPmS7gVzISMfUUHbgyoNdDQIZQ+xb3dmxdpENrrrPDMK
rGAoh1+Owocvmn9eWZxXp4hqGp1jMsgrvBT4HWdxqmbabit2yBs84q34zvnEmZkH
1Fsbp2w4DHw4JIP5YvYfH6N5vtumlP7errWcEQGHTXDkdq7kV4XKuN+np7trBUpA
F/9Go0QiypJW6+2HKtaaHUao+v/NQiQCwgk8RgO2p/iNrYR9zpefWQqxwGiqNDU0
cl916SbhSFPpfGVdUjiNBDiC4z9RGSiRLAI6zXMEa/mIj8gXZgSZZBzohycKvtyP
sx7eqS3/dUj0O7G42sOSay5hQT4k0IaK2r/2iJRqmN4zXSNa/hVqWduTwhckGf1/
OM3zuP1YHDIj+Gs8ssz3OXvIsR/+DBIAmACrV6VFNcogyU5lMww5A4HEHaWGynpQ
zqqs8LHvoPx5ekIn1tzvVA4bGJ7F4B0bNVqcG18fmEdVBR55x4ELVpYDU/euMOmZ
hiVEQ+8IjoBJsWAkISetmxvNy/CFAnZupfPdK4klRDfVHGCStbDY0ytuwWZWrbci
hx2eqMxSakkz68U1MvLxz8+RvxFBrPta6LVYjav4q762joT4ZFqXgMMOZzQwAIuJ
FgIieF5L3f8UZW71VH/7dg9khRoh9k+52FIIy+qVoN2nPccq3tPJa1VVmaP6iUpc
azfiOk8J3hHFtKmhGowPEvmP3RDBe0R76RG76wlUN2lbPh9Q/HOggc+/vAAsgGU2
fOlu1z0/9ZbqPlHMilk43dzhzxVl6bIkAKDPDmSlIFGoIJB6TZBstNeiE1XYvaVO
V7uQIW31ZIo09iHPe0fbUEYu+xddh7ntZiIuh7oU4vLFcjynDahuE2zMNLtAINWm
qN8BJmIkNmTC34obH1rkUoq1kUbO6U+VXR581+/HHLYMMGzW0bCb/IClo3feBHD8
SxwiGifeEYOngPB8IZBoGSMKqK/NanpNSaD2QbHoCfB1RDhfxQ9BEqBrjbEfhJz/
uoikaTLyYDVo7hCh6Vl5hzEa/EkykWY2wQ1GxPL5Bb3rLTlb3Z4WTaZI7fKHn5E+
M4JMzs15f86la2hUDG4/Yuqhb7QbCgYGyK1FwxbvvMQOy8KKHrhMRmjdzzqmoOAv
APF/PyvBjbqP2+jS4m/axkSTTipiYZLKKKPTAzgixSHFEdgE6fYjZVlvn1bzMQwy
xrO6e1FxrSkPXVdAC8CJcx/kUYHrMRvxofKcdHuO8xFY1qjcoZd4upqCn3GVZL3X
+zwwMEKSEQub6yHXOBQ0mXgWk7Yt92/RhOMp8SNuMB08fPMiScPRV/jyqeY6z2+F
b44s3tBS+UE6xc6lkxqMh8zi9iHbIo+PlHkIND4c1hkwWm2XhurHFXqeOBVk8Vqy
OJgPhjTB6NKhzHmMbzPJqMctaR6AtoDsJPLs2wMHoXNttD1ho6xPvmi22QSAzL7M
utu42JX8J9iyvEP4z4+RAzX+anbzM6FdIDPgaupsMcaodL4Yot6SLB2151SnVrpY
KM8qOr033GsrH+zbRtNpc3CoTLAmyXDeK7rAImC2ttMDMZ8tbk13VMT2D+A8XNrM
25XZ5cDyRYSzo2j6sWkjVd8wxQQywm6gpan813Oy8yFsOhPEN4brFzjWKqtfDn5l
CJa+XsLhnMC3D4ncNhl+V6MeaPqaPd7FHRYqVPys3bkiC29blyxtdRnPbVFZyJcM
Ak4/ndrTFmV98mIn8/EOmQjJminpfPhIAN74eC2S0b6zygD0U6knGyRcZ1KaAQ+L
8NpBjLmGVbhiL3VEuR5D4Uwd3cxOtnHT7URgS1kUj85CaXk+ZPZnxPJrey353pbW
4RN270L4zy+nd+p3Dw8M3aLK+CKhEBxtfwZ0W14/fFCARYfOIpHTHUxQawxp0gnu
ojV48Uu5J9Ds3drKn2wCYhMeZ6aMiUhbsWkbFVcsBZEzff8fuSWHOi1NBGJ0Sz19
DirMjjYJE3Z3W/iTkBtlbflEaWONZrAclT8pOsJHN8cWkBvgdLc1nJbx1BpY51nP
lCAxCmpfh8TNb1bO6b7uNMImL2OujhrnBAjFK9Dwgjo0KU4zRi7bYhTVbrpAZiAQ
CHAmybvFFg/BbTWSDMtHPgqKuaKaZs2SImHdyhKI88mZE6Z5CLms8xlucU9dw931
g2P9XETqIO4yKGuKfFPAyMwlM2yWj/s/qsOH0K9i/5g7wzC7VUQxx/OpqdqG4k0Q
dWTXHP+Q8WSt/yRjUK24DcJKIntMDvZiZwEkjS1tqhR6D0yY7WoujWncgl30oWTU
ESppECga44JswGESuSKQ0XVYcDKjCBC/iJe9elnAJiGB/2yYtJzIc82FfwJUuqFt
UuhWer7+b78+XEZuU5e5gkXIFQqRbjdpmikUUdqkGINHyopD0ZWTWm5awSpDoy+/
tIgkv8rZRcG8R63PF2KROGi2zkOojW0Ht+n+AtyAnF9dogKAIAwLf7iBOX4E8bKz
WoT4h4soIFYIrAgzGCEzY1bz3Gmig0E6qMFof6GIQQYSQuS7mTGGS2ljhlS/wr3a
Yx02ORneMhA1rNmNDg8is8Duono5BLG2rY2+FpkwwhD6eiu4lTMMv02dxJVbaFTi
vM4Uq42EqVX+oNFa+a/SAKCC8s8D/U5gklgO5wQELQZsETYj3rmsYzB0o25TRa/h
yVsfeOGDc7bCO3FlBV0JYQPB85W0pieqw73ZQ+DOb+LPwMeV0JohC4RRLKjAir/Y
01y/595TwK6d8smem0U2tmx/tgoENtjqSsdF7PSk2ZrtiSqBWomzhGv+MNN1rOtJ
k397251qVM+j9cLkY1wSRVIJI960mRnGV53rI51ZjcJTGxmjCozNTktr3JP1E6Xq
tTXrWf3RmGBPXhObXrBax7VKAst0STDrNOQ2PHKe7ZVJneXyttV/cJDdT9yrAMpc
iO+asZ92bvxfKFC/sS1kActWYkBs9fXTnZeLQ+Kl/YluDSp3vxRMs394twYs5WdC
BslUE+pMTpKB35YphtoswL1XEKhSAHkSh0C3SR7vU7hykC9vIUGSGpA26DR+53e2
9RRjwiN2WZLfnC6o9QiH6rC/NdaWxmu1bwRYtMC0tyiG8tdM8VSW4CfqVTz+5hXt
AOuq0y7ES/7D8QXd73oUwZYtJt9gobCOwgv/EtUttmRM3MaRVJ5sGx+qktQMzPob
iOJb9tV/FBEGug7LBZVEf1CRJtB2tVokw63TIJ4d3wabHX0gpc6xzQlQX50fr5H4
YBamz29RTUj3ZIL0Lym1fyciJNqWC1tRm4rJ3t4o4FdzrIWOoL486Y9USDLQkOjo
Yb4CAymNxa8fZsKaEJ5DUXFjIp4BGH5FQdvU1tUzKqO6APOQpkZJSp1JM9OHW1a6
4z135DytM/li8oyOvfFrTZWfTByWuouNaYk1qgHZd/7b1RpUyGZkMeU54GvsVAfc
RSjOL9rD9SXdsBHXtK96g4OUnwd3Tf8vhrenF1k9KIM4a1YX2jOZLhuWA2jGdfcl
+6gypENZN6xEdddTGv6yTqLMaZCKRhsovxbv763UPUuaCfNnYfYKz3o12FaaDiyF
gCg+5SUibOMt3l8GE1h9lVBF9qthuGl5i6Uizs7bDlMGaNW+pX0Uht8ttpVZGmsS
XV1ujy2+eO1nKs2IRM5RhBG8AN4ITZ0a7PZiN4dwebelUad2YAU/vW9LyDrvNMN9
mn7rLKe7d6lFFmqb7fqQdqn7AqFAdOquMaestCUU+Cjh6qwtim9K07JhRC2AajDp
xV2QxJB7YVnW6yW0uMNB+cuKrq5+DAShk/HRD7qkdDE1JUUG6DCdHV1ecNtETDe0
oUPUgdNcR5Aq/35Ai/YFj6iYuNScEwR1btRJUq1ZC5IO+1notOQlZnxJGlJhBe1R
vvfbN/p9kHU4YhJr9/qJ8EbfQKqdS1kbQ65C2pxRjhW9706EQq/fcXiXJVfhyaul
8ALPgcw/ctLjDtQJ3z9ITV57QGXXiRomO0/2a8Y6T9z8sTFCYbh+txvTiL6YOqtn
ggfDmZTe/cmszeZXY+Fr5x1lzVZAlukfX7HhHpwPLrjEnEQsZdaWGRZQsrleVkFh
0j0JCF/BBvDXxpZKc0Si4F+J1it42xxikwGIExQdP5OOtrIO9yOHwS2s6uvkX43f
uTxYpKW+D60IdwC523n78M8NZrHuSOifeGSghs4HkiMTfJRpJAK+6m2nskb/snpb
HzVOOAG7phn+1BRsn/2JPkOv1eKuJnLS9PHPR7CUdBCcdiosKFlH1s6lMcKL5Pq6
YeJZnMflr7EkC6dgySDgoQluWgp3TLRGP35JdlLP2g201lPI4M17OGBKBYiNIj9h
choaNHnSjuwja6tta5VV5b07spCEJR942Vw1mAid1knaUMDFfuO7sj4LrZgp3A1q
qz9eo/EaLwc+k+otxl4nIxDemP9v0jOYrGv2M4a/fx3GtP1R5YXdksjjPHgZp9x5
Z+J4+mOqMIZMEgGgqXl9CJLhCcdeX3l+TSUxvE3Q3bF6sR9ZVkT/T6w8w6Genm+h
XIA2OZyQGgAXs3bAOZh/yWbi8lquIwvzmTe7G8lEGIKROlMjrqYcK0EVUou+MwOl
WGcvdhi+GX+shUHvmAoLOVAJl5wroujgFCDIdVXSekd0DqHTG1x23wTbcVDnnM2A
r3p1rRgDj0jMcGqy2dGN80VJpayJnW/i0mpH4Ac1+JzPErtiSCSF7geOIJfXbXoF
+hGxHRHJ/itS39JVhNZAmsJU01qqqrmSmZnZWKvQbByaHVQBrhfyM02j8l3/DI5Y
l/zfSIvUEmA29u03cmPea4zMtEVTtC8VEU2gbQPLimAvk/aIZ1EKIT0tIYggQYm7
v0e0JkkPtMzzHDBDceDiWil9YusmOH7pLsd4g3fc6FA6T0umQTy/UgpxXV/cFwLj
m2OPRXN7c6TLH2hDU5n229FxWgfYJO5nUKiVEuJS9rTGfXSZmNMy0yg/2qCAYuOb
7qrWrhsM0ST19JpuxuRbksIr4x59yGEHOGtDXM6ZyGpxlV6vR1ymHdgzMil7dcs5
Gse+hzODo+8m8ygDOH1Loj/uuB9QLPRIeQTlVPLX3XxyIJFVhvrB43SB3/7WzSeR
kpOUSCTnRddoGESU35b9XX/J18OTcZ+hOQRy0uqSXnRDdFfDdHl0/w1wbK6durQC
IJz+nRccx0NXu8Owt+GZ3JniQ8OgniRPFifaLZjdEzLtjwnZ+q4MV0HEC+2GkRXC
rkPXSycpbtkBY4KrZoiop+tuBkl7uxduMXvjmbMHZUlDbYbCClGkJISuQHfiIRqz
A18ADHI9biAqKd6r4DmgN80OB8djq3ODv+q+rEnU+79TK4I6Z8dyBWsvXfh5q+Ka
v2JuDgzWatwss1+NreVLH3ujVKMGGwWmTtWSXz/nXCPp38Nnb3TrQmLHvY3sxONO
mOrdcPwLgeFZxsxSacLSWhFixV2GgNnji+F39rgSsat0dLnSusqzkBAmzFldCPTl
cUHEYdELZH27MRRV51546ilQ5WnL1efB4OCwb+TX7NxLb3dOHMgvwOjT19qb3fp9
jtP2Kp94xkY06jqsGZ+ijSBJiwtbih/C6MXZL/oXwdmsSxPDYOZeXvNvYImFl5x7
PUaLeeN7FWwj+6tyEBMN2PyuSmSmfjMGrCCfo3WSQqKaQbOU+U+bsEq0TG98Jpo1
w+zj7O70yoSiNtt9ZMiTysC+HDTdba/UnMzMbLeofNEMC/l2+9hyT3yqqkYWJnTJ
KzDtQ1Z42+4gALRc+68IEHXD1obYAAOvftGmhnSkJhToKVvz6Z8NpHCWQE4f78Qm
Yhoko1EbP8Q7A8kta/oAV4cW+2hv73Pd5xqgSejsQ3995780QYmglIGuIQnHGU6Q
ll8QmBxn9u4JWylBs7xgzaDth7Khnpc/WVL9PU2GVFV5FCBAINx22cf2j4Os6d7I
y/kAczgvczcLC8lVvubiNCMg3nXKm/6L+DBeQICPmPWyCyYxX4WRAdPSi6r7tUAE
x0W3zzlmsoyQC667aI1bm69ACY4TjGCsrkiBIHCIgYynMODrD6+jfMN5M5zCZEY7
jlsmFrLO+Cw7wB3MnPuRGwBXMTIbmmBDTM90NH5R7dBwOVTRIp/f5vFQIx3442ga
MIH2G87asfydvwAsYNnmzsznQt6GRkMOHcw78Yx1nHvgRtiHdcGyorhXkEKLq9qr
394GA7FwaI9uzT95/lFZH7kfFJAJ64Is3ePcoABvqxT2GBhgioakMG/b1zxvnM3Z
g51P5CrKSXTDtR6pfFH9zXj7Zm3dibGaDqzGMUtGRT6tUJYnz7XpMTLn1baHk1AP
v9UiOrrR+6jwd0Dseg6qSYvYpNJNjW6NzUmDzZqkEzSRQj8X3gfX2moMmJ8esIKs
SN21C2COyC/SYxQW07EfLy+CWM1zl3BsANX7M/kIMs1CRB4xoLsbykaNOIt87sTO
vqYWKzMXFq3q+rUG+4u3MWMhFE/d64zPnxg32Is1F2nVPW2ZxgLtT1LNWRks1PS1
X0uOuZybITPsqwFdqEgw+mFs9Keo2IT7FTnuyriWPIAHhTcrB+1kC/pxHfuYL66b
btUDaJ3FiUCNjqhlkcayEDsotep4xZGak1HRIo/E9Vc1MLEIWQ2Rj6HFZfAGhSIA
tIHdAh1wzajq0diRCQzRSMZlBxhruYo6IprJ1FpQWgsDwB6ReeeICjx0KGjIAAL9
d1RSNxqJTZPkyW9/Mfp+k+ZQDzMvHFsgH8gGa/0tPBz2VPGVaXbISd45ANI+LaW/
mAAFdBKM3Bu93gpRLY0ZaFRgct3xkf17d0AV/0gPKU0swGwovuyYw7YHpg4Lc8RQ
ATi7Bcxuz5oDmzPSCN7+N42jPT+2Q+d1Cc7UJWs7vGFmcWnXHTqZt+PIOFMmkTjh
UlZvo8ieqcCQKjcOKsJYJ85zAd1amTGBoITYuSX7Dez3J1FoTYFC5aR/w7VRa64t
1T5SttXXmdbgOpvCWSufFajKvx0nEv4L3Iz+s98FefTXm6GpmnsJb1bQ47drNhwk
UIJ3ZRH//bJ2m3KK3zjS5HZA5GO7TP+VQNCtvsU7ugj0ZMFd/nD1WMDG63Kuv0vt
l54wMABgMpM/ILOBItZPJ/GDZZxIhjSCuAkFwtOYb4TgV9ye5IDgrXUbm1BHFbdP
Gs8bhx+HVyJILgv8TB+ywaYYHMFYSAI4qexGRNtvk/yNjPxAIgVfinmDPpI5aF9C
J9NLyT5prvsUmWCVYnbTfUKObqwaRVmQ5Jr7QzyH4xGYlrRiME6SHglBK+Px3n1W
UlxnHagqIoEi3+7hvTdE+G0BAstnt1jNXZUZkjs4n+OY2NKiDXOcN1sHywLjFBy6
uxAyLPl5OC/HFLHn6k2RkswwYNyeoRs/zXqPf/HO/zL0jBNV8qzL7FQ7VesYL2bw
QIsHiHlCzyeS+1P/0YVVFkCr2PxBLuaC94gsItgvzRHBo0pZJUXhWxS1C54ymDSF
aLAzzY4Mxw/ZZVajvfSlHulc7KCo+suvmQPj9StmNu4IZHH7dhqTj4j2oyzMHl6V
XCPOCCJXlmYM6hWSCGxL1WR+29+iqk4spm+sbVDBV0XUHVMAHaA6/cG91SXX5k+Z
5uCaeQgsjWhN+ng5svxv5R2n2XYqW2aQpPyOSGpJsYh7aCwM90h+bGbmzvmGWiP+
3eqJ5vfg+dENNgM3VPA0UBG4q8Odqszpma+KyPR+XV34SxhWSBls6R8vjZpkpWdP
yOTQa89sBWh79lT+PKx0Ndr/PI93K19ubXw37b8aq2IdnV4PtGje4Z0nt8SGKlTV
5eGPRqBkSI5vXeEaB1fn3KD8uNScLiLwPoC3zshnqmId2jLJLoKEKVr3IJksgJm0
2Rehsq8tezDQijpO0SsKVzh6hN7Lfx5XEvOgR42PGKpHRk4msTTTR1qyjyp1vFc6
AzdJqtnCIu03A7PsfdDtK3iwfhZYaIWzyoCMrPJIGa3hGbhpky6MJ/C060Hw/MHo
mekYIM48mVroAIbiHZokydxDM8emVqhMpZQmfgegloASD3Hgs0PU/EjVpIFrtIIh
8MsXz2d7D51efC87ciWDl06tdFl/gBUgX5vQ+gFnvb98nrRakI+HCnkWsM0BQdrF
bNSheR3y28oR6u63yMa+zCv4EUY6YqFbVoi1xODVB8eB7i7HxK8jWe+sGqc2U79Z
WJpWix/DbKouTPpz3YteXJEBnfpRBeK3DhXvO5flrkOwnRB4w2cli16VvHegm+p7
R82TCi0WyI2opyaHmbXbO9I+CIUks/APbhmLbwEx/z5PUxgwS52ATOnYCG+SB7HD
2ZpxgKG4V/BXUgUrsHjb5uC3RAqCCEOlKgOmykT8bXVDEdt4LgbeLTwWL0s4IBGk
RQA3I9mc2GoR04Wl6qgxH2LAUAHRqILzi1Inmzut2X32APfiHtGK3+trFAigDwCA
Gr5gX5M4B5gvgr9VlgZNFlNy3xRIm14usWmFJqgKT3xJpGMXZBp8jOvk5G1uRjG1
N/9kCjsCdfHgCscUZkM2jHJSvnMZYQOhq+Xqa0dUKUVp3VG8QNlJOF+jDF0qDT8+
bhfBTNxc0ymXKxsxm+eXdmtO1BjDeVNhmpgILkgngGH6088S5SAlCy23g4CnaABt
8fmrweoIoeF0sPGiPQfwBb991MolJqYOuIosp8GqgujK1lDRUtVuPPc9QI3LgfVp
QRxibF/SsR3VXO0VZDlPmV5atCWLxYaWz9aRK8A1G1P6oqBzcVteRKqq+tf4w0Jb
sznWZvbyjgdGgNwQ7Fb23nYgygmEO/u1vtZGNMDjDIT9c7wEaBTHTB2eqUp24Sia
mFxhP1eJTtHZGrtFl10IlDc7GUqdedy/EqA4IzOZJ5kL1tIKFQUGgiKAdXbZO5M9
N5awrZGw2KlWNQjQoGhEYBDPFX3JQopzWCtlTfNLZl6U2TUHx+TxukrY45+0ix35
E9av2fq7kkBAB3tt8t6/VA7LD3tJBetWckyQl7x3UWgrDRf7RjwdnFbol/DhX4i+
MwNy8NXN+KcdMf9VAea9BN0+coIz3feCnoVXv7cykfvU5IIPngn8eCGxD1vWNN53
bwwJ4lWrVmr6exsJgEVW2UG4etvbGaK8OVmtmW7qrS4wmpjU0iudIdDJHWKiHcyf
9HyyN3TwefXJCG8YQi3r3VwnvmI50vM9VO0/1Yfk6gmhbFDuyXwi5b/eosm++b+S
byRaUc81QZYHb9i0dUVmU5MdfpAygNdlxz65qE6Xx21BQoueJU1QtXbbjDbcq+OY
XsNd/LBfTfuk0rRs7+opYPOrpsTKm2n71rARb9kqN+8Idc4fMNvMJSN6WW5ovnuM
goQeYXVkmLFnYBO2L+2RG+wd6HveMTgl28aEsyLx0NHYWNzso4rbhHvv/rIgPQqB
dMQ4qFeoo0H0xDa6E3niz9Dr1kV5rzFpduwz07EyAfKh2dDC6fO5O4wCVwSCie60
ibfKdwdaiwpTj4opDCdIhThqDjW3OIsnASVooUWC+vh9Yrr86CC7lf+quV/Fdduj
kdQ8Sq2sTUvU9XUfEhlXdUq8GlmjB+w2A0CbI3jP0po1ASLjr9PuHzvNY+hCmutu
BTT0fydTSPIHf85dW36GB83ll8ROHwTB8OJFJez6A2vNB7yyTCuBOXm8IYrbJmp2
2CMFAB5xHSkPRZsworungpHRXSEg4RNh7QdFF1QnpSoF9b4q+6rCQ5LpngXcnfko
g1M5lImYHQzYSbjCKJxBteDD/0vnmETu7VBYuj5p31nxq9FpIgByCPYZBB/M+sUV
1xcE+ukWcbCGYNpnS3ffGfuL2+F/IJGxTWz9yujiAQ6l67RCJzyFwlUipQeL4sKW
L83MmJq0KKzJk7adgx6fXRtJnnMNyRCvPsSANw7wa5m9ktZJBYW4LiMykJjiuTEw
PvyBLK+OIjODYfzGO5i9jQ1uOtC+0L7p/a0ClF1xqTQB2ncNyLBDWwV26lS6WoZ0
Rd3RY9CMQYmMpcKpThqpS6Ut4pL4vH3nvF3cLkg2e7qX151MJ3vCtQBzY990fJNJ
z0XdgJZVdTYvPKH8y4zRbPR9eVidEi6k8CMr9ysPDwVFmGrCPXn0uKC6KSnpewF2
yV97TJCbNyPGJ5yJzKVvlZaMURSgihm8rlD7BllOHY43q6ov+H0/IX0PzLE4QUuq
9qgVW0w672xqf5yUZ1U6MU528Y0rZ0txcEZXt0IAVW4t3a6hIRllLY2NwBhuMLH/
lheck+w7o8GbNp+QcCc8ivCjtYjxsEOP6hLFMpd/E0rjXWv9/48nGms5GiFi5Cse
iOgU9sOqXB7iClx2IFvm2FJFoanZmtrJgNPjSuXWP+QxFLBpZvFpNvMoBC5qHXo2
gPtVol5p9tF7N4tD6C7R9L+Rxrk4ZGyjL22KnUWWN8nb8ftyrG5qooh1gkhcIKJx
fF8K+/g4nNYd5tAW1unDDNGgJaMhNYqRhNujAMZRm2nyFNn1immy7GtQjBUCLZIg
weLMXdgvqjPk2XIVFrl7T9vTGQeWk5zNYUgtln3vAYACsgaS7/+q+HXBHzYrfOgg
kXBs1P9HQnMQ3RHClYkN6GaMx+WPxHV/12UE4iOCEtC70YdH3MQT17uIVlfP7GNB
I9Q9SRH0SatWNwoZNh+wbIHDd59N0zi9SneVC1EIykzq7pYfpcSR3OTkLYsWaYLy
C0VJTe3JuWyD0h5GIozEkrZWc+TvukZRSp7eejsws2p6LEPvfCcADIETa8CtsRgF
DByBDbHa/L5b8bS/D4Y6XDM5yOcMpJvbs7ZxWwdDYHNu+2b1i4+WUft9QTEqh+ND
n3vIPRUpjLb2G5lJ3U9OE/zT/3H1Jqh+XK9t+PpQDcjXJ4MtxU3fkaYcxni0o/fw
HDfbO6vqpQ48fGhGEZYMmjvLVXFCadJQDtYkMhJSXdxbrQd4K30SMi6VY9h1cNSC
01X+Milsl8uWMObM0UdBGyJj3ogr7IDIR/zNtEFKoWlgJPhYPOFwcUFn0pHiVwbr
XOY1jlensTluVc/Ke7yVcz7rWGASJfbCiX6IL+H6LNh77zsNO392NqrU8S3n5q2K
lNOdZi0DgTyBzjOqxu2o8EwX9vyub2sTgyDQO+gA2caL5FxxdPmDxzJkKqGgG+Hh
Ey5HwITo5Y+r1A35+vH6+Zs2YHX6vn7emw/MSn9veulTDCBKfTFO7MPovsed2mEO
FwA+PcalYA8MRDhrZmymw3Vgx34SegDJ5Ris7WqQxQDnUIcxwLV+3/4c14z+kugR
NrcHIGTb1QnkjBGQdLBW8BYQAvxEOAAcWzAMfpBKbZzHshiipyyt0lMjjUsj5YrW
arX4K+6KfBJ6LbCNbounQkmwBKGBVbn1LKYIQzwPRyCqym+i49AdqSDcbcxg8UZb
E7CGXT5z5BbsmAbhTeTwRVzzi6wzbtUwoN6doShCx7FxG8yDlPk/VrYBFAphS6rz
LEyEga/eMgPT4TqQEdlP2NR2QcskAOH03d1fi82i8ptsZLAPtR6GRxH6a/IbUrQQ
yOvxETwwkZ4Tw8K8O7CO9sRp6bGOQdzMCAuvIJ0et4FubF4c1Y5qE4nVhX40lHZG
13dG/fvteFzewGbEQ4HSgNrEA+nEAWX5623XkC1XL6JMJKlt57di/mrlfMiYH3EQ
1VCEVcYIC9C5aadiNMDU4Kn3sr+GCf6DlFO+yDvFuKH2ONSXkFYeXaHyFpu4L2HP
I24bBAagkfpfQxlZj1+rAnDsfRvSxx6WZARUHbrNBXNDoJTuN4ak8gbrpZZzcegK
DKmmFzjzZC42FIjZ28+jF7pCc/4ryKT/LmxU+ZkD/7GYuhciTZt7+uZLaVQs4In0
tZXzPzV09rcFtHgzSCmO9Deu0Rgh8Z2lr00JutMD7pSVRIMw8TP4XZiRTnh4nL4S
tHjRINsPvkWbzG9tudgFrWyXMu77pKD9N7FLb5s9dEWZMXxoX98rTfKaMeO800JG
s0IHyGFMhCe1smyMAQWy11WpMhkAvlFHLKWIP8HvDfisCQtmKvwUteiLpuJGzI+v
1P7P0Sfxh4kkJmoNpVLV71giEizSh8YyHrkB04fz82jfW5OBEjGUJEaj/C1GHyWb
hxZx0oBg9CYm0bcMw5H8ugBYAiYQTGjYzkMTJrgf9QKy/y94FBJt70uAfMwPE3iZ
virboNQN0D3VzY6/ziHTClra70SNB8qNiKlgbz3IFPEBhFHu15/Xv+MUFByWZDqb
Z3GLxLeAY2w9pWFNNasCGuj5KACaCThKJ8VmCJ2S7uQCVAJNq0M7/PQLASbHzOmx
WImtBH5004D0xFYqGsnsHqBP6syy9rFi0lKSZ5bIkhaXJK8Zdql2Lth8QSmlRiL1
1kK3BIE9+2lkRpF2hkHA8zRelXkiF1P8A3/aE5QRSXWMdSo0+AKjICxbYiXbTTou
xYkqIIVvnAMK1i8eZqGIYVOoKaJqu3Ho03F30mM4kvW7I2wx2m5GDi6ZAMtvhm8w
jU/3T6tk96Vz48HP+4BFR3ORdzednauQRDyT7Vs/RmXRD9aT8US6i1w5cka/EBqH
RglGvtKe10pyYfe5+a751UKxlIsGrwVa5/R2/gMDlHc7i9IBjmWKi9brz4mR8cq7
XzH/Rwm1xVOSe1HhUTW8zaNlT6Hxaf94iykmeAK8KOojisN/O7bKJVhEpIoLApOg
9+rm0/5W7r3Kme3QVq+GSH+lKfgmpqDylCvHbN+Wp1r5mBXDsB4/irZYn0zBcJA7
3ycyqsrSjS5E6mi1E1fyVIl8pbJ2oVwHTCWTplzUs7u9FYZK/dQeBiRGb9M//xbQ
fwt02oy5AAp+kwLQTQiA1oqRnsaWT1roxcJce1/rmePHmYWW07D54UD4z3XsYGSZ
IBFX5h2/OIVizraK52wLdqkez4bWxuj0Xl/PN/ijgPyTbBkYP23eT0x2197QeSra
E3xW/QYvCfOfk1rNnlv4j6qHDFvMWk5/KCPRb7Im2mIhMvD386ACJprOoTslIckp
ZVD7Z8Rd9oapNAGKUt6Aqxa553Vc6pIZAwzZSwkfgb0xWelIRtAsjHq5uJB1nDSI
mC74RyseldrAT4MST+ddr/DCPu5Ve2tmRPmf2tyTs4+CVygXKLLNZlSnpARc5kUV
QaxcoiMFzPbAUM4J3XbGXTI0Wm4OQcNKrXJfbh76AwmvOtntXEy3actYjpgSRy24
SWcxEDHGtB0IzeivZ9W9F3jM/8AM65+r0P8Q+rTq5Dh41Lxw5MWg3qbMAJZkzEzT
K5LUZtMplHfMaDyLrcDon/V5tRZy6/lK/nUHCl9Qth27sCbAGR8+xUPsJAjOApYo
9kcgsk36hYfYYevyRGTRCQ5U0gYSYKxLW2hnO8VuGwmNc9vH7xHft6UYNv9CPvZS
YQ5PQuHL2W/O2Ncg84ujLSx1nVDdkxm7kBUbb2iB8W9Ro56t9ojgcFdD7wD+niH0
Qmlq5E6Ct5+GjN2i1ZHb1rM5kRgmWWA93LD8CmEUNZ1Tzm3E9Fb+NLme2cbiNNZR
zodJYJLoUAYsME4vBaFPkYCM6YodCuMSnP4WXqOdaDg1YtXOO2Wcti0z0uovUVTA
HU690vYp3LbQQ6YSDmODjgEqi3kCI7IG+Ssyqd3f9VYZLLrCA/iv8Og01wKRPDxh
hiOej/DLL1MzcAqSx9AW7Q==
`pragma protect end_protected
