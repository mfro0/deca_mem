// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pz+fGb7ain2snyQ1eYlAyMcvildZF3Fq5/CiZZ6CSIjPVM6xkqsi5Px05zujruPt
/zvWhAT1z0gofGDDlzTjHHigsTTe9cz3P7JEcc5i53OiJlVoXBP9xb3KbGd1K8dK
j4ksJnGLLgV9jt2PH3Bk8n2FITsZnhFUWSiAEFh6wAM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 56688)
41aYeXyD9rU6FW6qqSXHPNhX7Q0/MuT5H5xMY5ljuLro23Xg1u0W2p7s1+1X4fb2
Kqaev6ufabDBcRQT+Ji6ia1EdOWMGkE/qJl/VsPGneoekql7Go+dvUkQxa4JzHp6
ZE/HbzitKuHZo32YxqYNJCdIrX+FYT7x3e7bRk7TpWMT1wiIyaNyrOQANJ3grSg+
IflW+DC4abvPVz/BM6Ug+vYU9uHCi/mL44zMKZF1YLRS/+IgIYAxh4t1lfpVO2xg
4jw3OBpZNbwB3lf3PI0Us8pPBUGhg6tUerfiipYHBqpFgQbs+nLjhVj8DJcyKyuO
WKYCdRWNeWeI5a2l/KuNuw7eKUrPA9/K2S6JwWcNSaLK7Jhn7qti10nEecLanTUK
yNVNymEk2DEhvXCGn8I5SjctEs6fusRfUv3Vi1XZqBr+PhKQHj59l1UJ5ycvvehc
vsk4MHOCF9Pw3DTKolj09RZkxcIc10rzTZaJ/WVxoufLZswjVSmr1fRhFx8xM6Ac
0NEzbDz1zborcB/ByfduR8+HLlrWV2WSluK7ciS1ClYb+ZZnvPSbtTdxIcYdNNwi
3HT9BxS8h9ai78RXMkcijKpXwE80uUyymS/Ef2FheqbCfSk0T+xiTaMDJwLPSZ+/
r7xHxhgy4Pbs6czzVSYITTr+jfBRvoXPe18Xs1NPnku7IBggK7wSN/ks9939PwWt
Cn7rqJGpwvTK7AnkRvHeuBi+YhioFfBcihDvjsd/WoSYjhddz2tEBRL3E2o44IPN
eBjL3xLZWCw4X8/dXsIo7bicu+IiBLwdke0HWInXMsi+R+BDkJHtd8UPRK3PjMvI
0lr1RRERTxdA7FXHQ9NPdEKp5S7P3OJeyV+8qmdoiXG+jAOxfU6Y38gNyb0bQpuz
3lP30h4vvxRzgoR0vASaDY4Kq3f3pqFHOReW3vXzZpcWFbKKZ5s8eI+EiWnSVBrI
uovQdRkON1u04YuXwBJW0THVQw06C08P9Zj7C0369Sc9bp+o0S8UjbKTQu48Bh4Z
FmOwOK13sTqw2/YWN2dMX3dMvt6l2vR02GEXDdmpesb0dExAG9hb4Y7VOcNmvEG4
4Ye1d5QWcXUauuhlboLveCYFw1RXcZT9DJ0KXi92/XtTeJl0wmKOXOpiC1A6goqi
phH3Rxi6jIlFAFYYQ4XXCFgIvwQhtfbqbkS2gQuY9/sH5b+0WWdmWh0oE6p8Ud2S
FRlA8z27JTuETs3vWeW4xkn57E3uKuNp3A9nMCyzkn11l4rvkzh/z42QvWJyQAVT
JWvaNdNqr7IKDoaxIyxk9+Nvh+G/cSTMPVFc1oqQ2PvgfvXxqnts8Aw9Xmb0GYhX
D4hLHNn02DAFVR89DbsacYfSftpGecYo9iThx4zKE9H6Rlf05RK7pBfgDBPo4Wjw
vcGbHsSX1WHgnIunwJnFcwbvNnRqUkFA+/UJf/YxBksWRDThlKoW3K1alARn21Ic
adqOUh5oXETXf+HBcD9sbEqNQMV27frkzVnTYCZvDBP+04iGbkTyr1sT/jeyHEhQ
eKqZ6X6PjS07urXuoLkxCsGHgW9FHEaU7xTHk2j1UhktdlWNsiyyiKmacc6OFYdM
AE9DSYSegQAREQuOqWmYq4JVwkfZ+K7HN0QYB/5zoupF2o8nOLriLYHY8MvNnBGq
seRUaTQuEKcGQY+km2ExOTXOD/OzBZxRkH8crEDVFo5mIYTxDGAcPRR3FWRf+V74
o05rU6O0lgJ+Tv5q2qX5VQf7QH6bI9HBVSzv3TEJ2oowrdGdOozvALm1GWSZjSc5
nN2+ktRrdbn8Tj4HVuJ6ZoleV0D1LADGh1BzrZuBSMEwtus3xWarVTncCk4NoJQc
HTBIy7g78cQULAWJcDAzuh9qrB7zXfOuX51TBVYpoMtvw4N4SvGm8yKSh/ftzryg
fWjPMMXXrC4szuHgdOMpUoCNDInwYSYrppbec5nBy+G3Vfpwwc6kADdME/BkWP/N
fF84IQ+pn2fkgD+HozwrO6xXV8JiJHcfpRIBUMukLV90W7Q3ZQhgk/N8fRkOOF+/
yCRN0Aue7LDnCBIv0H8pWX8/H0ZGLJEjtdBX5M3930k152UvXRk7eBX0d8CAG+fD
nJNvrWrLUB0z7ubO/nU2+1hyXPfoRSoh5vDATw10Qcr/GXhUd9WaVAY/nhhY7ZCi
zmZWXf2b9x8F7POYzx8BcdCFfcSIdVYEG9fI3xhu4X9hgD/1ePd9Rw+P4UzsDXzQ
nM8maH6s7S61INIt7iI8j6QDTZfiHIusdbR4UvcJvvStEdR5pronW7PHyQkLZxjs
4VqEJ6Bp39VFegP4mvOuj3JbBh9viZ6lBhZosH6NCVTotqpOGB6rDRukqgwhRHO2
avFcnmUa5bnKUXr5JlFvHCscyK5Qk2Lumd1HWXft/jS5D7k2L4G2ACVPdgwZVNyd
0WMKbZLCKi3DjBxizVSEB092CcIkKnGIoGCA4Tb8mTuDeS99nrNwhiq9Hb1XeDkf
gYh440ASHgui42ueV7yeumVCt73ThuJGDLJRgubnZ9Oik23UqaczGDld6oyQ9SQB
13MEewTAWS9jLUolSG6DL1GVF0yF3H5R0ev4tSS5rqtG010raFOur9iiydPezLEw
mdrV+SiK5j+/Q7/8d6hKKl3oF5jEeBphtysd1MOGUUabe39ZDPONOhz7qJLZ2xc+
gNsQsZMfH3LVDPuEl35RlitSKFbCbNqMiY/DoagNzdpVqVD5qckJgSPKeYiY38n7
j1H+G2P1cdGKd1TZ2DlzIaoYIzNKtPp+Gq6m386jeARrj32njMaB2M0UipbVL49b
GSuWr1Y4vjZE/BEqiFBkoXLmXpycPpa9SL54ongEIy17t66LUBSyPE3UsjlT65oi
7HXYm1Wtfe8wKsoHZgSCRauC+MgARZhrIUurVVQatH3e5RgKYG9rvC6tgC/JmI/L
QWJw26uD2nRZJJ749OpZhsSiacTNTkWvug2sqaHT3w4vLX8r/4sBOKOxmOmknNiQ
oz8dCOQpHC0L8qNvNyKGZXc0PrMGbPY0evYUlcVaIiwfZbhH5NhbI2TyUgHmNhkG
EsakhUVkrA0Ah9El4My40ZGA2M0OjJ7ZfBZBfGJy7BCyvItm+5Z2PRMz1y+mz/a2
eEJZiGweiBkP8ynbU8fNbm8jAT1TajRwGRdnzwDT1vVwghdfPekBG/+FYo2xBJj/
I7ps0Ci3gFR2KmGEeGqj300aHh0s7BJHmDVWv8fbTxqC+exkNw7+9dFsRvByAOco
uyV5IhzGB0b5E+FzM59Tw4sQCYkjp/BkgdE5s5SvRwAQ4MXyh194LAs7E4a1sM+8
Tzf8DvkUk2zQBtnZcScG2HVIWfzNZjPSegJn3gX4UdFMHp1HfJ5DQSsnHBEwjUAb
D31MCgSb2eLpdl+oeTHPpptCoqHZ2VyDCfl2duFxlU8mELl3qCbR4zwD1cMCJiez
Q3EdfZIGsesDutK89QseSbGKTiE0qcirLlxk+koiRjHfeGfbQkZEajrYVgyTQoSS
JuxVV1WMXWT9xlxKUDbBmJnDTs40n/lyhWfV3pNvitkcBWxawTZ7wKHNsnom3oq9
IFARcwDiqyiTn0wWFo9ZM74yASoj7OWrdcw4wo/z+qsvk4r9eMPYkHk5FDkHxDnS
z8EjrjSUs9eFVBL+l7MVffHpl/ZCrhlcoL/hAHnXHh4BA4VswFpK5QtmQ3BXBJJo
b46Sae5RYix5+k/fI1LKvSHd0xQUK9KbaVVclhvlJdBucGt4l/vbTFVo2rxqp/aJ
m92Yp5NPTGWea+f4OI9THb2h5H4g89ZZ4YEi1ODAG2c8VlCNk64B8Til58brn/2n
nxd6zxWM/QdeYkYXUBKaxzDpUOcbUCo++86OVk12oohVrTSS5cWZKaEbjzu+sseQ
JMrg5LLwYOi6MlcpSvy+5CHcBisW+oKYK3fvYkIe0/BSSRgTXN7aryzxftJ3VsmW
TERaYkSp/bwwBSEumcPwUG2DME2ALscXIfTFr0khcc8wn7AdtP/0SwwwXRUJN5+/
p8zIs4H+7ZoZjcW5DDR12YpKTHokII7ZqxTLfzccvo0bTMNAzzERCQ/CKwupaSNU
3YJkJRRLyW4JvqZqxthEKtTQ7wjK1oQ4HmUObUU+Dl0zrxEgBLiE/p7W2Ou/kMdx
zbCWGxIV0LmPohNUKfycsf9I9xEugDRyIzLbwrhbx5HEl9YC0Irx02SH1+6BGAEw
mgX3DmjUKTvZXyR8DLu92VRXF24eTk8J/q0spz//6w3Sa1Ub3N0oyHIYU/79Jmuk
GNEurtu3D7TmCCKs1DnLuLoqWv15ZQ1mk3GncuhAELgQXFRbnTHRjlTEIEJn51uI
19q3xDCrl9i1aSx/nCcZi5EU7Jn/PTI1RRWkfY+Tcp0Wt1OKeLNm9x7Ky7uAiE5d
eJ7UvS+m601vFQ2sjdrDMOCVZ9461pIgKfX61g4/c4bE5/CI8VTy2pA3yXnNDUGd
h+OfZnNMDjUN7698nk7+/8twgrs4xaYjO00yPjoWZp+OXgM1koZL3xDcSB+Kgwgn
9HsYkb61dvpW+CuDZM9uTdkTKgCR7OOGsV9dE2Li9JQCp2tPXYNU2jxBbGhdWP7Z
52v74BEJI/iUiz7qkURFUTPaRPj+/u0RpONT48fi/Uc4xqHp+hewsIozkV1I3K46
Q3s6B8Rm5K/EnTOpV0c0FbwKo0yg+3+9FwcjvyKzaP1JgFSuQa3gdHIx/s7ZQx5m
XPgfKQWXGUE1Hg79CDGx9qOz5FJxwoNx4jYaXLtRrz1HEG6u7VjxFjo1AjGvIb/F
VqK5uMVtb3xxCp8UTvZMcMf3VaQoOHkTbRNIXOA0c5/4m3HDY2EpKN28Ej2zIUV8
vxP18dAx+FMu3lmoQfKUhneWROLW6b0t0uqMaHmwQqnrSClMtDbnJMrBjqrWFM9f
G+gVqUi4TaqFa5BeUpWDjyRBoM+YlOw7PUsQBgV29YuxtE9Od1clY9ya51mDsj2T
HNCF81fwA4OpccNH5i9qPYgOKJEUNMq/v2TBL8GFE45KH56WjdL67pAgk7Hv1r76
xT3Xfl3l4zm8LRUBPdFi1jjUJk33hppuBP2hy6IM0amDFNdneN0ZHd8rqH9h65Pn
d8At9g0NGpSbjLfekzPUZ9O5rmGunRpAc26qevpaNDfZAYQCYXvPj15keJv+5bqS
jP0S7rmJelGswQ3WhFr5Nfk1v4OcmJl5dMz3TOUGEN0U/NvmieOR8AD2dexUgGMD
rpAAMymK2ZSNdY+F51pK4iAZI3sY8KDyE2fmU2TFqueAM7aJ6DUmbLgOLMvNQmIk
WDTkVije6UWuTWrWgDyMKvjpHbjUwiI+J8qbc1L11rE8EXQyALZyso2xAEvw9tyW
IKO6eM0FLO4Mxn/B/IA9mfSCdUz8F/KyAPHpsDQkmqk6CEOxogAP+Tnz9iv6GNJu
s8wfFQ4bW1F087Gg56knbdGBOkSvoayRUtJsfqdQ1OIuq8lW6rzairjW0LtvmQBr
8hr6c0+WuWqFs5mk1yjoIz6FDGQZLFYPXMsZSqKHqIrmVk/soBahEKBY6DIE6q09
VySNDxSq74nLOT9/1PWK4v79w7UHdkE38T17Scop9OBLUvNhc2AUMlIqTZ5vU2RW
48OpP+O2D9+ihBaMowfkKmr2EtaMKEa0u/yOx93o0mmjEZoiNiV6rJHh6gfSR0QM
UDQtt8lwIcwqz1aJ8d8CHEUM/7sS4zo016hTHTLAZTttGFKbSiL47qDsDRPLuA73
VN6cG+rLXkFA3mAO/WAlSL/rHlTgnrEJkgfNPVzNqEcVvEgM7elupd/nqmyEy2ZO
CpGM5tJmew00/C+rHLf5kIN1MoRf8+vQG9sPw+Zz7eUVJ8rdK7dUVahP01y2wYZ0
DzW5akjYQJ/eaxiB8zGJDRzFXe6WoHIWw9iVe1NRHnt+uryzqN2Noh5/fYTOpZQl
Rzw4tB7PoDkA5WcRgJLKDbO5NF9CwmNlffymLLL5PRNzzJicM1sH8T0sEMD2XPoE
WbluqcN3QU1sArKtvvSbKS3IoQ2dLuqd9CE0Zd3+Xbr16wTOCow9vVrnU0Z76at0
/mn5c9bJ1WzLxMMbPg8xh7NZ5K2VY11R+jqmzlBc7v5KOgl+3zYeQr/LlENA+ZGT
BbThku0drTFhbC4VhVes4QWJLj9s13DUt21xggayWd24jI4q6CENQ9O8rJsWzM6X
rvF6aaEOe2YIVEcwAohwnWMGYD8uFvftnsVH2/7io75eQdK76GYYsdyCbkHbHFmD
hKUfCGM5NsbIydgH3w53LWerUZnDlblB9rKeOO1oyQUonQklnyOU1XtDRq0xrAfX
+CmtKpOymCuFlqKjSW6ytL9bpdrk+Whd3GHq3r4cQJTC/OtAWQ4aKGfV7fhMeYtB
vEJL9q52TFqcfJ75oujMDiYLhl4t6nrfAjoHNUkgFXBoPZ+juomLxMkrQe+Bq42f
/2cn+thCxKQtcSB4CruAUKFzbjgmKlIp1Kj2AWzlAOdXmOBKzbdSh2icur7bUaoO
40xoI+sDzwe3kOd1IZ0PCB39tWvu2U1+f85i3StrGD/E6scR1PYwFXVvqmS+l1+k
v3X0fqqOnIAuXE016WWZIJsSI1sKoa9yzV1QOI4FAx0+tBItmWZul9exHtDCyabu
CEu+P0yrqbAQCfJ4c+HpL/fbNbqqKtyqQV53ZD5m1Y0DYTKAHiXA9WWCCzoc+cqq
4eVjNiJvEbOemYhvModmHEM5tMiN48pKf3dNRSa/31ZNz+uZySILi95SSW8+ukam
4rL6KSWVvTZabsq1U2qkMruJqNKbSsuA2Smx4UaemBJ+OTuRGE9NgnDlQwOdxTXM
N4QIQyRUK2JwUs3DQH6JpXIf9uCsLdZggaJ8mEWX89i9kIH3nUkiMzfzfWezTmQG
g0zOvRRX/7aOlLFboU9pdQ4mE/4HboMMjXkM7CO8VsVkSyR8E5GfZAjsFIPK0Gih
1owboZdtD2dRFCw2nM6ft5HHw0RDAs44xEQnazG/JiZ+FxUbvc/Z02xnqxXnEGqe
4kWjaxGoG1DB8NWQX4HsNpcN4nzO31uOaj39rUZcec4nZea73ZJnf7RnGslKcA34
oWJygkGjCuHE0Vuz0XPOGMld4I/qM6Vk2ibGFN9VR0jOcRTwzip/DMQ4bDB1erNc
USLbD5u5gBdD0F1uIudCNFcboFvLAt1gub9GYbiscQqU1a8OrMtRS33aUDWICoWL
wp8tFiBZWhWADsYW9cVDKDAw4mieQwmSRwXBVKyeUXJqriOCiTbaBw99qyzHMM3J
dN0e+h6tfa9nL9LiYI5icEfprlRpwOoCIVkqKevWJpTuL/+JGvtAGM6x03u9p5vn
e6UC58XKbPfOGSOCCUwMda18aeO25CHu+jXdOLtXUOU9aMVAcSZYlvdmeGkCs6it
IUKJjqsJFx5SkSWEqu8UF1uCq5esSKu7iag8gZu90JY8OhGq5ODHb6JwuCEEyFpR
LfNxXarm1P2auh9FppycUYHNCWg7APen693pHXpsx72ivMxznABUxqhM8XhuWbsN
DMpl8njPZfkjCyKW5lRWiK7Rw3ZDqNxCkvGnxBty5SarLpsv/+DuooK4dfEe08oy
yPQrKD/FHcHa5qtAd1YmnUp5W/rujiSFXqJs7Jf5VY7PZ6f9OAx5E8tqMg3M4b3Q
dcH4yUQsBXPtJLa7laaK/3Lc0lcRLsfTG+DBT827wmz8yl3/HMPj2CeHUZ07mNw1
HuapUBq3wbNLERcp012ykXDRbhJ7DBfVD+12FFgvx11gW6TI++/3WJA1JB1g3EkP
bs8kU4tzKktrvyRMSNjvUVmbVzH3Izg8Xc5heakFybm8mM2Md8uX7hZQVCBu/1nz
FtqB3YNpVXjohHF+yosEXHSjxNF26nqFQJd75mulxCwVD49Rb04BAWVnqBA2smzJ
UTDpyVElyHI7x7Lp6q9PC4pLyG8y200oPzKZiEQJebxQhVCHQOD4XhCqWupGz91q
tzwgF19j5hLs/awAEAoNOIjR3hxDP/h9UJ/ulY7tT7MES4/nlndorW4taF/WtQAu
/BJzf9mY4AhmPDFgHHvCFqzCufyJl2ZHj4GUufK5qc8ht4JO+GZ8OBz/nOyFhovP
qoO53HrjjLgi1MaPW2F91f2QMnSGF2SPlEYzFqKlsSPvBvPgLrR7i/ZBqwZDnRE4
cdhTPOj9BtBpDMkthJR2m9zpLeS+RGw90rVeBGTBUWeOtS/trv5LUdVmnT0bc3OJ
aLV2p0WymPJ+DZvG5lRwivXYc9N//KOctHYSUMsYtNT4MxZalSRail/TZDzKZ7Up
TXxh3Ic+YqtyYGydO0WPaNCX6RYWVmxbCuJZ1dMv1SrAN2wLLtDd8rzUl6FBnO7G
yw013hNhv8fdrOPlHJSTCWeaPsKONadiKIUEi4Hx4khkhRSmzm2ZNY62s8wz3Q4Y
AaA2xa4YRXyi/fFza/8RELh7e539GxKSxWoXTJETz+Er4i9F15pm2d7Gbpu3iVwl
qbvWAGqG+1O2x9orZ+bFk59HcyNgeSVE4bkR42xGszG4O0VrCw9nCwKJL4LpMSnI
fUi3NuWvId575FHB06MYBR9LqmrZebPRsg+LcnhmMaEpnEqPI0XPJnP/pTVkypx/
TGQPSJQNbzSsouf+8oj6Vo9fZNBH7UUX7qs3BrwQES3O6fDxTb+DOW+TJA/k4OEg
ZmRVFFAG53u490TH2LPOYnhCAi74SXlByMorTZp2e73Xg6Fnn0js4UtzAOR4FKio
3RS4I562S+OPn1pFEZ/Xg6cUbdh1OWEQ416zoh6H/mSXx8G0GDMUFlAe70ILoNPP
8IUiOcGnhpUkMNLV15pJWJH5TYbqXVfRlOaT5GmRgFLDqpnQiljOb8X9tyckzrBl
8rEIMOoHmJPeguykor8reIRHMLtdbNNsFAEvYB5YFVAzYzO1XddVFMWZ1EVgy9Hk
M5r7qMLpU6laVEAycrmBnYRMFnSvDhMOLw1XHuhs+LzvUUglsXZ85EXwE1zDHZdf
exT7ZN/WtxxyNVmB5HgdIaM4pvqy02hlasloN5UFzvuNVTRSyLoVW2vAgwdH81Ds
PG91BvQgpWuhtvJmM8sbWc2MM2138yELAxZtDFpfF/rEMDG44Em5uK97sA43ADZO
yz+BMMFkmy+yGERg9K5UeGTson/BAB7JDDHgpYTc9/6fWH3qR1xzPQC3QzJBafiG
C+7mparb7Jv29VvZA6uDh6PerOYHQzikrNm6wFPEn/t4XOCmdiwNh04g0AQTsRD5
CYoKA8Nrog7RB4pplHgZ081/yf3EkVcD/lzB7cc/dYqleWafRyiSAAVUdcMcEoA/
omXg6erzkFqUnQF+iXaO4gxR+uZtXdSpmSXDiLdWmBZxqzowcohT7w+lwsFNHknc
VBG1QSuYGwwLS3NU0Qszmw3DHEJd/3AEJgFW0Ug2PdSNxeuQv1cyYlUKOph18+eY
jbsSZSaPcNR7ck1lCkqpQl08yzxdxyddv1DuqCiTrmMc8wfap88bs7NYiN9/4XJT
Wd3QboKr2it8kv6JmJ5OdTkJ0ebLRHPKZiJaI2/gGiqzQ+/u59aKgV7WbOaWZH0e
CA1hl8iNQIlQx6dpSzZ6DYfCueoXekBDFpgIIlQwRbVBWr+cO8V+nd7lczj7/s5A
D6dgROAGjgJQFakEj8ouDGzJ2yRnbRgwYXZsUTU2Wfq/TNqmvJ5Zfk0+Sy+i4rMM
FOFruAs8GFvNKQoawr6M+Ktb0VQF2uKDYfS1JoDkB4QfA5eiNg6zrDft6V68ZKHO
oh9T2jaHvXQW5ygRH9MRmDrke0frOLmEepeexFtpIVylH2gj0AToItA5FjGfaNXW
luv3NaG+rifmnesOYqevsKLlgD8OhfEWZEhodDzpnl5qNwqywNXIftaPrC97D6bQ
rvdq6pFpdQIwG3qJRFA68QKOTKNTGRz4CYexSYDzeh091SG2ivy9Dp4TsL+8MKtf
c2ypnObNvp3x7IY50TEfCeXYWDhD3Tt7kawCH6mV1Qe22JJ4ftzl8z4o4KLRALzM
n1bopxwzVp+GX52UzKwlmn8F+EehEr3nhGg/vg5cbMk4wbLiZV+erXGz5u+0BoKG
S/s1DszVDiau+fAL1zsp9aM3DASRh/dCseTLN8sRkzYTVODJmDmAHYAsrWkUy0MT
cvAHXRUmoEJzwfx3EC0EJoORZvzhrwbtTetGRsgA1GugHUlzfJRS3JiNhLyRd0Uj
aDCrjADjUThbiNujEznk/dZ7A9bYKDv+zyZWwk0yKqpA0NAzHEh209S/VBhKyDHz
fOh+d6b0nMym1c5x0kWMPUM7/sQfMj2RgecvPzvCzocrQpp9G4B2wwxkAdO0rDi9
mOOfEDoPnp64PxWquWK0hdNgJT5IXWkWmkh2HHw6s89kqFRUuBHSy5dt0dQRc5ob
OT+qF9v4f+MCoL2x5eaOI6mVcHXOTU++o9kZ7uli6EYU+fnaOhNHATtjKmlalQPj
IoggIoPj1mM2Lrxh/t7OeJhIi8MjhyWFjDE7OpR3mIl2ttgpH+g16+eVBUy+W7wa
S7/yN8ko5nj23/IzR2duw1gvgliy2/vcHeEB8L6mkK1+LxdFPlFevBBFnVkrw3E2
oFzgIrxXs/lgWBsp6g8wcpNtFbOlYQhnZHsLzZMeBNkqbbqvwNdOG0pYqLhusVXY
5MSEgR+zzMR3JxfRt5q3NBbbr9EDlyH3c58MCve1xkFMqeQG+1wXJqOS4mx8rZ6W
PhPLYeJU0egVWHpohhBgLN5xk9APd+z9dPZuxM8Ym8tps6rW7oEoDqROD7yUBp5b
7EZEyAfjs2c9w8sHKVyyAT4Uo+uOxTx5aBeyNVZ2P/a9ocOrGf7Urh4lrsFOOBGd
Dz3ii1eRwCGl6mUBIxbGndPYz9lzvxaIMn8e3skQLlAGCqK4Vfw7gI8/udlvU8yh
t0s+/IJ9Odsp7qamQkIDhbpWIe2b5ry3wyB3x7JtSfV7lOTcUUF8VXkkZRfpCMT0
mi12PWB0w1NExYrMMTmZZvizASkO3anvMmEpyhuru2fX6+LxyeUJHRR3FmslTIHr
5ujoRMpEVgbUMoPYOpOmItdIArQ9kYPfWMGAyDnlaVJmbi+rJlHCCrpRvDs9cNAd
4qFG6oo2DvwhtD71zYur2WAjqdfgaxsO2MhYodFkAAei4LPYvfJp6LATBHTGtrNa
55VO0GW2oL2PDVj/HjlZmUa37eJnLBI+DiEk7IO0tIe6l0kT9Re3tOCUwfJRo1ub
0IGbCOjxIhadaLgY5tEU+lQESPMj5NeSFcAzOU8iVYQqnrhc9YVZR3Hr9QJkRAcV
B2pnSHmTwT84Lbg5/WTaUHG8iEW40/drVh//jKWXeN/zR5KMXa6hNuCMvsE4nvVa
f8c9rA5KpSCA3CUbkpb7el3a8usMhW4mRjb0f4YB6Ta5iy7IbDPae+ylYA7P3Ofn
Ic61MMsfdrcBdbFWqSc/41q/dIxfW6XeDpORnUqWbRjlKQnrAC4PBdSG75w16iTl
f6HiRGmY6EFazBe8wQWtMO6pWrZVsO2HKUzolU2XxxOOmWLgjaJEfF58N4nfzPY1
WomPL7wMUXrNU0KgHPytHMbpkg39dD31h+huiVF2Be8tNsTTZjLVG7mLyb1t896a
IEBy9miY+MNIdMTlzRSLnKLN8xb+uPRZ0KAiiMugdQdElKs2PMwJyjYjJunQ9F+e
GNcxKyz7WFJleipw6rQRRuELf3e/3fzf6FCAYVClARo23eRLIAo6glbifut6kX96
j5jBxSgP1Hf7xgt929QWSNUBtu5gCCleB6+1KcvJqQmBgs5j5R+hFGYxI+VWoqtj
26IjRbngTFwzAtFCyWidUSKTO1HulweBeFUkD2uge0HALY7JnQy/l7i6+eQJrYxU
Za3OADp0bABjrw7lswM/c3tP799hJbRVPw6QKWp/4HavJQf1ZsnFEF2OMnIW3MCX
lYVyxqn7GH3uJZZ9QJ5GObpCCG53m0Yk7/MJhntt4oaCfMXj4fYce2Ktio8TsrTL
ES0HjOzLcKLY9mqINIWZK5HJIw7CUn4Qi/JM9IoOxOAgsVor9Ky+S/On8TONk+h5
Nk/AbUVQsGrvIo3GmyWA+yuA5mHqZc2uHUYjTw+UG5/3Yb8qYYr2ZOJmAya3y43U
IsTmYzN+V8CF3GwZhRN3wJC1+vd88iUlOatsWCFtJSLOCbUSTHimcgij2wPYmmdz
jjBCCz8NxpsXw/e5jRooFIE8XiHknDqBLAVj0ozfgvla+Y6Rq4AbQ0v/+J6qPR/K
NGSiso/qxz2b6Ujvqk06QIzYoQ/AOSnWfOWGMqHV/oIChhtqMCVV5gpbeCdESG6v
oWUtKFQd5Zy8Dz4/JGBhsDdXRqWSDuBDhXMtku/eQ5AzmC7HhYWYuS5OLtSjXTki
aEUqR18uLjS9MAk+yCiuLS6dVaqy/WZLPlfguI5ndOFk3cDfs3jtVuKr9MkVo6Vl
Ir/LyUFxiwDw46Pafi6/Le2jWTbowrdUP1KD3+ymK4qTW/mUx2bSx0HZhhBbjubL
X8B4P7+C2dmSr2YpxN3ysKS9WGaAeSh2rnJNxemP2oiTsgEUlcu9ms/joHz69Zp9
CfC1lxX+4/5SevmMjE9aoh7Ilm1e1boOGnNGAlPOKdxPaY53bsAMPJrbms2We6NS
YZGIbxClIxb2Kz1gjnzZ5fm1/d8uq447In6XN5ynIoTqgG/yn2ILf6eA9r9iNFS+
0juVewqZ6Io8DOaTnaa8tTx1B5AKnIVb0KlRFb6fzjAzndvOTbg6tGmmhOtUN4J1
kNriYRvb4QExuF2n8VBXXfRzIFDZTAByyGFHr6isPAdFnbdGwhpjo+BEL1tHaZBl
CSfCJEChO5My+4K8lZ+LWjgwUV9o6bIM4UXmepu6+6GJqCq2Dvd0bgdK79LNaVMg
/7XmpmBt2lq/HFzmzezmz+FA/Oy9sQV2tCWrqPqXl8n1kAD7fqwzzj2knjdXR0qT
w9FzNWCWcMmothKjhVYSBWc0EfMWU0FjfI0ooulUTTgBQD0Vswcee7ryh1W8hP9/
0uPm5pIG5t9STVl3GJlvLmtGACv0ofRY92AMvKGccaHoXB+MX0BUXP1L1oRDHr/8
YJcrdGQolo5++ywUZG/40QYTh9rlTT9s7SYFTUxLnZk/zsSJ40HtL2l9h/G5M40e
fKbXgJrC4lyj81GOX7ehTOIlIz2/oObkbf8eT0xLjbf0Os4SlV9RWbfQg+fVFUDD
yHvyMdH3F4l9rUP3lVBGlqaAXSraOBGi4UVeJI3DOGs8nA9tCmKhIVKGLFKYcRJI
GEdk+jPnFzaaK41ZOJpPnUrrXAGrVO9W/QVLdU/NMMQ/+7j3mceHTzL7Y1unB7tT
gkN2QBKPveTCY2zoBaD4O4srWtO36bcLS+F38kZqsPsyY0In9fD6cvz3wvYAhIv+
QRjgTVvoCcfD0ss4xMx+Lky5eTH1i4x+I79l1X4DgP/j551kLtj9ZsPNzYZxApry
XIzQyUyVSOoKD+u0QRjhiQkT6X7zzdhYRSjKAGKzQF4FBhTjAd28vdyHqMwUGEul
lG5KaDr3fi71CfN9/Yu/N2KbSULU55EJGnQ4s7TCaLggmjxMiZb9AJ8HvxhMoPyS
Ty/XNx8o0WzrWE6Cgre7od4YWmzPu4drd9FosakMkl4D/TuFgTotQjcFR1Hk+GOI
XuCFxdOJVBOYlWYKsaTP4RDBcl1lL7Snc93fWISJu4cDVYn7QjrukVBwymbor75Y
DJlhpkr2bDDknDxRglYqzNknoA+2FnUesXKwbxUFBpj+Cp7GFrTvbWl3TcdM4WIY
f263Q/ApwBiOyGVdwx6KeFQhWOtPiuqQ+ZHr+Xu0q0PzOBTqDlUnm6DgBp2Tqg5B
5oVt80C9MywZXsPgVI86eaLemXUoDG4UcVePiRXaIUBMMTY8Vt0qJBDttGX3tRVn
TWQu0WPBIogKBAHS/bZ2/O66Q0fGS6UV/R8o/CsqHkJCPMQqJCWlD5QbymXU5sBD
LbraQcbuKG/H+3v8wuhms+gVcyCriOGpsZZdnR/MU/MMCe20rQzDM2eEnealyZPx
oopGposkeTMU/q6CuxIN/YogtDAgd2LMI7CI6nz/9U5IMcBDP016PFE7Cf5Eh0MO
NeFq5cJK5ftKeL17ATTHKQdhv47CuxrbHPO6HHtFnN+TJyQFuyV6HU2kIXWfp2xp
6szcYwqIYIgKgzZVy7MoxTjKS2LPAGRO558RbibrcMX9BiItB0tZajc3KxSybKJ3
y8xA6ZdDK86QckVkKmDdsb5vYU1JSEXebiOzeLJtN+qqj6Zj8wA/m/SxB2gImUe8
tphatUSOQc5Sjl1SgI1SaBbqnXxEVUWSBXZSs+pIh5VSQF0S9Ie9lDrEV069YlXC
vW/sxM8NL2mH5lsWggcRdasjt2XG1Jjrmi4urrvVrPEjW27CbfsUWDQdWL+InM2O
hulgrmhn4RaKYrBrDJVbVfB8FAiThTt8ChtYXXPETgL6F4jOfIIgrmOGkySDiW2a
n7rTbfay8WCx2bb7XXKo1tWI0X5/N7qXTolc2dPdthnmZJGTF8+mPQKW5LU9hHoN
ahTGWhpQ5VJIb0+G62gXIWuvviFO3Uxbk7Tvqkz7KxxCZ/FSRF3GXKUbixIiP51b
IYC8GsenK+ETiYp0BTFofYNrtDT+u/PgyE4iNCIJxI3jqOqOkY1lzIO8qzlpftjA
2X+J8RWsp2/NrTT3ZTaX6m2ofbL9uEnADAEdkxsaB2f/34h0MJcuq5y9+dDmQxSf
3zBVBnSd2IH1QXS8d6murYRsXXOmND7ua9k7lx2/2lYtwkFXIcpSNB1t/2i4bbuE
0+G6ocPzrXblP+x6kbqli5kI8pCtWX6dDg2hjSwwhYNDrnEcQCM32O9m76uq4sTK
6lYeAbcaFpWSDzkZYwtWvmF7+u85OqMxt8cVu+fFa8gFhkc+g1cfWNhxYNTMUEqY
17xoIxsaI9Co6kaxgV+XGeUmiXb4irntyZvn1ukqoLZ3WCBARxb8cpnzugdMEYd/
cTgAdlVZtsVnkA2E0A7hht5Z42KffmBAs3Um4I4sB6/Ud3RZEwXS/2yMlMkEDB1w
b18XX7dXmnnWo6hBRgFlY8DOOHhfcELV+eR+HP6w/1lYg/VuXEaIOlCbQZCit1bL
OczL+gTNZw40LS1HHtxT/lEnrqmg7cP8m0MJC3aEY3RHdp6A2TXOuNx3iLfBXTxp
CeH7TuJq3wkDgaFvCA9d3zvqWLToaCC0vsV8CaAhch7fmHvt6r/VDMHxBz5kejJp
Jn02JiGXD/5LoD4SzvyINMVc6sV45muSCETwLL5HClk0KMrduV0g97CHAPSx6SRT
HrGwCUT8o6UPPuHprXq85G9IZpYSynNo9E0hK5byGiPAPcDGDl/BSIIS89PwEgJA
XStP9nUIuigvuwSibOJpiOdphoaeAhL+f0ceeEM43U+AiABrvysPeDKxgErbeDkG
4CeTqvlZvCF+UJ862ujycZ2EWptIBMknUfOvr+V5OaIFv4qtbgieRB4oU/YG0EhT
x5ttcdDNlyf0jRboTgUsDgrqMxS+LRr3DRoQv7C9xyMVa7tYKlExhGiOeIFQvU8H
TzmJBdG8QcGYMVtOVDk6trTAe73kBygZ4sN+gyNtyZ/+9B+PtCb1ofekrYba4DDS
VghPJgDfEZenrzg+nnxB0omKKQsXqWg5pVZ3JwpT4hVK8Mx+/OIz0XuNXzilzjk4
NPGyXV7aEvm3gJTnUyT/dhach9tBENyB2hFShZiHCYl+uZwigsd96NuNaZfdq91B
lvbaiITeCJrq0CHpRwPz6/Q3F+k7hKeYtmlhwTU1NPBelpN0ugTbeX31Xt1gcDrL
WxU+PNo7SW4Sf7oCXJcBU8rzcfFw/kzFs6dFytmStxsvMzkNqIrA91+PfCo5sku6
jfbr850sVmHggjMACM+2HtsL1easca+x4R/qz0ZetUfNtgF3SzGs4tGu1CycIqbe
c26NZXDBMgwCoMazrkmuehdzf6DnDmhdsnw5RPmAm5uPl1zxfRmDuziKsqlpEXR+
7Lq73sHGDHA3eLnoEub0CWA4mB+QJHrEQWf0Xx8Ns4spXb5QeB478vjoRSTw3u4m
gcwfAvapr+XM/Z7ZFesVtPkZ/Umv3yU58vClfMhL/mCmt7ffVhE79GAcRElsLc97
EpdjsyOia1/ZKeyLhwsJlROLtsH0k42N+KBWHPZNpJ8ASePOofuBp+v6qiIMHayf
m9jSbstNlzlLYwHhfUblFa5NWSvYBJrP6SfODAeA8brRomKMJtm0NwiDrMLZhgnq
wab6UjOsRiKch/cjqHsG4/SXoYFUlI0TADZW28HGqhYpqp7/v1kRgJ3ZLoA2Qu8n
jJUok05o+Jhe7QwHvMN/KEG+KohaZkFs8zgCA8U9nL2UPu7Vg2MmfV2Nj0PVZK7I
pdGXarwjid19TiGp5eLPiO4AQufaM8q2TA2pTfGX4YVFVh/71L0071X4gCOVMLua
LNFGSsjLx1EGsHkvhLYnXD7n8ydQihbHoyDH/etEMoLlSPjwCRLqHNz6OdPVD0Dt
ftYItmi+v49EMmZz2zVpEKIIgWMJHUUBX5UTOtF53in49OIdTSQFdpaE009NTLTe
Y6BKsmbYf8UbbHUHONt2/3OjH/CfaLrI9MWotUbffHzY+tVIKnZs6r6yehpPSmpm
0JukkweyppGPNctYkYA0CBFt8yJuc3KxsvQ1mSNnY/103vrCJ0CodiGNqiajg46S
dTl141yoO7ct0H0oW6TjeQgpApBvYpKrhTjRAbjKTuwSYVhCGcTNLxsR0ZgnUrjl
RxYY3MIVQOrS0xwD2JVuO7p6es/q2FnNWbaScdoFPrYI5Ch5a3RVnhDHRKxa5IVX
9GoENyzhUHXc2J/qDSPtvrB5JYrxMvtllCoonfBSbv2LdZ4zi97AkvmXuIpkVzwg
hSbb4/IAK1uobMxJ1RtFCTRSPLtO7vQ016OHMF2kSLB+A0B3oorBdNxd2QVdDKwf
eMnXIHS/hD93/OdPUQWHzDFb1Uuy0NVU5/VYOKaKvIGAOc2F2apDBN4OC/PiDkJY
9WD3k2LB3sLqSyXUvE8WTGH/Wo54h+HAXSxCSqE7giSxyLFFiM0g4LeRjMNxCIrG
KcV2mXECwFG1ksQmVx8EH+zo3GwiKN9Qx+qd5JS3bgM0FBjwfK5u6P0Emk/3pni3
IJfRAV9L9OSnRiFhWHy3p5s5+vrBI8UHYnOZVTVZ3mEpIXenhuEGOIPCR97nltB5
3JNu0MievDyjw0aTXJBanJ1BvH04KXZ8V25HYAbOUJPER6OQ1+4N1HrOmSQWMmvl
Ph72VA1xyvgDEtU588TPj5jK61iCQgbF35c5FDFb4y058NMKqiAxGsO2kJvgUIFy
n/j8UDKPN3+ZmqyZr/udxUq1ibmqGpcJb4KQy9oUZ/6YJxjVNaSFkdJxTzNj7J9j
dO5ampJHuDy2+TTBLh0lzGXtaF7GMulMWo2I++kEKIFpbyAR7AGtBeHm7bnleGXV
4CWwouXQQ8oqqtLHkQLb9VAnQVe9kt6hEoRf2GMer0SCKnoLqEMSw1FMBLxKAQps
NND9uuycI0NaD03OEl++3WSE1Qx3vd2DZi8o0l3V/801nGvsytkAQgQ5/f6pZ73h
LnYQwF49kblBz30B5qlgpL5Wwcxa2zJOrEV3Mh8CzWcx27TBRoAUFyoC7ymzRipq
LJtWrZXc2Gep3KjZ7LsUO35VE82RzRpM94QJiTyFtnJWEYjHw5XD07mO2DBxVYqI
qSNA7Pgt4NjCta+SQGFxv2ZDwz4LCqfsPv+r5RMRk/tzlm2wyy0qzjTepjhT2vfJ
AW3IY8S2JYBdUlZlwbBtXTI+VfjI1xdyW9ICuhtPMffdb3GF4oo8VCxoCqY/REJE
Jp83tqRaa3UXek7TzjJmcDYBl0D7+evWorDXO8+7DCfFZI3w0oMFU+M3pCJO/dPl
JWrMkna90MKELOoDqS2Pf38UacI6XV7/jfJ8tGL4uJ4li5/WB5PVnlBt6XZ4CYWG
/yzswftKI3Aa6tIjjcpsBMHCfCmTMcFNj3yvd51GHNK/E+5ZERxPYKeB4awcvuAa
rWffnEBYiPny2dX7mhqwmr0+T/lKBLIUENk4rEUiVQt5B+ggFjC9TurTYvZj7Bf9
z0+0e4fHMUHiHrS42xRhVqyQL55ahAp0fJ/E1xjNe7Awy8Jaq+hcR42WIh4upiY0
huEtRi0I0xTvO8hDbFfa+ukaG2GBS6OCigLz+ehJnjSM/T30Hf7sxoCvb2BGmZVD
u5LNgdStLRVk7svefgA0F3ZkkqvH18mX3Ob1Jg/1CHPPOS+itocPsTeRbIGCkaaO
XOlkhT9eHqUIu2vl3614AB5X7xxWe4GW6XY/wK0Yk2tRAsY1oPWK3XelqKPHuc7x
9BuCFb1dpHAa5oIBQlOVUL9eTRxPe1t97c09b1tfDu0mnnKj+0/wteIcxC1Kyj6G
FAM7oICqS78DsPIu3BhlWocINzsA6pytNsqAumupuMMdDZypyJEY3Nz9/fK/pDA4
XnZxmfbdOJbYmHVxFnbm110SB148MkRBTK3h5PLb71qDg/biiyHA0u/BHLU25QJi
rtRnpFcpr120A77Ha5FdyP3UGJ7sLoMPS2ho3LmI6G48tXTOWsUNRIzKXd5dFxI+
+wZ1168dcxHynECEhqh3V6xJCY3KHJ5k4LsS+RktUvCGEa5Xv7kdt5QhNloZz4lB
f5bhpiFpMLub7IQjDjarBkOJ5UkTjJGVlMelbjMF0u0CZaWwwtIOKraJLJ97HDSy
FW6vobz2JGCyhUa1VJqwFRuQ/sNF2cQ/CzuYQCz9E4D/BqIoRK3AZ9chgOLkIa/T
1ZR1eY7l2JwfnbNdB8jEoUJ0nZhgynnq8a1d43yQbqBRcp0fhQW18qR/zN1LKpPX
UqOgpQpK+7JQaMyr/1ukIGi2BEbXi/aSVbVN/Fpz/m6b8nUYvEv58mEgaAUb4AUE
O6T/HV7Q1SxEJmNEEuWZrt9OyywdImicgozR7haPp6c/aXYB7N7P6uOCgRI3KHPG
qe7tm5Fq/fs1wI45OAK4zqdL8hld8QCJXREg0wqK560ZI0SkT7qFzM3t3DpcjWaU
VtVmMU15FkdnI0qrTM8oDSjvWqNzV+bevvyLdmYadZjnhQAXTY5enFMlEZPC0Lo1
6P08woZ4R442FBi0pXoionXgCYs1l4TZ7qhDNYjTU2z2aLFn9QLbEYR+nMGUs8ht
tsdFYg9wxXuiRF98oN48veSHjZZ8+GvnVNlLQ7NummhDrEWUr3VPFfqwhQv2tICs
CoqiP5/Bl39LG4T2yULGcTG/MsXv6O9lMZ2PEqMjkh8UtXgtSlbUpl2dU//cn7Tc
PE+cB2FJOA0aoI4E6OHedrWczplLaISDz5a6yIAggfxY4wgmvVr/z407OAed8lG5
zOHkM4Y58t2tHNv3mqI8o+wL9V5BDQNw3iBuN7XU06zzVq4X+fpgPyDaqyhAVukt
Ykn3vv7UKMFe1wp9rWdtPf2HSPrvy5cve9qn7P5I6J2XVS++Pov+ScGzswVWQ8WN
3gct74dB2Hc4UsspvdU912i+KIlAgmSIb343nEuAT+q7EErnE2amWbXy88cb9E4+
wB7o0OJVgZG83InC4cSsnnTsySF1yuHdUlDVpGuGC6VemLkYjEylYOW1lk2Ftuvi
91geNq94OIeSR9wLpq+BBl2OlwaD7BO7TjQL7EANr+Jj6HXdjIqQTrCwwN2hm2cW
Ga30Csi7ACKr6yKmMtQAAR4xu7zOgbadayKb33RBBQw1WIMWW/2VZhWYu7U5VKSw
Eeh9XvDe4aLT+6HJ5wLnRQ2ekdJ1NEwDk8G//G8TsAoMOTw4c70st++nPC2pVhMl
84sR0JViTM0aIgMARTusHmz5N/Ydl2grvU0eWOXQWyxcEQq7L8LL/7iDZ4EMo9fR
LoVSB7/S8xhYC57X+NBiMwGwmUTkAH81FYpviG4u0F3nkced4NRPWJIXRrIWpj0+
2SOcQR9fnIvBku1mCNLcWGTc2Po5H+wniPkOUcvvtTP8gmWKjBD4PUjIXWFeFylG
D310B/KbA6+vZAU4bAp/mxsIfjIymcGmqFlffQBZWa8Eo7EVpbpB+MB9aSzq1Alm
/9uRsv8ZbpXyuICgcxBzPuKC0CYvkVC2Ep4uMlv61Rov0/S/ijPE2dBPZLEkqJ+l
Uf8r+bm61AFswaNVbwa2ci//+Wwh7Z+7FdhfO2ZbsUoTQCOV7G6kuTT+Fsv+V+fd
x9Mz/IaYXBc0fU93FzsaLMY/iWr9/Ze4oH+dhHcm2LE1nc3hAIETsKYv6BB2VL+n
N6Iv6lMHXgcYO6/irMIkT+ZhIUb3ulOJdI5sfOTZ1dJXTsNoc68aG8MKPUXWDXEl
fNX7+i/PdsU5csg6KWFzqbQjYDVZ1dDrT1VzB2svPozt5qThW+MzZPhwyFeCmtxJ
Yx66Yn9ruX8Faoh6WYcVa4dkN3ncaxeJABFPkEizy3S6bawnH6/E8GZnuornsSyB
F/k6RO6ZrS4LyNgIqdEihcTcLthcPrHjah84pOiWZmZiLByzzW9Xu/fUSYSqRKBe
5WysV3TxQxbrPWShjKq8vDGI8FWy+dL8vy4sbS3BdV8vklZNVUVhAO8EzsUfs85G
oiYQ2FkdT1vs0nnGmIIRItDsYSmnxHZ9VzUtNeO+zMHXYphj0I2JzKcFeb8z28WQ
D0rOKbGRjBy4bzyReRi7GoO+ILz9F7nRMffcxj47WezusqCGdr2hML/GxKLXXfus
GLbXu9FOCaAIjrC9WlVUYF7gZTStqXahwniEoTwTVvavUhAJH+GCi2uAgnJH5kA/
caAFheOJkjuK4gWA+lfnfKiyO6It3tl5I00WH5ZUds5OBk3QrLK+jrnxyH3698cU
R2toL2v5tgLuoOMmFaFxNdLNtrL2DGWZ8ia051SpLgDoav87g6QG2k7dLJmyMKAY
bKcwDRI9T8JtED7PD3uz7HZfyY30PF3/lTJWYsgSSdLXh/fNo8UU5zzn6DVg80Lx
P8GQFzVDOfwhwuCSmbnykFVpOXp154ze39abosotluG+VAP+svk92xiehLWG/NLq
gScCBI9upnWmPR9/viaJogvRSFVfAXDtoN6nbIkmOEyQiFiXLm+5zJS70H1G/2IY
/R8s2QdrAx5L3DHTM/7ddByxGgLuvVUUNs+1oLw9cGhgAFD19nEdXHBEe+opjFAZ
umM6gsITM80roULw8dpxhun6jbiqJW01dOQaT07vhWZZRu9jIKMD/qGT9Wrchx6V
ZENE4k34GwXqtzPAso+5c+D+VH1J1npygUwoYio0gTzUdg1e8Vq8n9TIXXym38m9
VS5nkm29nsdZCaW1eeih9MH+aZlEC+u6eUWrq662yO3cxtNxRwQUIm6TXzsB73Ap
NV66icIun8/EY++2pAyd7t5dISRNHweOIPrHO0OuGFdphM+M5Z/5FI5WGqeaqWjT
6aIkdeeok0cCOkjM67RtBKZMV64i5fhzWjdN4Uc0MqsuoCcLBgOl+YnJTHipn9Ka
O86mzOsCJc1EEi3YCustyxK4bcjjh2hZTlHn0Vs0qzhHh3d/RJapRgrWYZi9CbAO
LyArgykq/VrrwvAqbqJlty8Q6wTbv2Y3Fs7mnJgVnOzB2NoJib26YdmUMOxYyEC+
2Yv3qi2JiAg6r5JDhVr9E7qwsy1UtY3IjjmRKOzZaXi5AaADwugz4fa1FF0crBF6
cVQzhpw+vA5Hd0D9YY5Hw2oseedH2vkhkGVmhM71pxQQuoL6gN55eY9M2Y1LTxrC
4U3+uR19l+kOaC1uDqjTGSZra+LTVudvaJq4ndYNCGvQ5EvHx3hDgVaaT0RSiVh6
VwoTRXmjfMx5AeJ2sVu5RbVTMu6rLyLVdpppbG+6LoPyGFDgOP+Pj3WyTnpXHus7
oi8HyeqMyF+St6rJU1VJHD9v6uTRJbkyWrfFfToOUPPKdDCuwDJ6qOViMRb+28o0
zc5oBh8QyXCpIBDfHZqK5Ok0CPcck4eAAoLmqg6DT1pDvhAAQe/XCdLhyiAeadrE
DaG1NVz0G9Wc4oPetjsKcHacLBNtJR5gVC+hasfXmBr74T+pKi75k+GG/6wmUuXg
gTrFbzlAxpnTQf42rikhGXtRnGu6Esa/z+IPPHtxcXxUmLFr/NHun+y9uG5zFXs1
yOSl3FMnyJ9htuTZSd015LU8S6txraYjYrfuFXPUIHNyx5tYZFwpnSSAMaRGPb49
qorv65AUqQ7vCYOS3iZ3IF/wa3mAhDFM8hUVJvTZQ8seLJ+tKvnPmguitniKGElv
+1ekJedW3dVbLMQ/x4any/rgl5dth8QfKJ0ozqPdugtZvLhWQjVZkMc9VZ+OIgAU
5U6u2m4TEIo8KX8a/XaKRuYCt+sICtQc9MkcyFHQM+NOpbycwLDEMgI4sbJ/+ac2
M78fA4ptvpdGriJ4MMyVEb/v4AWCIdDqiNUMzA3GJ5Zdu9DEoNMWwGB2/agb51RM
T2PQ+NGP6Py2+W87JQT0f+1PxIKV9ReFmOs+ik4K4in02ay6cORUWtTQyRPh57FZ
MF8KChTmxjSwiNF3KXWYi9kAXgt7b5+s6KrCRoMaXODF0ngPUbLgLqI7gNn1wQL7
+zVm4F8IE6XUhrBOCV9J1Rbb3I8lgrNaETPDsOeL0XK5SJLpF48A7jfO3HzWo2X2
CppSbr+eXFY1im/DmaxaO9tndbR1tZfmnNOhOgOHky0ZfG96ZMmhYScuMPXqrpuK
62TogdU43dm/9xgbb0WpzwE0ux6SrgCkSImKn8OlPUh5uMoJjfdmsZlGvGJApVmk
zBxl/rH0Od9NZ9a+wciJxTCcp+vlGNV3BAN0y5llPKroAjajW55erDo5GpLtK0sz
0CLuPlW0dDt5ByE4DsCxGVW/n4q1n62VginXoWaiIxghlX6vPMuUcDB4571kmbU6
jCsJOaK/i6sRwVrN12hfCZlxj939CWVs7LNPVUXJfMNoKholp4Xih/RFqH6txKDJ
1MiR+TKtszOwwqJxsfXTxTjjTmovqw7hzebErFVRsiY5awSksGoq5iubxx7Sn1E3
eK4pRgeXETzb6MwQlD/gRgMlbRelmFROoQn8LIuUeYu4LQrRKkg4RLHnKzCMbTr/
oLSy4HeHlRnGWtzA8Ms1VibcEXcV5sYb6JKleyvplJwe3RKVkdlhOSDPTzp1R2og
dQTWoGBTmlUvSWN6S0iEkIEh7kpGY6vbW41IzqzJzkHZ2Pcgq65JGNfzARvoGrmJ
BSkG9pJNKUTLoyS+UeDdMD0yvYyYgnBg8TWnTJgP5PC8U+eAr0emSj1XK4LvQ2Lg
F684Hpdwo7KLWPbSp2KjzIb8pU0H9lU81FAyvaAM4FW2uD7WyGWvWIWKIlx1gc68
eBOEcGaxvCqlzUVvjubCJEoUDCLDMWFuKpdN4h5Uncn8jRAaLcCaMCqp2bjLKuez
xNAMvi4/O4H92O7GhOWwI5t+F9dPAFPfEeCjp5o1CdbJpXgZWUHtmHX3sa4aA6BI
PdOnsXjbZKNOPNrUXPCS1dIED3z/XHBrqhWWJulZP7WglpaomNerJgIkWcwObbMq
tD71Xnxoz/50c/EBLzO3qNYbW140V/o6odj0552fFo0HS0l+WwtU4OugmDwjF8n6
dpuutVy7ZJGp+AiVki2DNH/Sb6iknJnXQqC5CXq1K72uK4ETPQlhpOEJQQ0rcxf/
VvQreMhGhrLVH0vn6yuq053kWvc1U+XDdC8JKk7GiWJtVA3qajnakCqIc4yXEhKA
dqOLBkK/CrQerYLWEt/MnMNCf3Cm5yeEIJaY5XhOD1e1WvgNUdkXi7KCYxRZVJqn
zbv6t1uwDqpbl0K2Lp1ogpviINzUkYQ9nKPCHIJopF/hJafoq6wKLhQN0vHZf/eX
xHXUSm6NUGLNoS4ngtPNPcMv/0P+gKfDiMNc+DWVtzv907DQ0eUpT2E8NN1YwLe3
SS0G9SgMrDWgCI8RJePcyNtqw7/cQWOCvTCEmCUnCang7/mLZciLA1OgtqFqNbvd
70EMariGKK3BU5klAo1s3R6kHOKpyDoGX/+9EiaK+8FpAr1WAMnFxqQHrJ2qCI2c
VKcnViJwhK3eeezCXBmzy1BQOUwz3Ymbv2usVDec7YKR3cAoo5N3cNVMLOVCTmsY
5605u8c318NZF1hkUgWX2bVOY0Qhx4X67zsMWJdpn3F0XIgc+rQtwd7LOfp4NJcF
27wPigzA8gEjxkPRjL85HCtBOpubdBJSJC0ldQ+mUJbm/iJMx/rrWehvDi9zO3yq
WQ2wJeccUv4V/KWXVXE1RkDBqAav19DjUtgNv9IjXcsZNPl4m6jf3234dgeAaLsP
OACy2WuDId7lcUEOoUp7XDCHQWTfSflG9m+B5LvbA4DKorVOvKQ8PGVu0E2uqHao
ymsua3ImXxFLGG0nkmK1x810RYHP7h1HcanQSI6z6C5f3I/tgyC7TR3Cif9maDtM
Y2sDfkk2fiwsSB7ap4Sikk05CZv/TJiZ0ES05U+K0pwuvRiEpW0iYFqX2i8HLyxt
Nz7LChijTZ9BZ5610aO1scN0nbyFSXMWQEl1mmTwT12c90uBJrp0q3dOQAQYAsET
5XtY3DOYpAgNLk3HBODxFw7NQEAHd/rG9KdGVvJGDWtIUUjKw61yPxzZxrdPChNN
R+S73kdo54IElBplKV+V5oRrqykUHWvN+2fa6Pn/Ncmh0wpR1dz3N1xgEX55uYQo
epp28hIkaWKZX93YhjCKkcnuXIDma2JFTw2KwCTRpahuW6Ur0LTKdTt2vBvq/xQH
kT3WDow3SLF5+GeKPUt3e+FOD1RzfqsnoqkH29tf5PKJbMoRn7vAUAyBHrdfj0o6
9qTHeVcAqtTxTEK7MlEHGIn7gJShRZ9acW1stWaK2C4iIJocwfvmIlRBEouwESDq
P+v9RDyZbWlUsSf0BAOkIMYlGw543BcC0/Z1V5QzpoJtrZMINFk+ll9/dneTu+Qq
YkaN4pCDOGVebSjH4iwZEeTNZVmSSFagNLSrIBvhGyDPNyWfYf1NspSCrxlspNJd
FwWsTvcgEsd/gnj0w2IJv0ZM+IvgZR8Q/N+nbCLgxImbj60O51/vpcZ8720hGyWP
d4X2fYX0VVeT6PYW1DNZhvKkeLyePEdsMfjLHbVvfuLYBOt5tzdih8YeWgRHlBf6
UY8s954UpLyl1hAB+r3hevzgE/S/DSslcKYjbVZzSe3Z8XTuT1iMBj/OZWkjP2pk
YU131beRiODJSF4ZnkNy5QhwNF+UewcwXGBB8Sl+lU6hH4RmNDsACb7SrhLHnqWr
2YfPb6UpcFSQsMQuRw7K/MyUcmb42/FAK0hRDNBHEXeKfobb/a+rPCk9lAeTYGPq
GX/Po9sAI/OMoJ1bPrK+0JTA65SjQx3avsEiiw7IP1iRaGJHR7WPr3riupE2kbMB
Aue94Hqh1XMkvPQTjxttWMzFIQkm0YOb5B+gHZXKYRXw/+fxzZaFsdzhGqHgYCXI
y+EqCJlqIB6bL2fqGyC9ElLC5O1ZXCaqAEkLO40IDz/M++AzbD9vrR/etmstJ5eL
57Dmf3EzH6KRdtr8lk28OHhb7Xwl1biZPzRENg8oEbw54fAllLRxgVn8Vb9deM9v
OtqCTED5OhHVdKwmiWfIltdNdu9CBMugFIa8vXICKw7p7uA8VZvitQfTwr7bnZ4W
Ij77mc4Ab0nWFvgGVLOykOWPCNkjsPEITPzlZeXdSXSabS67yX/Jxr5x8DM0oak4
6lV9Q5TJyBTWTSM5nbWt8DdVBlUkDFhdcgTnRWbwDhez1aC8cJBBFMul9bGzJgH3
7UxcIyKvzoVFlfoVjPr4hUM3R10F37IVIGn5qfiM+MzMTFj0BAaVXKotBKq5shim
YHFDEprj8khBSxe8AvPso5zTLbqwhm6vzl2MrXW5w3h9b2FwTVQicIVSJCrBqH8B
BlxutcwNEFSQb2/E8zQQfDeKH6hMq1Gl+uTsU8dMEJdY/jPjsxj/MjDzCFBk1MZE
tqNHB6TSnzeLESQfIcEq26kFqbKnewHnA6j3yOHlBXs1CwLadKf7nWQuQ+ND1w5p
g7Rb075JxkbRyqBGTym+O6CueBGUGBJGdRLpO1FKiKPDL/Iqk2KzDhTfGZOxsaQH
YGPSiidQ860hfGA0eEeqiF9Ho2A4zPFtQsfbBG78k3KniMXeNPpXxnVPCxYtixrr
lgxGM+QicDFNSaWlyDnZpq1iOKqHB60VfotwnTT640Rni0HhVJX718DBIiupRGDj
vLOrzuLJgiqwtRa1Gv8l2soBYxxp62KBFIX507AnYmJ7TUrtn3rbltQuc1iNa/bF
k10w2o31Adx+oby0laYDJXwtfn4hr6ql3MMxEM1ku+k+uSPk01rNYV1dBUr0rlYb
bKVtjACD232BYbQJk99MUlPw3Qe7/si0HHJm7Uv26uuGE9OZdrUFEdDsLp+SgdM0
RcO9aHQ2kSLK3SUYAMPkBNdeII4Ftlnzj6hlox+rNoljdQ5AY1EC9yNgxk3P+Gew
tuOGYYg1F8C+5RKK2JmP1/1JZTpgmk7uVAshw0DXa3HyxVaTJeHFjxt1hUpP+fOU
De2n7cYP+xwTecnO1jz7LxFfz1ATRciqYLiKJTWptwA3I+I5qAU+gigPXcKeNi0x
oHE3AHAL+mYjTjRkPZdzbtpVq2GRUMz5uoWYmeLikHU1mNYwcfsNOBhMV3vAt956
G3uYOYvTUdSuwMit5j+8C4TgqLJIi0c1+4PZTAB8yi/F1Ewj+XtdRzf6F08fNLZ/
BlsPlcBYKvpUbg1g1bTbnJ8Yjq/rqWBuETawMndWM5xU33RZjBii++PC84p1BnFf
8ed6xV/zxrsdqD1vfnFOyP34wqDITagoBwj58sTS3e5LhPmorXvgeLF4DmYF9iVb
K+AqXVwe21qSq6OOhvkRyhx1nG97azU2UEf5TqXNQjih/DUyAmvWl9mO5aZ+zGtW
zcuBOnxLjRmUbyjNyyRJ+g7gh9l3Su8rjRPnoefAxyt/5v4eE1F9WAXRRb8xqGHB
sQ9TpBBLCN42r+MLcTdjG2cKBIa6D83haEGqmrmAGXJz+91RgSCmpmwXhdICPuM9
0zMHu1wKS/Jh/Jt3OiBTC+e2DMoAf2quwPZ5pdXUALAj0l19SHuj/oEMk8qeHu23
g+7CpqTWCdFU3uDuEvKK3RZ/s/A+2HfMNbvswkKTM/A0V227hr2+661lcOJucFHA
RjG8fDHGD8fsfrAc93m7WcsAHc0aZESizCNPa2oCFn02cjNb7vbgAzDc3ZgdCO4r
N65IDKFThjPFJjgvwgAouGJfgyGYnMDhTjs7rKDhgEzY1f7uj30m6G8L5ZnrN4WE
W7DWrhk2uhs34xOmKWGcGDeKBZBq/vAnNRAjgB98rglkuuhtSwiQPgN1jmFxDrdH
e8V2tbQB520hPyOB+JmQnAlwus18pWp10UlBtevmICQhUc1GKpyvVoOo0n+xlDIS
VIPeRk6RxIqbxomC07gnnUG9an/EVLAZYo4jecRfyQhO8RfIPlWByTmrmjBMykBY
8584DpCJ52Krm8vBYhNE5bFthcZtdkVGlEf4AdVOZSULceZcpo4l06LQUNoTbe7C
IW65YFpQwX/AZENXcdLDzzA8G0qy8Y4QNwxlqD0eil7hkSOjXr4TLI5eGy6qqqkZ
ZX61OkKgXguymJ7ujVzDcsg/QHBfLidSqE13qHNPU4tBb6jm7SPrxpbYclDGjmVT
wlVLIpYXjpsfxD7h0aIhrDeVXstRicZdnLK6C0e+/BomYP9FGuOjZ1T9Jy2fLZP+
35DH23hFjhWDF4km60fqyrMjpT81AhcUKY4gcY2P5NEwAApMMxiff1aKZNxSmfC2
vvGKAUTUWpPpLKPAtTRo2NqbDtpIxOTbnnnFWiIMAR/wt2q/rHpN5Oo25EWc4GRL
2bXrQFXOmfiRXSd9tW/j1rzGjcUSmgor/opU+WP0nZmpnoDnGMf0Bs0143PDfjmN
YBz63NWaVwlRlzNYgYUMxxj0c4FLNMt/Ndt8Qi5D873lLqS2B+QGvK4whSAhh53f
uN7xgyAZukiPuogk5oXfx50VsIIjioJJU9txsiFZRU1u/865kJlMnErnEklHSXdu
QmtFaJ1Hk6sWT3nwp/efKdPL0MyYBhTULOvrjgg9TOJ4AAPs7+JMWRTDs0M+syUG
auBnP341/oiCFH2Zjkb1oaZ0JYQ6vIPjL/IWiilyK+s7kbVZ6eTFNFc/JqMwbiPz
m/PNTsDsvt3r5QwAd8U2BxlNCSbHDTPBG4t+icomLgqnRbY5L1ObmKa/5k48lfbj
GgC6uojTm+mm83DOi/N4VgrJmyKo+QL73hH1GFOVLxVW6RCtI1oPkLY9Y03l79U8
YsZ7NXZDDwd4yB9Vs2vv6PV0G1It4c2RCnLmQYPM7iuGgdmgKfy9V9VYBEQG8Jzk
C6guE+rv2AMF7sRarbm70lZrvNxGM049xuhQjNucQqaaAQ8DhELcbDRLoEQKnwoA
jQpyqksfHv8/jIrqIBkL1CNCnFOdGjeuD/Gfz+ekmcqZpeCpxvdnmH4VZu0b+ELh
bye6LiywIOocpXXetjflqBYnDveZrKOWVlKZQf3+CC1w4P0LnPn76YsFx8YxltE4
qVEfzkDCYdnaddeMDx7KW1AuYA29YiDASVaqbkSWMFiql9myYFB8zCSIpOqJermZ
2Ku+0vowcIyuzhQLmpiMOPteznh7MdPRefYw9kgbJI4g/22tkC3wVdaB2YUO8EI4
Jsvy/Dos2u6D7MjhVA3y+AGfr9ZJ/fljXCbqnh/K0ASve47hV41Xs9JIUmjIrE8s
K2CoalRtlBuHJVyqJu9p8F36ADJxtLx2bu1Lt0scqhBttBWuD1Z747kKXPwnZIKl
kplCBsblMJH/DShddVnxPfXQGkmXoRBqK9eIpnkMiPTdAuYj6xBaPF2UWLTSVF1e
Lag2+/cWHDbYqMMkxlyctczJgfr1hsyGth138yicYW5Eo5Hx76Bh9qvP2qd6nH0p
WMn1JlEvT792RYYbpiNZyGmDGhwCSgsQQvki695RPmK7KkWKbnuQhOG2IVwC330B
fXw/RI9tk2BFXJpSBsn71yKkNg5kU7cjdNPwE9SV/C1wPAQ3qHd3kEoDTM+7ZUw3
nX8Q73FWkPSNrwTJs2ZeO6QdCQi+XgNDubmb016viedhbJxfjzJwACrV8yLvTS6p
BtYSoPgHccAv6sBRz/58zw9Wo189Qjrul2G1Bu59U5KhBlbi9XDEFr4AfWTu6WuC
YcUlX4oBa19NJ/x7/55pbPGuMFp2/FmNhKDnG3xHE/Wwb3TJTal+JQCVxeslfIq5
QOi7LGNXjhlw4mDlkXDmFYZmN4MCJCZfSq3oYd8gYKF3gr2HeQSDWqkx6VhBxsNe
aTmw8Hp552rkzBWdrnDWjgxPeB8v7GQ3a9/tYl8ZNGbXfcJBLZ5I5IGqH/pPDL3f
SPryNssmTJgNY18ys2nSHIx8wBBwkrtfPpY/FyrONMJ6zMrvkwaVexfi4Mg4PcTh
JSgL1ODjaJKZu+uUl6QmqoIfMtlWkbYfhtvdCDXY0VnNb4Vjl7IbsLFL5W487WxG
zWMYjA/nMj6UNeyiNMnLy5KTYXZ8dgnp0uI6PPSjHjcNq8Bnr4FmtZHZWfaexcG/
dCJktQC5u6hKCUtGz7+4XzLx4kF5V2bRuzCWcMKAtLCONVKNvxGTbDE3bCyMvb6W
cLca/qgAsI1LJhUimj4Aq5gFdTzsFZWTHR6r3OKkPQLRj5g1HSwwzhYaJKjyulP+
WJNij4yHEATh9nqlVZ401Ub2WKmv3BK1NZgvKy/e7AbWYhjjGasdnA+7nF55o2iX
Tet7qLVmMcy/73ta+ML6YsY52Hdd0mUoYPmP5lmYlcl0IygQ8qQcMyFLf+Y0gsd3
3xxdKA2ECzcZ1exKRETN9cC+a9HMg4SDDWpEvfLuyQzy35v7U44ruL5Kc3ZgFQNG
Dql1U2twdHu0YYkoWKW2vKulnjfzscKUqDYBPHCgvBU6s274rCd8DkClMmxzdPjH
vldtWgGlNx9nJneMAY/HnD1Ssy+RfEGEEzbkkfXzjFgthFvh1k3sFWTzisR8GrvT
/T/dfSv2bzLdcDOrQ7mrycJ3sg5oyphPdSg111fCYaYbWjittSEldhr4IJZhKFXG
V8iP5R1CJAuQXT+uaJmf9yIxGkZgZeRw4TOHbg9hEfjgBO9dWiYv1A3rn9SJhoSJ
Ygla9SaXTFGGOCQ89uWvdJ5P949VII+ZmF1hDAzbuvo1QMVb4Q3m4MbDUAv4LUGn
xJFJkdHEfU24U8+E/SgeBt63yAcGlJytqcwATtIuHCkqAOqaB5U8RBlGZDI/LH8Q
NTmEcLksgsvMZKHKY6uY0iZ1FXf+HvkuTFVI1oGt6gz1f5Ue0LbDfQmbbulEFZmw
rR7V9RQIVDaHs1zGYdR0C7ekexmci88LwAd4dYbB/jDsuiB6sMnXye/OiyeCLHEl
luLrchdWiXQKXRw5Jwow29BTEBBSm8ESS3FJ6JrYY2dxYrQGJMDcsTiPkJa1db5l
5oa6e3XyweVwrW5xpYvdinXBilSEJJMaVR8lswDoE6PdDl2x80IIIZ6uyPSWC2Uc
VqDGuDIaZrMyZ3E/twDLxWBhZuCISwqFQAtJ2Ow/45NR6tvDraabLxRkTzSdEjI4
8aehuYL2QdTHgX/3GX3scAQyoT97wO/+IFT9D6EuzLcQmhxGxomO1zv/sCAgVQ+3
F59CTJL85hgULm26YTHYXufgmwWhuRCj6qHe6Q0g1BZVDhak4fc9fRS/LD6osEU3
3LYICGyzSbDBWi6Ll9jTGtUP6RI7ImvCR3XZsY+lAPG6eNcqlquVbIspbqfRqiSP
0cf5Q69yj8j7EwOmYAEszRb2/D8ySPwxJRXaOfxf0Ul5wIvaDsNZnCG59tQRNgYJ
QEFFTNdT/EIyaXBy2XlMkoNT6Hn1iaOpiFQpQFEv5mGQ92rGRTxvboblFKHNW8Jo
pTvL/jw4mqOMFDqKDKsDr9e7br3gfVRnyfZ71/UabfDgWWdtxa2sIjyfyYzo36yr
83wyC+JLQtp/NgnbOBeMZGXHe/1vTxkibz8ylwqroPmvDFw22t7tu7vFF6xXyR7Z
VknpZCyedm2fhdrIqjDVqpKg/63sVAm5AM9laKFaRO6OMRi1vOqZX6+ak2iuvLnp
D6HvqkW1Ixbwupkr5t1cLByhzTGa8ga0dUkPXA/gzK9i+kAOPxaCBgOvRLYXvJUF
Yltk0hKpZQM0HeeWmNWk/0zmm3uSKK4bansl6Qab5u21NSn9BmwhyBm9EoIUSXmt
1U1LWfCy7uAcZci9CY0xmrRnALJL4ISFrI/5Oal/eY4u+taczaQhUe3+xvjbCehL
QR1bVyLYf1q5REJmYvzP0DMIG3grRyNT7VDN2sExINiHkFNAgmLRW3UTqFJsvOET
UsR489mJShtU5mzz1e3cci73zw0/UO0JozqImCa6Jun+ArWcVaq3rl9nMZ+7o8wr
lJakAtVpfa3LbvR6+gheEowndv/YYr00gSIE0oGWOQo0IurJK7xPG2VUaMNIpxvd
NrCvIxQsi6n9OAKgno8S2aTsMclSn2Li+Gw6FCqiNW8tK8issRGlAMu1Rx9X3Bev
jzuc9cUThxh66XuRjs3ZlDrlnDP4hBc/699AzLVpSzz1G2GrBDiydbP25BZh1HiT
1ZKfs/Qt+7nRFbTwWvmgJ80aQbSa73Ka/smIp0VFDiwICfnZY+sSB2a8RYfdiNij
WiWhKXNEpsFE4Qqe6rRkAW869n58ByABHoyr7ChiO7z/sHqfFBL8Qtz/d9xDwulL
aC5v/q/9tqeMJJ4TxboyvpvwxqcuUKQpF/JAsOgxfy4zAbOF7YDMi/Ggnk+zo+uV
TRc8YcCheHch8m3nvvXZ7yb3Ncnwu4HCw9pTwdEr+410yTMas+s+d+9UERC6x2gj
2B56cPtCmrXUVYkeOPTjD+2VxKpi6gnzgV8h3UI/4V13PI/eSyWTmXsds4GhcAxx
YJPcuk+bbNDfdi5Yul9bemYudiDSQ1gHcVJIiHyMUNcNA7zSMMJaVhwsmKN1wqV0
yzTLOTA3dNpJ8OhL55tdQ1CmR0V+QrJK1PiYZN5BkcpW/0YkHFzKwumUI/y1ClT9
kSDC1WkGU46TYp/lcflZfFs48ppLeMT60oMfgo7N1gnEEsTwPAOV6UGv9qdBH1gS
X20I8Xct/+3FLyhTCQ4SsIp02v8k3p9EXPdliK5LpkJHNOc3ke57arwbEhBXdjPw
rZdZfiT/PwU1IiHFASSiJ27PJLjZrz5nHuhBKX1gm/Kohs2mLacSSasnF9PPLpdH
Q1wfz1B9zFr2oz4RZfknv3bsjZJscorZAgPQOd5pVnP6HE+AlM+yZWHwUZDY7cCn
ZkDdXXn5L/DuMkUZ7hR7wvv3olCxATy0e94fJiJsG7Lx1d2ObYd3yJOckvp87jvH
nHfHYwu32wHLE8Ch4w3jYXYXU7qmVd0IMIwhfdSI0UvugTH7DZgog01e1A//+0EZ
1u39D/FBRlnf9Ty+JZim5bVI/Btp7rz2ei36EmCFesTBbxjaUkikiqTfpNTHWcA/
5AOG6qjFCeHY5Ffumf+1Phr73m8wC641xYmiZKqV65QE8Uaw0OTULrg3dMYRqSwk
z94jN875lTdiysxGo8p4bYHbxPEl/Nvivz7CXF915pR2T/Hnt/IgeKCLSiqmmsqx
rzqn+pMQUuFyidLguHSI/dXiUScNx8SISl32V6jRBYDKMqIjzetYh0OENWHDzw2S
BYcceaCynN7QGHnnY5DFncMS2QjEjMD3C3w7pqx1bJ2+JQUfDfLWggqK2phoa2ks
6N4AVTq2vyAsA+eSfL468MxAU0FlLgzrrCh7WNXP7bZ2P9GSnI0zIPk1QJvRtVBp
Alg3bvtduOL+FTXHv8NdU/g+7wddz1g6cJR1ZK75aE1GQaIo5xLe+3NzkplkGmj5
2HNmItlRwHF47EO54juv37hBZDdub2cctnNSq005SuBhk5s1ccKGB8p3C1HKyji5
2sVVSIyM4W1R6rMVkfGp2b08nEmA1SfrQ3f780LWIvzrJ012sHuOf5nXDYXxA2/L
BT9BYlt0HJ5+OCEK8SiPqecOysctwzR7bSNz+mkOueE7DhERrhpCvc2Uj/pPdeFo
BMxO4X3nH+Tbm+c8HihC1a9VAiAkbWjts+u96DVpbD8n5/zkferKE/mMk/oBMySs
+l8n/7WNxtsl7JYyQG+erLFNbwsHvD6m2x8ic7xzKB9qU+H5L8eFDOQb5EV6+VVT
cY4CawFBU1rtu86sMYD+ugw9SE9Ax83P+2lwUPSQolofHY+jA1X6UnNpIAgQFf3L
B/PLQL+rxe4+ksAM9LU9LqiUutQiLCRf5CkJBKcHu32/+h46JmhhBZKlQbnSeaKT
ELdYeqObfwm3hoOARdEKsiX1hHA3vsS0PLLJyEqxa3fvTl5slnXh9lc26RtpV7/e
GoAFfwOV4CvcTbK3Rrn4KYYo8DJJlG+Q2lr6lbQ7fxEPvbry9qkRjBuAohPRqRhq
/go9FCZOIFL+wCOnNGUy1O5/1V6cI8Nd8VeSsuxNRsRI27cuqPUuyv/FtmhVz4Cn
6/m8Mm19J70kjv9aXZbX0I4cCG0oQCrxuI+f3bqQ0L9oVwU7A/EVavwNqqYN0bP2
zXNce83h7dTzsYPa2YIpCjiKnU3fJcgphbsGqCrDAv6sWRy8grSIag4dOoCeFXia
SfL9BpLMKf3id1byQuzvZ+ph/KAulLak/JQwnrWIcx67SrZrdvl5D0AOuZX1j4l7
R+5MYgvGkGqzsqUDFVb5YxB5yJgEVimcOytRd+/yanS+k6xjuDWTqdzxw5r4WpLX
xDSY1i4+VIZE7OiZIuZQTm/FStkxn6v0ax3U//C2kIJ1WlNQOlmGT2D+TaWjQUro
K5BRSmiFumVEx/KiRFMX1sNtJa6igiNcHatWR6J+MlfSmrQD5ZZMZCs8Unw+DTq9
Kl67zHELAbussRnNI6tCnB5oK33HTONzzF8ttCONZ8F8Dzv+ZOP1qTZsypiNWMOd
4MspkYvbIuIXx59kDQWb+PVTfQIetorzmBvFpxnK5DJfi74E5lyEQEnL4DcNLsEY
PXYzSA7g4wMYsWJW3u2b4q7HX9vSXlKSnii+78pkJKJFyKKE9oarmVT37h+DHGvU
eHm6DJfxJIcDQJ3fil16Q8HaGKavqZqA6NiBPLbiI4bsH4LOde2ZQW1s8YvW+kj1
ZQVAJD6ZqGha/Os3m+BBwSRmaEMITEcUL8ek+JwWtPyOV4ef5+nU+0tdCK8UBYbn
YZebykX2VcrlfcB3I+z3wuD3c+C+I7VZSBfZizoEDhPuXZHrQb0P5zBvFlXGVSJL
yjvHtvpfSwTjq1gXJLdI1Rx/q2U7YN/MM3DXP6xcdveHiUjAmkuCnv69AAHupBJX
dTdedR4U5U9iJ9Tukot/0ED7w5MnqdJTr2QrArU/drWIikCnps/4WVAYk23TaFcq
dYgWzzCEVGJn9ExlBog5s867rO+g9cAjxwHZVSW9bRIzrVMXPCUE35+09dPrs2nr
Pd13bNcKNoqHOXl6D8G+lzEao43FTx3D0f5PDGgwlSgiltPJ25DYNmUySXWnqUk8
AY9KeFIzfYwTqAjkkb8sMwJPbRWQQpo88FoXop7YCA7uwx+igcnrp6k5tpfY8gQj
proSaBSyEDAalw30fyp6fPpSwZsBoGhBEqjtewIa5vb0Oi0Epx5QEa2txTL7MheT
taLSWA3wPy8w9HhHgFgxeC8QtazT8zOBuvzQ4+9zDrbHYWa1I0qqUVhKvY3ULpy8
pDkk6C8KQOIcxbs2rMdj14gYKuWZ+YRohYScaIUuXVg3xtEJMDyy9e/k4oTRlqjZ
gla2pouf2t1Fi3cGug8WQOQ5LIFnbJ02fUsCd5jjLeKHmWMAq9Ewaw3XFruN6SsB
6HzF1asYg/VKsVc62u62iFLs3dLSng5Ju08nQ73zjAslHdb5ul2/r24h/FLx5TEM
VGr/QFJSI4EeDZzyPoZ4XEk6b3hyUwsfexDtNxAet5ADYhKfy1bWCsQGcjoeDTr+
xKuk2xvILpAZjwE7SEGtHEaG92vohz9jtGnouCLWgVzEKP+U4e5WPtR89sxMn98y
2UcXsLXWU1VDhtFNQbj30wdYKWgkszUEDEARgEPbFTJGxoo8WIBBUzsrvLdmnegW
MCSqb02Ar7mAoX5eZynysxLn3QpdGa+D5/jTLwTdv59m4XGn27pIPZV+bPtTFfwm
AW7PUP/1G17JgTUTSUjnC41+eumpeXQO4rlsv01MTxovjDGMvVBOxmx0SkIsmCyM
beedEDFBwsOqAPJoJbNuuvcf2YE5FNySn6ONdRsQXftk12j0rGtjjr4QYhuZvVEb
cCaxM9EzPgrgMLRNHk5Bq9Bsrj9W7FGmXtQOkoDKhZTuvVS73po2JhNLRiBwgArG
Q19Sk7jbAwFS8ienZKcFr7BF/CD6rAlYarn9sIci83g0p5nIbhh52h0VEtDzjf5T
nD381NEuwViX7r4g2/g9ptr+mYvwhNpIGVHjURE6+Cmk96JQtQf0/KAzVmMkP123
6o3s5PGMFepDdXbyd5m2z1R29P8OVeodEy+k0sq5kCHbHmwGVhjAxiXEwiWasZFX
UW0xzDrgzgdKoIHPXT4qHFDs2Qtlnl8HBBxrHkSIsmPR+QNFZv5Isk/mAlMptMiw
lBizH1MUxd2MJz5+SSELUcVqokeG542XOKVyyMG5SmaB88Wilw10OuaqNGFHsG6z
wr++XuePNWCPd6UnOt1w5daeXOZFXEH7IEZ0ERnIPnsRl2ssck7r9ADJQiYk5HrG
OJD1GV76qgT3L8FEXlfwS5pghY4zF4ZaP9DuM1HuLbUv+dbYYic5WB7owr5I4dSO
TCMYNO9hYyoABPMnxogDww14YnsQytzefci/1JgaaY1yYxfMAtxCUXv8SlnIFsbo
vpbvfkKSkFG+tNjcPcumJxNunzfIyKR9F4gXECx8cWkisHvGO9U0/2f7yWdU7pWk
5W4iB9vt2a5K4ioPYgPMNA7QSu0z6i2qxajp/pWvv7xWKz24pQAO94NvMi0/Yz9A
TdlaOpqvYFP7Fx9Ny5gJggIZlBBC6N624wwre9N9vDGu/sL2sU7I5R++MH7G9izJ
Hlx0ECzG/pF4QKv5Y/+3vOAzm9wBwMqGQNRnfe08VXMYZOoQQ8ExwafosM+tGFKO
LZdiW6Hdi1cUSRvTy34GN/85I9CLFG6xxxbak75a5oCf+NXcEx03+rgqhq6wtSZ7
iIFTIzdR2RDyiY4BFMzpHdRajfZqXOZO/E38VmmXtaOO+OvqXd/p+RSEOvR1uuvi
GhpHQaHvgtvNhH6hBHHcRxvvXUtOq/uA3Mh27srYuFACPk1wKw+oaajAt04sDAOP
0AHVS0sqdkJetbDe2pM876DdwVKsBY1H/4gGp0R1/0e6oOdr2N/7VD89hp+ppQCZ
h3WV6Eqo5kUujWeF9yFfeBOwbH2Kycs+peenA7VjR36yZo3NqNPFN5N//TDfDJjp
k7Jgrx6nbE2BsA8YzFgFLdQkQHxa46zwAGQYwgJfK+JtrV97IEOh0TSQ0e6JnwDf
J8cyoMLLkJ4kaPjL2H3ErgmXuhz2AK1/fuYi1VmhJDglwOmdq2C1bcYO/YGNe/Fh
8tXE112fXbzNcf/bCwyOWeE8tSxdz/OLu+F1efRh7GE4pSkdK5BjNjcgyzJDkEd4
qEDsaqHw83I8I0MteJ8pw5C+PivQUGWX95RkUnGFL1UC0gvefZUxlxe0p/qYqShA
jfwPf1kPNRj1X4kktbLIREJQp30FcHt7uIARF/Y6HiOZLwzKVu/WJr7kY3EbQ9K9
qDfXcE4XPkEhsvR9gyZoGBv0POLyJ+PQS1i71mGTaMjfVOa8L0yyIg9/Yg9s3jqF
ndoNV1m8v4ZdA7Hn0upcojGPTOdUfAnrRCCDs1avBQZhFvZs/Iv9nmU1dLUgrnKn
SyDES3mj5SiXwz48MzAvYs1ZeIDbV6eVrcCuGwOnaaerEMS7cqtAndFU7lKLLaNy
Pk77rFhoYwzQaQ/e7JUu3g+gPr9TmvoZjT644YtxDe0Ec2S1gFaLksHNHvpC5Uni
aPbGIj81DTFGx3n7BwB6p6PVvgumkj0BlfaAcUcFj5A0rsXsptCrdDDCdl/qiw3S
cYNFlH8Xww4DiTM2jyOnQ0AfP+cErUrfo5gC3fatX0v37ZrKP9DRtTDZMs0HSB4D
H/6F+uB3BPbAf/lg9RdvaGy6EjlmDB/o/CyuEwbW8a18uLN4PPu244Zam3RsBM5D
3ekcG6FD9iRx5YVp9nvPO7fZ89kE006Tl5su9eeVno9O70S7HDn/sgc+G7L5cwXX
W/dkLSr4qqb5d1Oq3uuGHSUEPd5N+VLIke1fj/4ktXJ7Dn5O4O8EPtRZBDtVL3tQ
XQgTYn0p2E0sVVos9mYMhVuc8cOTRNLWLkOCFWtyulZDHtwP567wQUwlny4q4pSF
yjUvNYMYcIBoAMRr/jMSdoGF7gr1mmn41lwSC6GXnFu5OL+k5HZ8FBdJdCiVKsJ7
H/k9TYRamCGFxCta/4ODHC8Ajv9UA3NlE/PU9orQ77vFPG2BKONx+C9Ip32/2hfH
VTXinV8kWFxWNN25M3OMpmVfalNOozJ7deJV+H2MTDetTgI0T35ZNOpnlwIrYTT9
Gnd2dXM8jZfLnSUS0gyqsPnCsCWX2GFyPRzV5BcRnEC2RoMVtRNcL9aDC8Hp8Rb7
yDRrN8eaSYwvMQ1ofiJS+JR8sr7KUH92j9ixLP4CuU5eJ9M2gpEimeljNxkZEfaS
tPd9BSKY9LrOrtbBeUuP1qrmUZ0WJWnjSlKqyuxiP3Oky39Y2moPZvhm8wfE76mr
V1MgNtHaP2xMqMNHUPRn4Loh/crUpcTZVeOu6p85mEEG3NnBRSYX4X0WsmIgImJD
+9KT77kTOdaueVSM0xrlV6C1zmsi/MnwHcy2cmj9KHj6zlL+UNSXxpMsfhd++YsY
E14JsFvstC9WsIGBWANvamCEOhgu2d8Qbo+T1GdIP+85+vCbVpSifUWGIB3gUqxY
/YCDKUgPXnF4NRYJhpM4gMBwtZOQBYIJurfFN75XkK8yqmiRQOHDC/3+Zlq+IYYK
Dn19T+bAxdqB1JaLJCkkgiEydZ2b9ei1wR/lFkyem3A73MCEc/ysiZFxY5/teBdt
BgRFLv7dMsEm2AtXt61O+SNZgiWpG4AAVfbLglTyzC49E7UIh6/0kvwiYgw+cLRN
Z9WaVL7GzPLUlGrypTniv7Xn6KM4pMUGKFbGiYAFK3+aG6nddAjpJByJ8q16rV2I
Zf4fgOC5i0Ca95tbzFYDPbLrRa9gt+2zcl6QAnkB1P7M56lRV4HD2+dYhTrW8uW0
Ws1mDx0AgJht2ecECDi/A2nWss2qo0wdDzfUjKhZPYpRrJ5zn0YWkRBFcQAgWw21
9Uw70ZTpOVbdDlC3ryprkDaNQ6VQC8r1a1fbmPLhIla42znyM178/uofUV23DqLq
AxRLdM7VTUvdNoZUfWmPMiEaPy/+obiH9ewtKpE1G7WluWlAlnnGFpSgqZnQhnIP
TG+2fy8xXMLu8V/j7XYiwK8iWBheFs85xRvrp8vJRtGuaWJqisjMA6X2xt6tRtPI
mBY1ZAYOXUlhEKgrt0KlLQCZaVnr4NYiv7cwWeJaR85CvaY5J74YD/KbylQ6WlCq
0PjJbKgiLBTU2X9lXb2UqOB/8lcxq5/2FmIvUQLQj7Urlvu9ACfv6F3YfxB0jBzD
UCSex+QR4/MZLhc2nrJ1+6ig82b6T3Phtw1l1OGJgqORMEeXBgG6QONHgLkH1mXL
OSXOsvkm+5duq8H74sancadKtJhi839QLw/UVm581p3S1v8GlsDM9U/6hWh1ABHi
DcFKhdeUpgnztRTbyckUqTsRsr1KAeF3hY8yiH8RxiOTosFfrZoUMIBlxtjYVGUk
8zeQYGL8+SubEYSJWiL7U1FdbIu1pgrM72PcAyn2T/0ZPYO8urvhhyXYLvJ2CFwc
rQsJMyG3S2irVlt3nLQoNN+Cs9Bp5lQ43vs+9lxvTPWoV9A0Kog649vDPxgfsAHr
04Wr0P3Fd4Nvq/VJ/8WOgsY3p2iYAP/GTjv+utQm7SQvWZ4iYYN3VT1h27s51+e0
tTs6kT7qQae9tUrnP1XQhr/eqjhTLehbJFz1vj7USacoXbtXuPZJgmXkWt978NEC
BUU5UXulp1KnOGpQegWqDCPwpnuyifddmG4S2f5+f/S7KWjkd2Tfc5nSL1k/ga+2
cjkgzUX1lEGjVxWmz6fu06q3GpRYJKNvLyavAH0pXPJDJzrT5034X44s+7lerzUX
3crpbRn4MQwVI4KpImK0L5XyVT73HwqOpVqE2NQ0gbsSgmJleRwcwTCIgF72/Jfg
8wHUpTUR9SWEw/k29sjpDelciBdPJ8kzRdamaJD1f4anQeZFMVyD35X4vrQqWCfI
HFL4Gwb+MrREyrE+b1UZ2vIKlqkm8sNtvcBAErD/1z1hGgVGObqcrzWPVbgqGcud
Lj3O0BX2bdSMDxrl/PePQh1kUSeYWAykdBa65cXQBSMESrORmVw7SGNTl91ga6QB
NgjVydUYd0bo/5jp6M28vqr07VLrs71RXSQBdmE+gs+TWlld6oZ3mcuH6GKbiwfX
qsZjbuGxDf87qdTW6t9gStO22gtW+ZVc+kgxb7aGnhetdg/v9H+dWAYDnY34HY2A
DANBdL2PV4NKbW9YiC1K+D5SNZ1ytF2BP3gzLbQ4VtoSffigRGMp/YAH5wcquD0A
XNAzmfw+p0vnyUupGQv81feNLByJLq6Un5Y66mFYqqhzSQQmLdZhMgi/47I54S7c
GCA4zFcAw/6AVosIySvu0oschZK13ne2YVArRgvtqUMDJ5PqkgrnqcdwgkAZuKyK
PAzJvntDdfz8/rzkukY3Ie1Zi1bWZsfz3AVPwqPkRKSurSvCedOJU5ln5IR46/QL
kYDCSkKKA5KnY1vP3NRgiyiSNLSpVDmCe5+mnpk/zfvrvD2bZ9wev4o0qP/F6wH9
9cHTTlZpO/s1DJBNpz1H3Dnl3zJJQZEBhvu0MSAyHzOxGFi8VumkBvzJFHt8dr/g
Os8wsHr3pm90a9JI0HMG0DvTad/KuAi3Rj7XPUwiC/VAogssEqWt15ZXJ4ghXA4u
Z334OuPrjDf0gF8tMOP3BdE2FjJv5GOFDtzP5s3Rajr8W0WxrTldav2nZex9E1un
V9AcZwxVk8UmRALZMYOQqf/COHUBTX2FpyN9j3NYSbBaxiz7YseqVz0Ny/hun49s
1JYYvNQj7GGwTvjKO09j1it7eGOaRSNnCRMNaKWeSb8peKMlgW3ju3YJkvDGmL43
H0iuhSshOXQEa9pxZZy/F3h84XQgP/nBDTCP9LNtnRZb/HgzKwTan6nncAIt0sxi
0gvJb8veX67u2GkmT+aGFGnPDYgJIt7qovm3id4jaMat7XPkOhlYM7rw4vgak08O
I0seVjDOQXK3mdmy0y2k2LtRq+smgoiq7vPj7+AKYRx+Yb+Eiipto0Yxosn9FYHV
IRYu1YASg5Q71QkqSBvQ73I28ihgn9yXjfLDrWsVYO+cKZTUU+hCw6cezhGNhK+M
v9a32QxYEXvLed7RK29adar+WnBoEzRPjpVvQ2w/NUrWBzrLvF6U1HZNLiZc8Q0M
rb2wouocZt6ZMOJ0vNM71GKnjwl/YHHf5r2rjwLnTvxovoO+t9wLCvyffkc/tzBN
R+Urhy2/BvmzKOG1h5dF4kLalhrqTwhGh/1K2lb3LTDMUpk2eSg46qNTS/3mbUXh
u6fm6mB4XlDP2x8Qwm1UgcHrTJ6PJq59XqSIp/BoCYypq8io6M/QEpnMwpemevxy
qIWaomXNwuF50jf1SwjSnSuZcPwVZcqr073skbr7o46UK1jA0W4ahCcUrk1yf6bS
oJTEeWbanBRAaAq4Q+orRe66RHPPaniddQNH95eye/pnkGDNSG3vXQPV/FDwLMg1
iItEL+9Z/GcLS795LVMo2onesluGKnflLEoOTIp2EXsH3XVdGDqEwN25vkUKybyZ
PtNWTe6LIOLChiRHJn/fLopbr+lUaipK3tkUZXP0eVtYpBLDMJ1XnJAa4zkjXPIK
EqsI62Tpk9bCcxIjLy9IrytmhiuWldLswP3mzl5bF0tGGZ0y9vNNASZqm7H8DfHo
G48jGTa8nhzm1Iq8xxTWGN04uq8f7iPDu+wRPvMVb2zPUIAENU/zXXuPIS9RNkDv
JrtZW8zbRes0jDVQ2fCG4jUfpKUCqQybc96h4wdI8WFscwecsLg1O4bPwQOZ7A/e
eIqjmun/+k90sFCLVoR2QyWucrPNorQS0qOjh9a+wui4Gd0TB2biU6VMqbvJVIaK
1I/gs1b86dNsW2whKTUgZvubUXfYkGhEzygP6D7BxUEtX4ZtdwHlCp71UPlyZf3Q
2mV3ZAf5xj8UgWwneeq2SZEjIM833aMJegqXIhZhDAwMcrlKaGwCX0maFLr+e9Ke
aFWc6NduZnTe2sNxyenuoEQSTsyT+YffiBQilYnwVRIM1vCGz+cObkElvGBf60uU
uBuepl24nlmv/qgeLNKbzpHLbUzFK1PBZ7jK36HUhprozlTuW/M6ObSrbK8WNYv4
HKfM23nOUfQAPp00VBXBhLGBISegEzGyDJEraxXVaQG8U/SbIZ2Y4f9TIc74JI2G
HRbPAFemBPV+HrK3H7sUymJCwgcE7GV3/C+JfB95YTFxkrnwSV1Q9m1O4QCQUiD4
DJ6tpK6vnQLnOzUvhBrjuSoEl3BsWJ9/jbIKkRKs6eIcBNpMCXjRVhpw8ZFKP0bd
4XUqPkalU+A/3wH6tA3bHvK9OZ4LYQC8e6eywkN5mhyADAXMoMRanReGzQgWT3Wl
HC0JVF6+sVHPfQWSHWHsG0uNEjrhiPj47oTFPrm5Zbc/Qg0qL804Q9dRGh1ZEmbq
dOmuM0lvWM6UlGzxVSRoQAcgh/UGd1wHykFh0mGlBwPXqlms7iwBms53kK+cBhFj
ztJH7YeeGvQuepHP2ss4un+HrP6ODRH/Wa3oMwBbvV2IkR0WpagTyG3dWMv4iPMK
mXExnCUP+ZBvXz4KFEriz9+1RS1YpnuVvbtz9mUAF+97Gv8+6c9a2pep+OQVwjMW
8k8WLLdLJZWOW7/6lZDbSQ03ElBfvMAPdaAOpfAjtRQwc3XanQGAonLSnRA2ozfG
fg3yGuupVQheITKldbRG0p+Wu+yR3/MPF/gUQnQZKwp4oRGZnoNEZwB0kQCZSvot
67jaX8DT3nMdZ9RiVKwz2Z5KFMglw34Gpk5RiH8bKftVTzVSKXHN9+173v54YpGh
4ZUBwXrTNTvrEm+Ar+6jr8bVseAoEDlmWvnqkmoKMC3pqk/ubio0YxXWDQ1S2Mw0
GZ7PVnyv6xlKrpyePErqCEhMrPb/Me4Bg7b6+dG14nCVkKchhEe1gRAMJAPi1G4N
cjD24aQ5NTsR2vbQ/mMHhap6OaEcie8Mq96tijnubhqU1dPiydydty7zUk2qL/ZN
Lana41oB78xOdxOe1ULBwWeeD5Q7zWrmGCtpwNn5WYonG9hZuRZQPMIoOlTb1o9v
+nUljzke9pjp3V6Nxv7FJjToTDNVzES8UJq5BmgLnjavAArxZ88SRWsxqCThxrke
A/NpwvefZZJa1aquVdXkbtVd6b5HRf2+iSqjPOnfb3T07AhHI6kqSuyTJJfjiN28
KJW/ZYQ+gI4rrFegb3astR4HjGEQygq2YKN4GpKiAcuH9dsfmiSNxBBdJ0WvQivZ
iXeG3K5aZMH275hQ54YSbFrEiCf1wtAHtASoKAAhwK8KNpSZ8D4aJkUWHkJ8shS0
/QMmRjCRqsUDfL7KTPGd3K7z+rhxO/sEp6MUMeksa5j3Cs1Eg64DYxdSCn0rgQT9
AmpID+IRZHaFlh4E7PuyJmzXdXX4ba/Cc2CNS5ZY6I/Akdek6NS6PVh4TQgImgPa
g+YhY8TUFlSjpFrcUYYd98w7J2rtuyVDaU2YbEte0f5wm3/c+KpUzjhAjUfC+RP6
fUTZsUD+SOM22UI5eh4PRcVzh+8nUYZUkEbsuddNxSILMyI+WSd9IWR8+qqKX/oB
ytyhhhofZMBSzyFHsB7UeBHzy0LxPPaMA0vwjlLY1E7YLvhH8rVG6IrIFSXbw0XA
r3E1htAUYnQs16AA1uqlpBc97iqUs88bwUHwj/qjeRPPLIDF5t52vHkysTDlDyt3
oK1Soy97gherDs4znGd45iSf9qLYGQr0Uyl6/dNKFRnHb0IGh9EMEbkhiprXmiql
ZLeLov4TeStvfsar1kpE3jma2R22FqImml3DRddhGD9f9WWFqwLYB2UlBpF5xV++
NckqTozIIoZlGNWUJ6aqvaMeQlMPvilyfERUb4RpJCVRvISiPkFKRwF4oh+D56Ek
pkAe94WncmT+SpFCR5zXmktF+6HtPbbfrG4gkQo49CVjOktuV3KaEbu46kHwiFyS
p7Gb0f2QJOAS7IfHGlXDCKBx3guT+yT1/yU/tnI3yy9pBYbCup+a7ByDbt08RzOj
cZtTpKZlq7C/FnI8yZ3KeNPnFVmK7ciRAkhRnD6TXvfCAHMTuP7VDm0APDaKK8zz
VjKYhPbB363E+Fw0F6C0F6v9zdSmCO6ejznD1D4TImRQbBevKGbMV3ZGdbyKB8Fq
jjbOKtODYCZfBqkNdO/+BWDYoMw9cXkfHXyOFheMwRtTjrCK/kVRX82yrINQlGnb
YRwMrSnJAXapympfOxg9TzCHZSFgb5c2mUbYC2CreVA8Ox7kUc22mQGDChIjj8/W
OdJRNaj1GEwaL55FygC2u888YMbeu0AKJEA6Myqg8xfp1t3dbYMGr9Vte3JIvEmD
NUH9owQQ1eYg7sM53fBMr7tig2OeYcdRWg70Vkz3EW1lcIC+ticY9E3uT5emQhQp
2LtTKZ/Gbn8ojBg2zGOy48WKxVThZvTyJDCn5WJWfo+GJQCFKiX+QpbAiLkDuY1j
lFCpKD6k2hpCybpTB0acmKgXRNBaR2KZAKiOHQpU/ebF7u5UHPOa9JOVp6EotDl5
Mh44OehTpMcKVUxAhs9tWoCH3KDZXmibGZkHzuF3Sq/v/91H3GkXbGu2ZF/ljdB6
+yJwGVcOEKiIV3D07iBRlvOiMA5PKpldPLxJAAIIzXbBH14ER/XEkm8v8VcBNs/Z
r1prtjAmB175PPJhns9kt4FREzZwPPRYuJwztYYZS0JImV+uke2O2IiEwplF4A7H
EHYXLdqQ/xL8g1PiTpN3oUg0dhoGfvIHN6J6LZzJKz74qVxRLjgjkx4CIpYIog6C
V7x4gXO17tfgMgT8dYOhbyqRU0m4wTd8zNnuQTSPFXyQI5fYana6mPYL5/HXVJlt
XK3tRekcHM3wTUYtFRb3NBbPpfY6226N4cjLjorktMjmeLgtdBh2m9Hx1yAPTtiW
BmdDZNDTLwpEomPqB6dt8Gjj1wwyK+/Ko7OFIOwbyNXbjZ2nPwEHjKNxs23h7VIV
KM2VSqob3BGrSvbi5DMuGJ13BEPfqMYNf2otb/VRtRYrLCOCe22I0iF00OnO0/Tf
pfgjrSPjLjgiXnEScNmsraK6F/9D5wjj2JBF9SmWCo+SsL1ngjzqLQsg0y24Pw65
gifRWhOwY/eluVUY55pY5Q41sCPxECORMC7c9MNFD4i9QwYtIiSYc8lTdgRM0rwo
7o45oQed53dYtytc4lJXStfudBQ96F0pbqbBr97z+x+OKAIe5nl0mkO+7sQmvx6D
mKfZhTVKnr3ZVXUQC4i5pHGbpcpjQRtHd8BWbkN6F76+wjnQG9qdVSH6CxNEcfZV
IeA0qcNfAS4b7RxtYpLy9FGboJo9hNhArs3bN+WXcxQDWEoYVZwf3be8zJiBoJYc
sEixxlsin58FCbAN2ZTuYkFMpn7JRamaArV5A8uqWBP8oCOVs50TqXp5btc5MQQp
KIpYr0P/BbGHhy57CgkeuV8+mRLEUrrXFrqbdK0NVSMOemBNNfp5iG6b6nKr3ExU
vqXOa741C2Hfb3itU17DpC6aLVXC4G1rv4MgtX7osDArS5VarTJ3NW7nKF7Zn6+X
okC0v1/5t9nQyB/Mjjh+lKHrOYDljlhD6LSWTrVPCUPZVcDRWg9eDP3H4eLqRDZe
1KjtitzS8/X1stGhLgabibKD1oSfy6pfo9jS95VjV4MV8yo1T8MRzCvZ/163ECt9
G5yqvOPzXf9iKjmDRlmckFGC2Rjf8EFjGgzzPJ/T8W2Rl5RmCCW+Prjn3eT0uKxa
h2rBC6Ki9u9YZMrteLl0Iz88o+5xRXg7WzahXbXbcxXCkjddGUmx5ncQ0+4R60VX
T3JiO/4WdhCukLnoo91+PizHt9hOh55ZDmShAPW2nlogDjUsSECpqbu5qwKDcisK
mcOeCxgPsrA7MLQla55BR1w2Pz5a7eNpcTsMKjgtG+rMBmpdBAGjQxT91pJc0GQX
U0Cx1ucFnJg/UXAgTs06CepdwcSfd3tkng+p5mBEi9uRiiuZdIHXk0nEmekBOcYN
Bn2RcYiHzgLnDmYl1jeqKvwx+g+fmLmhaDxNioSROu6/wH1bdLF2nllgaio6MMKT
q9E8seVWKXoGEr1pWb7jeWOY7uzkn2QEdJpGOh/ZZ89me4l1einexOcpiM+KXgBx
6n23+RW43o0F+ZN79Y4lS/gz6YQDUWTiGRKVvdbYAGr408mBwBdx+r93c7VRNpIY
a7l9vYZFSyb6VLWAG6QQTiXGVwnUmCfJMlxAbs5n78nnu/XzH2+49Cw4wSoP6pqZ
x9BO2b4B4ZyXRpdtI/khHkktUhdZnOIBW7fedGSDUKTyeFi4r1j0klHdAvdeoS0j
cTJNfMAgWtx1WXafujMSxfvxFip/o1cx4Fp0cPfdHwxZqmmb6nbh+uSMLQgdKZZE
JGVxsvMDqgxD4L6yX+gxCblWFfYT2cpeMXBpvrfg2FSIxU/zBSw45AFHX41L7B6K
8RkjzqSwdcEAexK9Ko2rU2lA4EtOqQnfUif7tsEhmdOk509CJ7xlgBtrMd2GWf/H
Fn9xQvqdrBFsZ+EJWEJ8y8mcrGSBqLdWt+1OvSuHeuFFzAKTPR4QyUBlkPw9WRM/
6VDlobBTmZa2MXcDDItFTygZX24FyBvOTdjywCfF5dmPRistdpGzRQKxkZlfAlrM
x+nvdCnXzyIo8G23hcTpzuS+OCGKyueozHv2RXx8HEj+mSTT5p3EDHis4H7oi8TZ
28ilPXZ6447s98HOVARvHVMmhjua78fPsKI7zdcxcEimKYhGte5njLGXadsdUjEK
VcxdvLux8Pmjw02tzWZC8RiTmwtZznpvZVN37YIYW91S+vOPE3zH3xuUhTmuU4ps
nUJ+E7ICubrGEhzzFVXVntG9Otfu8w72j+/m9kwOc/5Y16sX1zmxbZCjujqJMWuy
G0zxBvE2d3+3/BFZSn63HZhdbMGz3fKRoOx/QeTIaNvNStbysu9kpUUD6pstoElE
CKSXQYRznAoNEmYB+Ob8n68GkutOaMAQPdIcHJnq1Y+vBFHyJDwVED4ISmFitY6f
2nocl5wa/No+4D3K9C5NsUCttY2N6fVhGf3YHUGWHyaAnSwe5E1Kl8FIZpulCYD9
21aHGa2BnR/TlnDViG2M7G32SIFX562gy9HjOqvcBaN3shcUnp9c9dLxarKaG/B0
UUS2DjPM418Dcjv/ofYR7e2hqo9+tiuN6e5f3CMJ7iMYs3neVqvYP7MgcPqPLKJb
k4m2BwLmxaNoFtTD0kUi26v4glcJykIvthr6PSKL29mYFk2jeANORWcDdXfVNb5P
4Aj7JfavrcSj/I7E3R2ESVzcKjnv5ZC8zltv5vp/g5BD057Y0bGvnc4kzfccqr0U
Ah+B8tjrNmiT1e0kjHqasV3IyKJdR7oMdBlPLqKyVZAXZipL4mYhclSVjPS/lXPy
KAJ6isoRezIexmIorln9++XfcrpxdJzYhAEGcpRTGZtR0wcCBBq9Xgf7Oyezd4lj
sSCtflLspNtPmAt3TBWhulHD7dZXexqagb7TTKtH7gZyON3rSjtqYebEdR8vHlmB
27rAC3eallqPn5kZSgc68CP6dIr6TluAYziTMsAn9VajfGpoc/d6J7CBnlfn7spC
roivlpVfJRDRg8jYbKlMaHffmNzQXuX2zFxIQgxIKcz07unRbZcd6tEkhOB3Gh+e
1Bf1MgbtQ3VlknB5L9CIUHOkuwp6OA84PUmu9mkVt/eIsHh32x7yl7rVzr8D+cpP
9G0Ousl9ulJWnAup+8HMgkz//uwbF2IJqUJvSPY7JBRvrXlFDe0zKHI5WaUbJlPe
irypEyEsUtd0CXWT4mgXGBex8JUDUpGiThCaImlis7gIIFoGZB9aqD+bu5QYYRR3
BriNT7yEhjo2CdJrdBGdt5zMoh88HJGxNjLd175CHBxtkQUnL4ieE3D8lNOrH0aL
JdypEG6suQwchkrYjaJertQQ7I8X0RqVrgv+EexogkL5yMwM0OgSgacuucgIaQ5k
j7IR72TSIRvg9XqfzJpRySJmw9zQQ1Nqwr4CpVXGtuw6H/+l6sgTkEiyuDjnzdKs
bvdPdeVuiJNI8V2Et4bM05SMpin25j6Cj/UmWgSrt8vZoERYKWOMH36u0P9DmStH
WdoDyeR/P2zZyXsg1AB5yx6tUvUfs8LRGvNW7mIRJNjqsDd/vsbxxrbuuvvkk9HT
gNTljjMEU0yn8I+0Snu5LR6ZPExsdJTFDuCHT8E9eQbfP4fFmvRosZGELyYoIz+f
bJ8TLo2cL8wLzeuGeK5/izp+Ib0SFkOP/CLUkfCgrOB4Xrrx9N+8vuB5MI5DNQvl
Jq4Nez0HH0fgh9uA2prprk1IdXzqld7PccwcZQ95ZnpvMJkAwyN/FhjVuNW4a3V2
TMAUUJJdFZKGrhfMhF3o59Yj0yxAbLgJMmVnHkcCI1iZst801zLL8M7NyQrN+QeS
xCSOQ6SDZG7GHWCvLlIyAjuO2gNwImTT+YarLUUjFtmDHrw5r9qWdhnLkiEdtIm8
+YMVIc48gcRoQJz3wCk+3LX2evh5qCNsDYQrRzFMUzIvezW70Tt1Qaqmb+pxsRyZ
ftGOi17Jr/HuS0YLovNrNcOQJ46sLjt1bxT9bNOXkLnKS5lSQ7jqUoHpJzMFEYcG
xpENlUjm0U3nrg0uKAja+HTt3g/Fxhmee2oB+n0iLwbK4JXd2E/BXPGwHZvNpiUe
ZuvRseD63CrD2ycjh2cDkMnUYHNXoq5x2hIf4x0V05ax+RWMJnJievdWyc0eW2D1
nHGJKqkQLxn63DsCMiOvV72YXbHDoxYyGwwbBzOUoXGSJYTiHbsM1ZgcVWtIqceR
5UW/HWEKv4IqVqpUUULFP8YxQsuyIt0EtWvgHK/Or6CL8gsZJQVCgOIwhgZESUQF
vTxCnPLDyM7XkPfyvBVUgj4FhXSkS7IEQt1bpGGsKcBt7i3T4BloDzL0+zr+bnBD
I8OhB8evTH7jB8Mup/lWyZTtEl/rEnZsHsXbmpMzPU51DtMysu/N4akxiHsfIABm
AN0RXgsk8GrYCUTYdvkBfp6PRXDjS0iGPZ9eJlJ63HTKUIPobQeYo/4J+2WsjcW2
whoD2YjksaJIT4VmAvLUVA/nRnZe4qYqOT++8EMrfhB6VIp5DXoS4RyHGD7hMXG+
bZ9Cb6p55mUtfw2/lio3+fqQNyW/dJmm9BC0C33Sz6tmQwR/ylcLTBQk8A9uDUt/
JnFdlZDTa6WQwBY0fWMw89OPX/vtsJFe3jDmxGo1UWsAYSw2/K5ua03RQ/TPgV/K
EcFshZrZhQc0bU5cA8nQQn4Lcm//sKgEs9wr9CvUTcxRpGc/SKI6Upznfp/7yCzM
75Cd9FTZEfM24JG9In25hNEk0dmxoWbq7Fl1GFoxQnDWpmuNETOZa5U2otdCpp+t
4//gzdf3mZ5Clk4LJwRvtioR7P2wHdPaMnFJG0dy3+jdYtW70aNHB/FpxWPNC5iv
Ukqr6M8Dju4baDN/ZoxdRRYbYEo2G4O57LoSe1gxAxl70InfZlzsCavseM4i/xjc
G3/XAwYL1231YbzsAouS8VPBXT/mPobSjujtIrKD+QK6MUmPW3PxecpHOtjv6Yn8
PEhnuwosB0KqndXGal+spiaA/Kh4sI9XawcAwI9kjWnd7db+DIOfXg2Id5xV/iSr
x4XtPfmY+DpEFwUW6AXd1mR6insixUxZRZkdG5vrJ5yoOeUh0HNicomXy38gdQQb
+2tSy9MpCbA8ixWs6LflGbQ5A9aaH7fLkHrwOOSR/LGrYe4/qKpUJ9+0l9ajTaXj
Ep8HFyHfZco5oaOJApIl/awxrzaUmtIj75Ufb0555WZ+lQDWTsbnQ1I4+0k/i6Kt
AuabIEsFsHbtQgGfBnTSZtUhqPIaU04Hhy8m9DkJW2wmjPetMTzyIvRXsee8Z9aF
A7m3W+7AXsT3QGDu2r98hjFX20qPTQc4wwSWAjTYXSimHuYdHirjnmITnBWkg5Z4
3so2DFM/XgKFo/VR+zg1WY9pL7cqCo4qPdcLLgTXesESVh/ethjZUl3AuJgIDBd0
+SyP/DrGqHnuFI97zs9D7K+EjABvRLsRnOI9ZoncTl72I041y8eqTiIE4dGJPqp+
rHE7Az3F4uLMiH/qbAaJrwZcagkc8oIAiO8DG6ixh6XGjDXBzEl/sdjCo8sNqF58
fACPg868YEWxKcJ1diD53cdVYg9TR49PrvIaj8jmLlmTl/va0RFI/Cx9XdJQNnlq
i/ILM3GCGnzXvZRa44e28wX5/lt3mFSN7xTXTZ0fcUMI4TE/Wwwl+/MSpupIr9zs
eEfDm+rGy/UkqxVTdeUS1/RZVdo++4jcbF0LEVvvMkpKLQcS81TIqytD8mSaR3ZD
15pQ+HU0txKgvvtIhmgitorppPLPNxCeyGycHS4u14MAFSVOKQQIx+sKaQZViGSA
9u9ND7Mb+jNapAyUEQ2leHeRpXyDHndt8XQCRCtbUyCE1Q8pHlJqHw3PI0A/2t0Q
w+MrB/HUtY/XwItS6Yql0MyN+WF2DAA2BXF1MH1n3JGjFTJ5Erk0qWmVI5ZGf4xS
6xWzGLIKvWDskzRoxJIGUgjoaiCybNkL07mgLsSFnnrcuJ7NuFRF4h1h/huE/Bvh
dID0EyeOCGElSWmlh0xF4lh8aWVh6m8vYO4XQO6YhQBh9gh1Es9U3TSCbCKiBii1
sGstlCjp0UaLvisl6jrb6reNsRkxhjLVyAZd1prmS8BO/M1aBRUjTlFVqAxAvg6l
fDyH2rV62zhbzQIIlo8C4JYn7i0l8LmOhcwNYqhimfh5jhs0hlye+/wTOZucbOKr
Mu2pzYXwD8wQ6kzR3Z7geq0QKtxrkb8vCSq2LNCyQCGjtHF7x805Id4niHveQf7G
e1tP/aTK47NTNarORoQ87wyK1Ieq4PDiPyhRo6Uk8V/oVj32uBP0RMpWCIDwDznj
jzSiSFTkdfItONgE3f7YQ3h0PW60D+q6eSd4CySJkJigRnWJ4bB9rdLKx7C0pceT
rwBM7y80GcTTkhFyIFks4wrn5Te5O2/+6PCMT1SaxlghafmtxEA3Fxa8fXWSzjeL
7uRh25dyHc/ss1wI7+XU2gDki2j7l5k8Ygar6fsIsb7tQYTD5sJ4+QTAqDfRSxNq
VMPiB2iucqU29viJ6QeQjQQGTyD/xMP6Q7e9s2241Ctg4r8Ja2D23cxG2sAAmRCj
zWUJWcB5AHvS0A+17Lpj26426dSZCCLL96mVVeov68fbLr/sMcEow8QuyMeZf/pZ
HqpLABxv/SRJGqkVQRcj43SDdmtoll5HLfFb/dqD11uCbJeskzXi4xAQATJJyfq5
qYXrPXfkGExajZbmVv9/F4pZBjvm9lNF1igGfp9UgK7mIAYJ7hkIcWSvsq05CftP
n4QnQGXa/TniGAvzP/g6B4vH5t+uRM+rDjpEMySZm/2NkMzn+Wgb79WTrKGT4Bt8
3iB5igsT0F13BSNarJ8hKX7yMixRXsGaPbHORGSfVYjk2w7PXZPYmP7oYGC71KIi
r/JEyJnC1wrD1tfIcMm2B+oWwrM3WiuPWPF6X3w61zsIpi4qfih7qwRal3irWiEP
i0vp9eRRnpVDPQWcsJyPJFWwSBdj9thj8GhDCIiwRD8cG4ZdxDn7dwA12iz2ClDT
1D57oCQ++3YQ5ikU6/VDbTjsOCgJgh0+SqcvoLlHLiwvzerDB08In7COFKkog79B
VZXpCou8PLT/+xOdYLLhBxTanP3+4PvFR0Whgfm+eBRzHtVxHioCo9aMdD3jgIGz
Cg/0yUuANuSTE1FL++2xmnuvU0B32jBi4OddiCDdTPdhrjuCAjzZ0HnNDLs/B1UI
nao2p/3IVH/pLv2rmBAQQju/wuR+r2CHWdyx1khXPKzguO6CT+A0RcNxGSDhbiKi
K5LFzqSqJH+7S4aRYjDSTaIcKKmHnUS89DxGDpdLnuqmUlJgyDehF4718oU9SRVX
FRBdfckYlGVrm345adzJ/SrQgAJQrIzha1jX0kxMO/f9y9ffqU0B1OBlCNj28DaD
JB1BIbUd5Z1kHOXURbX1BqiofWWrsWcS2PuJX55l6JAx5UYZx1V6hJ1U8M5/4aZP
NcRs3amIn2GqrHz4svBnaBKMukNhNnK7eq2UgcQJpRp0SsBDquG20zjD0/Q7M3tR
xLnx0twDHYfGGqFbEDevySvW7Cwsvk0u6N6tZmj8hZXq0cWq3Dz98kK2RZ1lgNXw
8PnBqhkZZmXrU9spJIWJGeieaiUnPHq2rLh5GckgKd6ZVDjePj+68HeQfekPA7ev
cUJRqKfj1jwolZ/mrB7IHtFt5EmKEwbuikSXBuc+fTPtu96/xGuXefE+qTsQK3LJ
KjRcl0gDZTfGQ3J1g8w6MjrRJyCvJTLHbPrjxh2doX1zpaOAOK69XEFmwiMryMlp
14xjDOz5ibENqkVBzIPLR2zUwwIfTACNpxtSo1BdW3Dd5TDKQuuozmp9e18cFFNK
6GyCMMmifw2iqN4kj/Vb9Vw5ZGXYXfKsHd9WScxxr+4ipxRTuLtBE+UxUSUjlLxU
38B0L7MTAiwN2xKD9vWssoBUkJp8/kG9w7taBNuBvdS1i0iXSsFlwCyT1a4i8JI6
ff+P9Duv24uskRhD56z5LfJCwTqpmNXFT+nW3DtyrHhKcH9qq3vrVEISeyjq3tyW
s7MV2Da9HpYJ5LzxmxqmXu4+et6W5xS0EWA7mmu/gfEbEmNhDu3bahQks+wzykXV
W/dVnHbBTxTsDijABJlV9C+O4W6l9TO3DdJA7z5GY6vIK7GmFE3yyIwb7Ua7RquM
A+b6BbuRtjcpLBkggHtZVwARAjStMF5lTuRUtRAi49SpsaEvWiEN5rnf3V82lwow
bnkUnk7Flz5Hb07mCaGoIKEhHMxFTNfI0MiCbRI+xfnise0vqQ2nkiGk2RYN94fk
AOcRXMVbQt0mw8Hr70wtHDdeC7xooJmUJ1uC0eOw9qMj+yO5eyFT4wnC5eoZZTqS
vF5Fovykpnl8HABmPnzOZ1kW07/kft/NrPfb8wj1poIOU6kdmQpdkb8vnr/HKQ0d
Mw0issdudcP006Qatai0UZ5tuXARoP6dMdAwDVe5Nb9tzaqrlSyJziRD55qgcEqU
wZvZ7v1txLAU8AJn4+sTVIczTcmkmK0uYpxlx6HoluQSBzPPcKUR1fZfLfBfNbgI
E9TFJr0zcCM6u2KVe4vGDpl4vwjc3j/ivULHzcq+dvPqUboMX7PUJJSCDhR02LLx
cCiJ0B4whWNbqTZXia+irnFQntnbqq15kiF49+R85yULpPA94ublc6ccuUKoCQAP
EGqg9m02vjl7aMaapXeqYL9pQ0S51kXmHhLxSaFgQ0EIdKUYjnbloKS96btNbR1Z
y/MqyWFryWufo1KEBxUUbaa5jAnno6DDZkjW1mgOCni7kd5LeRZo4nWnnpDO47yJ
i4HFdznwOB4CUterPXWHiQli2U4RAtuL+KNpSO5/qW1i3XJFtNpepfF5vsvALQVX
htH5baP1tWJInCevUcyypFTO6fLvLAe29mqojkjvmakios1dBBEYExJy1TRgoIj6
k+3aVlP0utExnT+BRIdE22y3r4mwdy16najLCX7M8qwkcaToWjBt/t3ttVqGEdfN
LBtQ3iSP0tl4ThvBCQQGJVtrOE0tGESiqsWptUOnLR/qe0Tyqm1FD6l5tiieHOuI
mIZz6MJY31BWfjr37wYaD4HrvkoqSfi3LaQeqbNQtizfAxBVuRPptdow+vpbwJ9Q
YE64Q5xpgQZEHdURE5HZcvGAIzg1dBSL9/G/52qHPNakp8H0bk0k/hnvp1ck/eRH
wqgWTuZs5ghTZ3DSzKYD/PM2Ce9QioqyflWmN5m8t/c2M6eeZKqIAdbIrjiv9F6U
kOESJ0XYPnhqMneBd3VEh/796TC9jdc5Qb5ul00WIbNIq3hhTq979HtNRscyO6k+
Do+V17vuLES25eOOqFJce0HQZfauvrWOEfzDM24P6l0GCvjtTjRbptN/UzryMF3l
81ucrPRFI3j1pc8RUEBWOuP1rnaJboTL2AFjjB/L9ba5Hyv+VLAZx7vPQs7N3nET
gZvxd9YNMep+Q8Re9swuj/2F6zb8mQvkJ9q6t7Fg0uhiGxo6ayLITZ4P0EKY18kR
668PqZpb+RjpE/cZP8eZ7SCeEUejRF64jtAZEOnVSY8C4WzjgNC/NQ/YQ9Uk58Qa
WqCXt50mbV4+RARYv2ZK9Yn6UKqB63jEAB2pI42S0Dcu0+XivuJtMnR/cBIAfbx6
rdrbN/NJINKaKbeA5ckt9iXUFEhFU8crU7V0ixZt+Oe6up8HJKJogPQLbI+w/0ME
Ok2SKVjLrZFBGot0Qj5pAS1inQjCS3061n5InBml196wKro2cGU2giR9GQYNL2bn
UTPO5zhNbnFYIL8r55PUsU+M9xp6eIq70DnUGvFfumfZdx5rslI4j7tTC01tP1P2
GnujT9kqiYFp/kvJxYgSuTwogUZ9ZjWgh9VgVjgoLDYkD0YEQk7scp3KCqaLQx7t
JhaKzUYhkIjPypLphVo+ly/HCGmNrhy80M8KpF/AqdgsZHPFQBrJHb3coKMpJcH0
aYwmgmx7oS4YTkqJScGM4RtxXJVCr9CdjjjH9otm2uPrs9H4g4cY4uNqRqousJuA
vnCRpD25spwqtqAoPlIoVTMyx2c34m9qlznZ4HLQDuDT/QvK8RFh93mRwHz3Oljy
YUGGSflHhx0OdAltsR1SoSIW2+cs6PlUbsGNSLuuGGcf1D1warlMfmbQ9yhn2pG3
56wdckhqs1sLJpXzmFQN6SAv1vEZI7Qpt4nM9t/Vb/vogzMBec8uaOcA6+tumrPk
oRcd72eRWwvytDkcjQ56BeKmynax2bIIeDkiPZgP5+pdbUXTSE15dKLVSWDW9Msu
4GkDXDfy6HbsF4ftkxeXboTBSF6r9Q8w9ytKGT4oycBooiMCSvvxsSOVYss1wra/
CeVQ2pgdHt86vV/Vh7BT0bAz3ufbdoVLhKEqA54YjgJ2hAHMovVOf2TukS1h0kXw
K0b+SIke2qP+jseXV+LdREQ5SlO3mvjqtkQ0QybQW5cLS0J1yRbuqWmGWZ/xquv2
kr8sdDs5cRTJcEPtmeYvffNePenV/lBQQh6C5ilhUgLmwVQiWameqxzAovei4Gip
Bg+di5HrG/B82+VWTsyIDWUoBNoATipwhXv9qObj39uoDQd1LAv88gFhV/xlopyt
Fx7djwwJLpxMiJk5QzigFHpm9gIVFlxfRqgYrsAtcVT9XLAbRMSS5O4wMolFUYIA
vzuQ7EkzT2uHczqqchfs246YB80rrDHo9OmWtrEgwBzQYyqdaXYpOYCXsUYCVlHe
9L7sz3Zs9bi2iQHNO7djhmr2CWkwcjj98wOMsYihjiobWLBIGNcLwXQeh/jWE6k8
UAtKz9SKb3OUcldpT+wV+igjCjTqebKLe3ziJH84aOYWlr6gitB+ooSfSMDCKbiq
x/T6gp9BORqdC7uPASRPPWOSh7+wJNSbLdEKhx9+36YwGWjmqHW87nLJo3CVuOdR
xsKkKERrJIvpD//Uo3PTXEWs3ZG6G918eKjTsoGEBzxjBicvgyfUXSh0EOJg82pj
WADouqcvMaXRmGuHwb+sH9RZSwntU1xo5cusYlyG39Cs0lytwtCjFrgxS/sn6N5R
hafVPN9gwwtZpr9X40qeZgo6XbwJGwImzbc2q8j6Q6nRwGswSojejIZTUlwpaP+F
A0Bxw5+t4cqfWwHQTgCIpj+KigVPP3Q9CPEKB9dZ0Om8gutAMWVbATExCViEPHZN
ngayQXBmjxDRBB7GapjXbSuqEoAP4UvfUDDrWpmPamFtsKXwmSz8n8oaHjMlYno2
fKmwH2pqNM98O+UNDjhSPWE2weR55HLbONUFhnLFwcMHgWAOQ4xMn9I6VaXbRDN7
mZnkuoLNcjnNw5TtzjW0WutvFBHrVvo8t5lSwXfy3CKjaV1OCn/v4QUqk3eId+0E
sfo7oOr60flDUaaN0zBSGld0gaIZelisa3CazQZ7QqBS2CGVb4se2IDKHZg8ZGhi
5ztddjG4vmaj5NTUxIMnmk9KtKAD4LL8qjAXEe1ZEWMw2z6R94OOhlESe50ZsWgd
Nn46uLlPecp0C5XtboQu170Eh8lsHDe68Wby1rvQf7xQkdAko6wG2ljk5XMiDwcP
2DM2QKklpwYCWev/PMr5HfapbuxAh01MMr6Y3v89aKhszo973B2SkEfY0UF3sfPz
k3HpR8pTu7UJL79t3BEJnE/OcoCL0tJ4Onc6vroebi27G4Se5+1hfNIISoVk4K4+
ySyvfpZx+EgyjrigMci519MJpj/eIGR60jbPFs+0+xLoCM6dhnZI3RcQFvCyoeXf
y5k2dy+Ni2Xp0lTfpwWnqB6g2dwviiouLf+nSKypLUXZOKAoPNIxh1OIfttcfaOC
fv9pMvrU/G7uzCiNvuJFLTkJt6gpueG8zB62Zv6DWQGHGl3Ny5gtxUjZuPH8KFe8
g8SmdyeFgRv8+VYfxQJVEpt6quSXEgSnEv5agA37j4ljVcMPpc3VrGRJJ7yIpPsu
EAMVixwfy6JFLZlH4xj0YEY68gTPQt1j+Vz2jUDY5UhFx5ae2pMcByJvdnm9Ks1J
AjAGUxp+IAXqfCodvvgXCwA1bzNcnZqaF3602zthL2vqjTuhk50x52l7W+lfYnyP
Vx93Oo30xDlBJJEsURRJQQ3AwRxbS7/TLBd7pEiFTwox8Gm9RalerdBCFM6M2cpX
uweCJn7Hu9Wj6k6VcqG4m9TS2HuTgyZMj88D+23qDMgQcjlUedODN8wPYR84Nakd
ZaFVzkiAuAmnMWLIqLteyoryuu++GfSKO92MRXGNrftJRDoHGIGJzdvzYPgm+rgF
7C2PJgaE+7FXJiAOPj5OwRdq5mflcg0KMhy1CmR90B17jbMMeK2fa5sBgPJ07mGh
/0E72g7ajzyG02ymbrUuPu/3C5UKweTA6OIqFOhWaJQsq03tGS90z1D2vVuLhO4b
YApppIEafg9gwL//vw2qtdARYPD4QQVydFnUQMkoHcB75EpayZr/E5J/JMzKARKc
Flf09wnGndNBXXEem1o9j6fV4W6M+tQ7UNa20sjFWShvIOpPy9FWjTrjhKf4boPH
1WjDxuTQvmP80IKCd56gwl7WfuvC9w2MEGjMozT1nHJ89Lq6VZ9WkNmTZx3A1E1g
FcvODt30b+TCkBYJ6KrCEAxBlTH/hW/kxcTFUu7dEeF8dCg/EbbQmTUAnwx3d5bS
Zu2jgaVPuOLwhhSLeViY0JMlrmBXNiz4Yo4fsYqwkSww1QeZtzt4PFNrYlbZP6sO
RGBrEyZ6tguPMbzsZbhfF8WEnv7iPUXP0mrEeYH+6IE8u3NltD7yO3zyHNmmdg+H
Rseoe8wb52Wdk6RxwWqt2faUEBzLqPzYhM1gk6j02+4m9dOkpmNgeSm0Pt8JCTwN
IMems0fvFAbm1EVIcFv43XKUEJkhAdcX39hRMe4KD0w3hZrrHhxBdHXzpoJNg5cq
u5zk928mqdSJuwB6rO9+JmBhM/wJqeN7mfdUfhX1fBRSxvOaHgrT6guzM8bQt8pA
5RiiURYQZYzTm/2Dq8ORSj1P0RfLALGWXtUPddfj8cbYN6OoUIkyI7bwgI5KBMRa
eFmcMRTrlFAdO1EUdD4VqKl+O3qmFXwUT3vykkoQuarLAVYrv/OiEmljU5xsH+Ky
JwLxo6jr1/K5BgDPk4ReE15vA86E1teqv0DqO9F5B9i+V129xYZzel90xhYmew0J
BDwdOfwy1jN8axYmKDdFtthKDYI8vleoAQe18QSe/vifI/ckFLOJW002zsmO1gA7
aCThDgagjwX3naNKNTPOryZVVDXFfTHR7uI1rfAedCt91YCT8Q1JpdVycHZJ/GUc
yKDlGYSCDaxqIqQCBnWj2FuQqXhivtuDl8Ap+V6PZ4yV9Ef8JlQIuLnmQdCrGeFo
kqB8qdMKkgLqfbBwLpr2MEck8p1eR8HW7uiLKl4T+pSr9LNWYRN5db9OYU9IzTDr
SAZb6zbsoCZf0OhUjuLaGLo3mqoZwnb9sVf+f1KyBaGZBF4QTnz4P+/i5jTOXg5m
MaSaqvDCdBrUzaC8TCPQTcXdoQyxR/aA+M+jpi5Ri437gwAyY1t/NNZGieykZdBu
0uRftd6jM6S10gU8+mnzbCgYwg2rXip2Fb9PLL8gBfBHZP8Ate+t1ybprt6smcNS
psvKSImrdyWnMHDXEJhDOpZQudMaMXyRYAzPTqofmemLs5c76K3wEX1Q1EAQIEst
yVwWalgQw8ezEPg15Rlg7cQ+xn4qm+KenQ9F6AgnFrbcFsKLjRQxTGKUPCwd+2KM
J7+oIj4mjGPlPAn0PO84lgC14QgNF6IKyeizoba8RkH7uXCbpOAlJAz4NPrVLUOd
R0ZCu/xyJdxjGLg9Gh3fdO1jZwzsZaQOMR8+f9JOlnD1PQv/+fI1EHoTqehyuIQS
Et5dXS5VmzQuj6er8IhDd5s/SSGd1VNKCNM5lvoH7skqSsR44OI6MJzdCLfYsSJ6
W9pETnhUcSABzXxowoJhFAKUdgP2YuZ9pM18FyKjv0pzQP0c5+oiTm20r9RMHixx
mCA+b+nif3bYtohpdx+MZeWLbVdwAC3PQzsQhbjrZdco+jW0I5Kz1hM+PAjYpvTS
P4s6cXSrSpRKDQFVQNtbrINfK55GgbsRerwZP2eto9SxiHbtFJ7BOM5h7IkK+v+4
1DdXq4ywJVfMlMFBLq/K3tdaI/nHdR31uqvG+3ka/tGeWZdAw+Mj4q3cOW8SH8Sd
7ANzTtlJu14NREyKD2tiR/RlRw3W3ihVFC43RwjqyIl7mNmfY5Do/bAvt7CKW4R4
ZZHfO4PWQn9jZCDJWizMAY1qQxdKLqissl0jxpEHljrOTBpBtmVN6ptKiJ+bq26l
YU8zBS5ncPgt0+X5Iel7a/OGYrxEBgqacRbTpi+p5nW7FOOHV+NIm3izZuPzR516
0cN1ZoLByGuqDfufkQLKm2/BLwNHmZ3wXZWI3Btnixrg4dPIAXmIf4TBBDboj8Z5
ccGo/tSJ+ljpBhcA6xxkE2WHPLbAuGMN+BiqUTJ8uyfWBgHFckfAnxGhRTKdqviI
/k/m7wRJjLOEujID2P8wvy2K3UudSjOvH360xt0/jvXamX9WW75lRMTx73Pfv/Ci
6cS4V6xZw1cvgJDsdkD7T+4VWc/A1/mbRCEeeJwYowf6KTes8kHJETX2SWK1+86c
OHKuerqGDlOtdeT69U257j91eGhbgwXQJeSEha7xSInrG4M3pbG+sTWF04P6PBKm
MitRr8Erl+BBPwWDeUbxS7PjP/XJ1E0OUXjMwk4P4gOFrkFvcPZ2j2KfgLC1WarF
EIbxjrbFdMm3e3/PIs9cwN0c9qbwuKTRjVOHuZgZFEZ0NfvE+PILpQmmQ6pI5A7I
lr2A42A9atQ605Cn1tzeuao5wJghbaDElEq/ibAVyxbxNvjQsHAwda5BJAcpSpmk
my7TkyRCQV9Woz0qeBeTqr1FCV+PafnzotHN2KetcsD6DP26fFisoZdI01oynfI0
Z7ZH1iQ7gfVJAZO2iKCJr2Uz+h+p6T7eWaidkFt5do83TIPDR32+dDtLcj780UiI
Qe5BqvhHyPFLpHKXrJz1xowS5/O/MUnoxdRpp4WUL5Ur9WIHQQ0oi+Ih+4vXMbXl
B3ILFBeMzrKR6q9lYNo4tcIyxUG/UH14RlvdbfTqzonL2ULlnZPvV6TqaVqr7cnG
ZOlntmiE0y3/Y4ejquorqtMn/rgA8On6BKohSV0TUSbixX3alDCcVQqmNROJD9Rq
X2jL22G+qJY2+eoH/org39KUvCp7CnYProjtXoZgZ386nBkIdOdhbNMPFaug+aVl
3zN+KsNGeN6S5p89grIuwFJlCrm3/wOkFEKkO6a+5vVGnqTYX4wa63MBIvHNuq5j
9u7+jz6rEXYA1upk2kznaQEwxvJnfPILeIhxTvKHAXGxjI3lEShvSfZmailxYKqh
FUYzsTeH1HgHUa5CXHd+c9KK8zxMmyJnCAYrRc2wovfONzglzdmm2i44ukQUHHos
laN2cfprn3RssuYo/9nS5xBDfyqqCiXicRKO+EOL5xJZJyaPQ2A7VGQ2ef4M/+tB
pXhLCmFNqLCnMyDn+DhGeEjq47Nyt6Ual9jI/m6BpPunxFU1vjM+fVTIWSaBLSPN
1riFBN+2TBDeBNdE/ve0QWpYEpMC24dFcwYvVls37k0xd0eYfeie16apsoIa7eRt
/k+DqZjxR828NVlIqLlEf6a76AZa3QKKaygq5Y+0u606wlqWxzSMyS4RnIKsQxrM
nxWSDJTtQc24p4U/8KaXkx08dIAszEF4+Dbe4CYQdOjQJFkeAV2JtAh9ZCt1Jsgy
+mAXKiMibauij2yM6ZpLS0I3iv1dmZXz/0EfD4uhPgC2D/+LP/rpCmrlwRHjumds
780Q6Vk/gam2tn1/UIy/2vsr04OjgpHc/2sojcW0DnCKw+iN5Zw7QwulRCfCwKj1
fd2qm03hima1Ubd6eJqSGLNq6BwW4O5RhjCjn0ja/Uq97vm7ru+kois0KIYHYwL4
eWNh4AnYoAWeYUkSP3CGmI7l1EosDPJZLpWQwnvw2cY0HcbRrOO07oeLD7uEP/xx
zMIkldwPXTVS0FdLjWld79T1ePDWxgoxSsrWhFHUXiQRq+YfL4Icf6hKvQwsQ3/n
RtB12C7fC81YcNS8BylwDtCABt7KrmJuwRKpdv72eLLu4hw/DylYp2wwzrrZGTTy
ilF/DSHiCHaiXG/Qj7TrlZo2/Lfit4AAaS1XBBIaKxevP4Af+Ka7s+qUS8pFZs/y
avHNOWWrk+5G2QADvRrHq8n/RUkYeZJ8+x8skzWzrP0L4lDIuSULC6VfAuXrMIba
JD/4yWNcPw5uaZRI30N/yir9G73fn4wtjdvyPLi7FxzldIlqGRWsZGLm8elVREUA
sXRK6c4Qw43RVmmKbeAKBvhQR5r6hoNdfmT8aKkv3X8ag5u4wHQ66OGnltlEH002
i6oA9a3TBq8nMYStUIKmo32F8c2fct/KSbxD07teC3km+arGs39Qke7NZX5KNZGW
/srQWeIPSVsSau10eWgQvy4vhCIdKcb3DhCnXrZ0HLKXyeLdpkjPl8DoRddH+SK6
5ZuunyRn1lgn3ySP3l8nN5n9A3gmYHcoxykkz1+Sej6zGunu9mHFpZ5Gqan1MVXe
/t5EqQzj3OR4w0fOd+yEyidjzmTfeZ9KDakH2u80eT46DXfA1gIELIt0N43nn04j
2msKVzDq9ac55R4GjFV1eAeIFFd2njorwvQZzuaPNcW38p6/N5C9YtlmIhB3sRO+
CWfkyam1zfPh8lTPM189HJBeczSagesohaWFyKhHLenM98ANRwuKgGimeYTPlL8C
IiuxKHUx8jvGOY5qN9F8C8e3qC8kKTLE6NMTzRFPWnlGfqMUeJzh/mUPrVPzaxGu
BJ3jo6HEOKynUCzjjk0DJxV3yyotcbAuuJPPVmj/bFMyZOvzZ+18vWHsNvq2YVWF
/5wz23RHMznmP4eLOeTDHgbJ0NuWLNh9ijjBYwQMvyh8MbFffqY0llfbl7nQIyH6
YiqBcpz7w38b6+k2HzEmcgmRbUbEe4W+RSMwOWh2Hpmi0wi9YpyEZKvpkydvmT6R
hnej8iBtOYj81CkLAJSEn3I/p6JJTLa9vjiVrvcEwpdGM343SPPDNAiYJugAUoUt
yCGvizhFUYhbVs2au3WuXmm/QmlzApJR9se8aNalp9C4FX+Ugo5BXg8cJMeC1nMr
bwRm/5ulngms7sLGSn2LLrCqtk9ccJRjhG3uGV34KiFkFP036dMi1UZgmbKGkqNf
Dfs11mLcN/O+GWNCSzfsHHySx1j0NEJf+nERw1GRmfCis8WsjJZu9x+zjpuNjE+x
KdsY+nMWXSPuGkt5cIq8RcdH0V/O3f+IzMMHMvc+kEKAnmBnadZL7sqM7fcAn5Gj
agAnuYoHPwJltVdYQt1gxP0BUUNtcIDiofJIPy4mNyEpNEYUkuUSf+CzLCyw6+NI
HpulfjmnCHfH1WF+sfbpp+cZahsFsCLDRIcrUsDdAdeq3yJnQI5qNb0lYvdN99nU
EQ5QWOoeaBWmQ4BwYUj5MN5Ux1jbsNihMcIpTrJeDLz7EFqHemycRld85GV4bGAY
2fXsgsdJWYMDhJ8lsLrT/Wk8wMCv2iVCV6gPuX0QY1kThOSlWWpIjmNqzAvRBgx4
/Id6jh7sauPsvsDqhJm4cG6XvdQle3qB6Z3ybrXLAWZLWYQTJllKnlIyZKYWMloF
DCxDXhGUMfPniaAnHTzSRd9FclglWHQTnHK7Vu21ifFo0RK8hl9MJgzZdm2B5scF
HwQfvz73Uh8L74ExXnITId989OZyX9AmS6CUXA7qKXYUr8/GMkJPXXH/XiNcBoIc
wEV3H7FxOzyaOhGkWXAZHUvHEuJdb/oRuSiddHbBkIIUPoE3bVoJtJnUCSgvYn1e
qOvQdwHyBKImsxSzythBaJiUtl2kBq7xtO2Ov1j1+VtpBjRvxiVmTAXUt2XzeMAd
R4fwW6J9X2Q5hqfhMd7zmIwgltuM0ZCy8X+zX2Dn0JMGiuPORaVm+kY+k4o5bArJ
wqRn9z332IHKir9WvW1hJ++yPDcSUxbQNowwAOCjklVdBblDoXZXSZfPPF4M9CkF
pw0oiv3mUOZGAxMhyuSXMyrPKvkTeI6fBkpMFXkgwsQ/JBtqHelyH5/TyUoM9Iaq
FP+haFez0LlymJwpVuvwwNbw7Hsmbookc/xHA1hDzbkAuXOAoxy/D51bj5q4Zr61
PWPVt3OZnmWjwAMJTL/mcSAiyTHb9zQC6B/Gv0cdpivhvEuCmIwkd1DdU/gRrlz/
o4+ZXK24443pseG1K0nBilK1lXqbQ2ed+3702mF4l6SSdnVezEwgKs9gdZHhVFOE
hcEj4bw933c712DwqZjrvuRzZDl3tiUgDF+KoBCucsXL9Pnh3zNSbKiUycjHD0V8
MbdyDEBYUs9SgpBsUZ9wU6DIlCusR9KFNIOhlwuQUiJMjpfmYh8V+cPdKPB/eB/p
fFDWP45mN36zLJ/fYh5aT7MwoOakl1/J9N+KrBiYIgqq+lYOwvR4bPs7Usa8phOj
oU8sGnx5Jtd0XWOPKVNlxBLVbcuNixXJBa6/umE488IC5uNLMEwKi7wrchmhWGKm
QWEHT/6A9lPppN7Ycm2c5iMZk7tXlQ+dCe57e34cbjNvH9trWAuFZvJ6vw+Evl3F
0piUB6TtGaBQ4qrCKsi3ZI+Wx1lglIc4D+qMORSWDYoOC6ZeWC9lRDi8xtNhZvNj
tPH640tYqaxxVUShb34skWhLe4BLgnNFq2N1myN5FkppVGyLZeprtwDlpovsiGVN
gxNPPqMCL9QyrZcK9hjOb4OWuiwunwprl927HdlcJcE1YldQoaC8ljJDeCDp6sJ5
m6YQ0yY+d7MtCGQ8gJIFciFWV2TyB/AuLyvhdKSHyEm6HvI40gZrVxH2nHwNAAGM
oPjp8e1n/RPW5Rl3U1x43IorAi/6ixoAAEokHHm9SSDTTYPF6R052m8Fu0brUPIy
GRnnmJ9YMF1geV+RWtC4D3/JE/1mWjXJzRWQudSQIKhF0aVktBO+OeeTdte61rui
jk1QDPMJBl9oVaqesbcFGNdCoFaBfTTdl7TLAZWB/21N5f5ZxqcPzLqabCnmThlU
YQjcBBj3+B3/MuqzTiUqAZd9AjyKNWLeLvIHOyIsXa8TMTnQ2oSlVcjw2RJ8MzKI
IqE6s5Kb//w6n4SFX/H/rScbMXLivdjQBX2o6HoMeKY5nl5QWOjp5FJLkfOGGGcS
1XwW6uyqXv3v1+2dUBifShPyv23it0XfAAUh0UAkiXPCeP06A1blsrPIqjc5nhPP
COYyPZZit9ikWS7Cu7b702l4Ul23Mpuo8foMqFijDnEizkiu58HNjfQZGzFqrKFg
+vJ/WgSTlEihPl2S5h+n7i5HvXzj0nncBbAgK/V6yB+D4uHgqyh+2xz39wA8J5MQ
FAIFMzxTYjCaUSBHVoIe/5J2UYRKqKXWhLJLv3Ysf6SjM3icuzYm9//0fXWXC4GM
Rej4E/exOqa1TZocqU40u7jioo+1JcY2O+H+Dpe+V0BbvsTewoiE0dldmcNcyGba
0dd08CcWWUZpgAku4308HlLT7n4IL1dsz7ulPMeX899YgXn/FLbGIhlLQSS886yW
hTVidiYBhUoWW4FfTReIy278c+roWdkq/GV+ie1twf0kLNzIcJhXnF1QjZ3WxHk4
Bv64O31xtNC/j215stkv5An17veyVmm3jRY4K9OJxTb4K+jLjKxtiNczLr76fdBU
NVdxQETfxQjucxxWJuKnaz5AUi2WYwR+Shhf3L2AGSwzsr385u+Yr8AlkzhP9/Lv
HX4dU5WsWYPhcwFoULyFry9eCHG6tFnMu+59ITd10lQHiHiE42XqbtKLG26XHGQ9
e8Y8DpxdlqFM3jw/2OudlWRd6xtiYOTG+s/TYaSi9PkDOyJ6fqInGiuWTOaOb5bq
WFpoH7F6YUX1VgKnXki1VtStGmk2+dGrJ805RGtZkVzs9sc+zKBlUSfGu+VqFA3u
Imw6Jj8qWY6ILPaB+nBWRHSSvt2zE4PaEwaEmcJSvhtS3jv+lkclB92C5wdqaq5y
z8v3GXd5kuPZ86O92MUVP3SdUuyqwtkYMx35t9V7p0V4bW5EoYJkp9bc/XorpQJf
6MwjP9vETE2Kl39yhcFXuiXjOZID36TasVkl2kx5P+3ThX3hQic4hpDn/Y6R6xy2
wkMvvK88Xm0tSbxGUm5gKk/BuH6zJGUZIII9kv4t6+9lk9zcz/Glpymk9qZx9T3r
eg+IyuEG8KZDxLb/W4uDAK+t4JojHz1MEa2/95tnHFgESHd8vThC4l9KJtX2BXHN
T4lITaTszJYi7RbSrBMgw3MBvMXXpkwUEvYCZgDXNJGJ4ZqUe+hT6t48XJ+Dg4xa
ASY7BB9SAevjSaJKaItudF/RSuw9/gupU9bqAIGM12sEkG91lGK97KO27oY0pNal
p1As/KADEvNUE7TumxFQLgCRqOFrMzstPdiRWpkFHTpzcFzHXOT8/WwI0JAH4Cvi
ei9GB1l6AoVSOjfE2NRg70exg5q7xk+QqAcNuU3X4b9ylx+MTXZZ+QKeaKJaUrwd
/NOg+WSSxd1OKiGyYE1wsp0zdjhSPFYlFdr0G6+3582foUfKaYhM0qV7t1Irx5W1
MEeLp2A7Vw4rFtNK97MxwuppXfy4OyjJd3WQoVx/mFIvKN761dmrXaHqVs5GvK55
89PeE31l9NMReV/bygoKRnf1I03+KM/iCBbhuUlHucKyylIER6XCB2d/N2LsLS/d
eExMaMFukeDOazC3ejhxnE/IiiKeSxtcTBmazAYoUhU2tzjHm+FeVbCIdT/MZrqt
+M8COOMPHIHIKT1NCM1GCRZMB7NEXcv9eNFRqOR9yIr+5G9llx4dgVNDABnF7nSE
BawEZISLDm3dtor8bfAhqnGb+BQJ4XGJrtjyPAwkVqlFfk7KeYt4vHbTyrjzlkTa
dvdoUFJ0Jrs9HNY5Qn+10tsCy7PbOiLqazEFcU4MR0ZmtoWPQySUi+qwmJCFUdX8
uGONAvvGU6WxIfvDi5eaVs/xY2RWFnHttIM42GeMNs2nYB4wnl7LRwJJHS0OM0tE
hY6wpifAzTMOu6UAJ5mwZaJwGS5ip2Vj5obeoI5FRTxpkaW4q4PzpEo1Jqufte9n
gx3bRZJNeUX13MFp2mZK4L7dFGIGwwdgE27HVgoF4ANgRFdjDyL8X45+qiJQdP2d
Z7xCwsCFcjyjhVcJn0K5w+N+bwSkAdGXdSpS22Oa3MLdXH1BEim/N+3xpHZ7S+T9
uu/EM2fYRMULzlv6c+vZ3gQ698QQCCz9jzmXKmFFMeIlvWMN+WSpZFqB7As12RhB
RvHhYcNjE+3e0Y+mrVjOncAMbvUAv9vyeGAtK6X2/UcQz2OMl5I14krjC5qaXd9p
amjlWqV1hKzyOyAwsXQNH5voyf4Ebe8FW+J6SdFSuupizqg9Zdgm3M8Yo3opeY+R
HBIufY5tS22IG7wT8Irs3KuXy5ICV1HH+MNNXWUZRgeAaReOKC4vGTOGPYR/9iSI
bAYS1iYibhMlDkCpC15bYegkqtLN4dyXJgpnvl2jl1v+OGQJR/1/uNSXwWCY81+b
iaP36bhLvlAkCJ+IzG9ehrc2S8EMm60IZNJ+CM8Vwhd+YgKDa0qsD2jXq46saJRC
0hQMOI9FmXfWwa0nmyMbxMxibw0WT/vFMxhnjA/EdYF727odbf7Xic2rfiVhI0aN
rkPbAlvrWz+oFCH/6D1Byfazjluh/2MptDot529qLn+0aI0AvZ94AoA/oASCW59h
eQyaRAyeQSXHGNICf39Sdt7qE42ESTgw8yGI+a2XW1H3ip2DP3EPFEy7hynsIMsj
v/hjANbFaWhUiZjxn5oXNwkAsuRmU0eifz1VE8FDY93ti1/QYETblEAPjA4/V3r7
5tYSiiiC1IIHxeb24k2fW4s/3UaeJO8iZQWHg6gWGVh3gUDhg3+Hu5GPPhfdsspL
c1n34a+FT51DxHagOof6ecaJ58YPB5DugcOz07AxZv9JoLBqk5zeuI/AeqdCVuFx
GlDJCPmNUqgpxx7Wy1CFCfk5n1PeLIiZl3tRM+lyHZozzwmEWYJPkS8mjCVNFrb/
M64Zu1ZoGJJtJz6wDI1msdv6NREEhikjgA/GBIx7xfL7ZNNlGm8IbjmI1BqLLC4d
AqzPC1NbUN/ktTg3bD/Dpz25plfBfs6Jxzmm26RQOFgPGNsxZ5ILImeAfMZkqjk7
JWl4rPHgSsLURoWb2CP32itK9fcWrNk/Q0fpOhum1DJAdHNn0gpfl3DsPKnfmLpI
c1Aer/H1+4kGI7PrrxF/hNsCfeIPTrn9z0kHvBErqxDEMskWlHu0oXI1dG9pjhR2
wPHBNdP4ZrmP8NGH1LSmzk05YdzXLbjPIua1S16hWxNj9jJO9sthqDJjoAKdiNd4
WhuSoNFLm669umsoTMwpu8ZMj/H5nLkKtmDgt9qvE1LpHQCWT9N6ZHzLjYxKlvzM
mAJ7LGWovpRv+8j+t+esaynAR3/XSSXdLfhyP0FyJwjhlxnVzkEWRkch/MUY8Yua
1RoIJcYNoxyKu/cpdBMv/1nIxF6nng7v9tNcJRg7uM3HTtNbqLvFtSMVriaQX/9z
+TaDLTmctg9ZPqllntwnu+s9KSp9iwakjvhMqgtTgWu6YcTjW6kWxA0RaiWYEzNE
l2BqbC/k8CfxRPjII9BmYu0j9GMjJqumsrAyZPWO2HipoeneYYjBB8GVs7OmbGMd
evagZ8HOm4pZW2CTRiMZ8XoKlkZvffx9SddKbppxOHNAl1uRCgrbwrlkEWxUYHYo
Rv+WMYQMq/H17SOmDKZWw/JFzkuUXK42kWKwRkUmVGJnd5ytEErI1OKvoCqESYZE
3+bu2S0h1Xzn5WK92fygDsH/nHeLt0DqdXec7J1mkJpiVSq6g3iO1hHqr/reCoRX
TQjy238sHpMKT+uXcRMkqwirPqYAu6grOWPQslZS/ydfTGnhZ+mf2q97eeBpM9ba
LZJ8N5Yk7Z78H1FL1+t3ROWTfHZHcH8wOSWyyQVpylrLJ7wSqvXZoK/W9YMyXiSi
Wv8Mb1Uh3EldIjDnioZWT337NPPIfz+AiV5CRHc1Yp30JPBRukfZrYx4nmTfo1ti
7hnIlPjCdTbYxrqDnt1dFi3orUGiBovkzbKoIxJS2l+32WbTIn95aQmK3SnH4D4z
Gm0Ki4BegmADNR6/a5aaFaanw3FVBf/e4r/VODKJvaBCZ9Y3DqAxsH/eFW9hspeK
jBbUm+gKAjjAXEHtb27I1WC+uj8IvSFzcXsRHxjYko7bGAW0CBp3EH3jwFJFvEqP
sCF3Pp3uZYnEVed6+qUb+4/ki+q5eV5bWppx5XwFqShb39vgrgZWvbDAODlmm2VZ
LcEQDYslSidGbye6KwgB03kVJN7QkvN2GlGI7/WjBQ4Z+UAfhFjvXjltxCqxUheZ
JRjSkVgBLk0DR1nBk9r07fMwKolo7n3XnRhZObVvZnAMGFxFFawVnlTjGpXBlpW5
lavxsoEpnQm56zfRntcMb7PP3/AAOzE4jAfra/C5ImbRMAFBu+ktIaYi6000IP6O
dDTLf/V0dMFh2TEmka1kGVdf1ROSZMACQUpn4Xh/aKsQjH7yvpiVNbJCS8SjoRLG
mA6BuBP/LrFzv7b8az5d4qZp1hw/xxD1ci4lyy/gJbHkCwVgz6X6E0O2veEjWl3q
SQFXNyEed82csvnBY8OBrMwWHm9yux3iocR0achkFRCW+ev5qOLMb54CCwdbt7Vj
HOPXcTpBr3PqxKQuhH+GikJgG1F6xA8yWD9zhEDWIc479CR9kUhRtgFMhcjhEdku
IekdiZx6xkIZSxsNYeHx5PgJZuvOkeiXBauj04imFKOeUy5Fx79owS/hwn/HgMTf
p/+10Sx7LkoZinENV684TsSYBnhAcvwwPGBx00gL6KhJa/4glwUqLnwaJ48Wi218
ohp81Qc7CGD6Qk4kQySMfHwfsiKDwZeDcE1tgEddgaN/YhkJh3/7bnMscyy4WNmA
nhpue7xNVzulGEWaD6tdht/GmwZ1Q+7xMUDllsgsnAUW00ZW9F7VjXf17bbD8dUQ
Gzo5DFGqfcdUl2eLjvc+zWhT9hwXLBGA1EFmXuVu6l6jHGtKkuwB3jQDKijo28vP
SQ2iDYEEbwoo9Bg94dDKB3RCVvneYry2bmMaC/k/bRgJq1QII3AS3/G+6Fd9eO26
HDUMoczDEICN5+7acXY5lpLgP6NjtVB7f4aJfi/4Xrkd5J/RCFJ8I23EmiFzBMFQ
XTJMHh7Dg2COIkzQ/pSI2SMNJy4yPvtie2quGyIP+4E1r57rTqN9thwcEkWBVnsJ
z5dAtfztBdR5mwc6hzy9PUhJLkLNmXO3ehEQBRTWOjmhUsPSmW1ImBXVxo3qWkaA
O45V193zbzt+37oYDnn8tbmEeXGJfeNbN8kVSY3Me8gmhSK5PBxgycN2uUWKTC+t
3UjUz7TB+pO9MDUkYTI8kN+AVHS/zrSEYvH019hFcFOxASauZkhyFMFihws8Vbx/
gq9v83KF4I/GCr5SIUnBDtWB7hc8WLnI4pH05L7khAsgyuBqscc+vJVYcworIxNx
Vih68VoPWOWIIRl3xFSzA0Qu2LI0prUPNRdvBhVPlKKPJihK5ALcPPCS7EEAKcJz
SOR4xI0A+2wudorrV0KU2TGGvpyrCUfDjnfujYkvWJL3Tqc1HYKmUKyn76gNB6fh
QCENUJMOiWliHWnn59PGf/othoiexYuOduFmaAsCzVmCFEZsPqtdsevWcrNVUlkM
gFUwQegPZcr/0ajLCADJCuMOlIVLGWfTBO20mELVtYiC5n7OM1V7x+1qYDagiEa+
2ivkvPAizZVWO+/Uw1QqRUzjCAnC4ySqKKLEVYXeiG+ftxRb+SszmI7+GN/c643a
xTwP6KkVuS6pFFxUTughd8Ix90sP1t4PguPouE2as1yOXGeQ/dir9MySbdSSvnuB
dvzGRwOEMp926NCKs53RQs3wHvNFHrKZoj+hw9BZCB6xRTcmWS4KrD3no7SvG8aQ
wLfS4LQ3RGstwgoCLvtlhXLP/+khfkaphXCtWJ8cnneHqHixLF+sXYnJ9CcPEiST
4GQ2yFQ2ALHa28Gm/bih5KA7hQL9egHvtc2A2IIxF3S26e7D4Xf86yS+wbPjKL4h
aK7a6T/CkAi28B4mdsPWVhfb90bRvrbyxthDi2mS66gchWThdF741jlpwhx0kgY5
xymaQAmgfjTEEGwRHOPWlT6EnUiAFDYK9fUtrlVejrdryKcpTQBgi4xETipa/aOT
ei/aycrcNILWi3/kWFU3Z7icTVjY6U/QQn5gC1t98rQtTm+JmGsWmH7pfD+iyVCE
LRKNOreUcyTltSqGEmTfEjQB7PPpOx+TCtCZxITsXl0KnPth21Mw8leswg5nXjRo
c8XH64o3xmvZWBwjMqUeq/6lt3ODuXZnr3ebM+zn/61+/r9YpbSRclrqd71s9MC8
uKC4NjjTjWdVcTy6FbzUb2YEEr041gR8RobVy9lJrBPqF2RidswzOGW4NI1HYe3C
UIAS4yjc3vkh5gTYbzSKY3eWbt0QRdVWPTmssnbqbu66m/phxNjL0YqQuBPB7jaN
aWnj+bSr6UD8dQ+T4YqND3uxDesVPUjhbu54SCzmRxUWPVhkU45GGsCe9sx/yq61
h6ApGIWiKO9uH9/7NbNGZRJFuK1drAnl8QDPUmFedhvshNWufRTZJkZVULQjuuQA
4QUJUyl3Begyj6o/l/wuhsxLNGwq8pWcTd7C52gArsrizC4Pr8bLVWgg+D4guru1
mQ/VUDvL0yVCZS38kMxS2LUpZPtaYPX9jdYu7WOH9JQhvuIrY6rX8yW1V6tOX28x
MYYeMdHH0XMQ2rXHfSmywX+Yoh9GVbK8zKFJ5bEeSNUawXqtdgm0oNBZ0bv6fKH6
gcIN/PGLC0tFOHEBXEvZP0NaObpBv1YXKflXc3aSfIXobjWcJ+uKtwzc/PIjW4Zo
A5X6pJ6kpGikdO2bnpIJBjrx76D5D6RlEu5CbsGQlDGJEIALOT2P55sKCr/LVca0
Pr+txqNRq/Fx2aW8CmTBmLEEsXwvhhwX/KV5vh69AQhl2iKwHgBS11I4rlTQDdKc
Zb3v/MY1Cm/qz45X8Tsrmk1nnq77P7TAn/MNtMSceRg6Bb4hw0sBhIrefbv0M2+0
mx9iTzS0O48gP1rnOEBeX/uxQwTnlo6DsA6EgKuXH8fVWnVqvSHmajfHT42QiSI7
7CTkAezpIB5dYu0aNBjnStYlC3aU3/ySxJUdivQRZB39s+VHKK9F6Vvp/0autJWd
kj6BMzvQoWyU3wjBEioTbDWO1wNyDvGgvB+bzjlJwwUQk0yN433vcjN9mUx2wDfK
lB0/wL9zlrP5vdV73JcDcjnzwnl5fteiCZJCn51qM010JgVt/WzMbr7TeJS6EQb9
Pb/emJ1+vedOBGTurN0d8OQIlLUcpIQdWaVr63TrBpjACGVnZFyQNw0zAj9/iVpY
cmg+2nOevWlx77+OmxmOE53dO6NVuUWWJMJ48rU37/f+lpzxG8veGpejNSUsbvJ1
AvqyOKBT0hVChaxXngx9zMMNrwt3/hOw/yCKNj8vPuTXKZEUkZkJv9QKx7eZEVxW
HqZmdxjdCUdNcgHg+MawVU/9bygrJ74R9PsLFVVmlCKk9NrpIORGX0BkSbXda3kv
5TsgoZUZWnfiZ3BTjEWuJ9nMmGgy8rSGi7QVdhPkx3lY2CpIUXJ67WOYj7RNadWl
34NAVPc8qyb/EeW4pvc8lMeMJ65fuEovVfUc/PIj5fZ8/eaeZvmBQLFJUhb05Gok
vsovyG0VJb4rH0WPQJwp2uXsaNaQAqLpnIDF8V2D9R9IbcrzOJNblpFNiuHunEAg
i+gEgPWHmksDgE9b9XFQ1m9zsbG8l0TQxbdeIKqibYCaabVIu9GnlnBlMom0F117
OJTO+zRY5DTA77LQ+Keyi/nMnxTwxDltpXIxyE59tR/Yf/o7itWC496KSVzr8BnE
SqgkajfttBJogE3oJ1M6pUdSc5Qiy6AVZaQaX3WE6oUc1anaB34XfQkU3WjkI1kt
Lf2pobmDUD8gLD0YUoMzJabzWGjjKoVygU9ZOgb7EnDgXSniGqn/mitq8EgCORft
MYKFO4zCy1FsTxUubrtETZbUyJUE3Kd+SNoYRCRzdCkXt5hRwXnqR9GbQlMNpat3
mXTIPf4SplkesW1fvbU3QWIJ6s7TGHB1fFW7vXjuSdm0aFsotA9XWzwJmAZQ/LFW
P6Chi/It3+YvcZIk8OofMsHIkOxaUmC+sBYiGi3kwdCWUESJpvzOIXJuDYTEiUIu
Dc50woIVgT/tZzgZHMrw7GIAGYuE5qumvmYS0wjp4c2F/UUKgmzY8t/Dw+zUgLij
KWR7e7oCs08ne8bRDMCgqXjC87QIinQJFSQb35CWXYB43AI+JG84oEYjJIXlVI3L
502PSbw/8NnJ2oyO8xc34Oy2q43TQGF4S2n0orzN1/hmKvnWdsdsCpSEIVMHtpor
r46Dq6XYlrhqAtdHBBac9Xk8BzDjw6MyEctebG4GMcH/aJfx9//mSU1hL/A0YX7F
gg3aeeO+YUURv33/P8JjiD40RtL/TemApEr/cKvH/qW1ewrzkiCrtfCqpylf/9Vk
E+HPWf1V6+Kb5sNjy+XIGrUC9CyBaSwxP3SBD/4YifouYIm0cmrgIMxtoNZP+TpL
EeW2Qn7mdrWO3/OTPvXha8f1F4MFrKuWa2pcaY5knypeEdoYGu4a6/UoenVLyhMd
XDoffpzO0jx6QUX0oEHUg4kMR0gS5VEuNbW2pc9Q8D7BxWt6bSpgy0LxXW/dZ4Nu
cuTkGWFI8I1Kpg4RDG7iCQ3CGMvB2XXo6fmPzsgfGazo/cQuB+nupfZNC7YpSk42
woOLkqeF01tknyZbJXBsiNoyz334CM8FrF3IxhkahLVcqk06psTXFFtUBgAGJL1i
wzxlPhhplNYf9y6oLqLP6Nv6nk2EECnR/1lITr7V2daobo+Zq4GL7XI4sA9Pc7o5
+mzppKakZ+Bl/CLhlLc9j8X6HMSN5YXEYvyxtD+MxOURlm7OlGCX4jdeppyyHnHp
/BhqnqvEyIvPj0G8Iv8BEB6Mkq8oi8t6KV6J8qH7WJSkn2ZI6hPpJZGxYLFwZ6J0
zVwmtjhI+IZD6OhlKkZQFxPIB6w+XtSxwOZ7HnT1gn6zv3S91CZPcGK41jeLbQmt
1e4xGJI/lp7hgO6y8E1OMbSep46mos7P7uPNqmysKwgf8WYeORhmiF2VuAsEF26e
cFFm6PQ7SMcfQcGWxMLB3PG1IM+he3APa+YqDgX4iK7nPjZxTkBQj7V8x/YZwWei
UiuZlgrJcS28mY6pPvhxB3N+3+R36il7+M60azTIKqC6vBF0kV7vAzsT6VMiGmMf
6HfLedgGNXOO/bn3X+Ul8nM+5NBP6xmKyfhvSVWXMsCPZiQDv9XnpmgD6umvxBbf
08RDoruA0Mr7v1rmWl/xMjoOg0kd8t+gRBdJMVdbVxTXmHlvA/si6dg/lSE1u06v
4zmj/RBzsp4SlEC+x9zgZrTqHU6TF2xtadPxJashJ8M8YCkMwB94AW5uBTZ2peUZ
Xn/HnSbAIyBXVICIWTINrhZoN80nX6BEY2UFuwHYBTMMvIkYcUNsc189SQGkKYUu
aTGSlnNan+egcyg9T6zIPy2zsJd9EpZifJ5ODPbG7RsqIK2LBukUmec5tYSKEBvX
swLRSShrkhnPgjpERJWzLNJR2b3i/LjuYyOZvGps8okuWFNF8o9529zDOr9pu4aT
NlexuvBBW3IEOQ+Gz0He3B8g9h9No79Y1FLxKM/jwq+2FjifAIILM7XSgUBtQNvy
9v5OhuovYS+CL8GAtkW/f77wkxz6NQwnR3yOSPNVTsq+6WQAp5cMacmqTgjJAV7O
QQvmdD1UeIoh/ZROqT4hcjNYLtydLvcTKzYSMiT2DvH+yuGZu2LWkPoOGZZQVJCj
HmdXt+DWvGWOVJPDR0fJPtoWh5mLajcqIskShdBq3LA2YCNqT4euFJi9/BfL6z+a
5oE6+mUqYRNq1KWlQtEpgPTIucO7PSpmA54rz1VcZNqHPx+r0+3/B/xzBLd7Um0B
F/wy9TkPkWIp2Oomg3FwxDuYXBrg7JHBHBUJHAz3V2AS6aHxq4XmIHClE9P6FPcR
IXq8rlVlm8RBLqDnupJQyoz0S9SF8F/R2dchSlwa0rgfkmi0PbIRM7Zosw/bLVd3
h/7qLaFv55txGPuHRHnwqgMdW01k5lePGobxmrDI5PIC4t8mSfK1NEelxHWdx8yx
m1bihOjyx4zPY3i4NLhb4vxksdRa/DN4L3sBqqlXofguCcHbAk2tty/tVyCd+pUz
J0J/nJOIPoq+BxiAveWHSKYXfvYnBHQ9juZ2oJ9e39l3gF6xx5FF232KWEeKoQmA
k9tR8odH81FXojc5e7D7gUNPt1HHZyjh0xChXkn7gWjir/HjHTnDJC7scS3eASx+
adP03/RnbTOp0ZYBviRJci8Huw2erAyoBwBRXjV952knYbg6zcewtJjX0tAqIEh/
aBuNykS98OMhSNuQfMxtx3jc+L6/nKz7Kta8kWbyfp9knQCLRcMJLmYqQQstfqwW
eubMrhpoXgukGPPrk440GMONpzBOlSN/BScsWpaO8UEUiYZc8LeL2z+7bMSLp7Gu
b6Lw38JwHnZZgyMROyic4zVhvGvMBdQ2CjTB/fuBrUQ/LPYijcIu6dBWWSyQTC+r
XghJWjnDEtkPhpOFozz2BYHHxGXHJK5qHfT4K40lwKVkspjzngVVLVm1KKqtvYL3
OeD/AaEP6XqLzXJ8Pj/uCEAyMG7ENWw2uNSxEf0Kf7CCHk8rrshc60dWa79eerEK
bLbspEKP6AEFRdy1dzKTV6ShOm4irsSq8weHsVhri84SmY5UmKXWHRRyVK5T60Lq
bJVpcTUl1OlxNgWyVTTx07Eau9EuIWi1pJ/59v0XHtpcYX0EdyLAftYXczcKSYXm
GOi0RT+coPVCCxGW4hxhBqHCdAb1TP3hypWxquwUB0k25uCYOSuDYpQBfmW+H2hl
yBstfGRUxjiWkQU41z20Ro/oHEg0dCsFbjxCnt8FWHwMiiaVioZTYpA1xeUfh5zC
KhQ33SXFr+NuZ6+ZlWJ6iq8gw1ZgXuK4ih5XEqZH/nwensmfv/OyMc5Ry9Jdzm4l
fmUREGKYPY8JFvJU1MwmdsRZ9SQeyGMqJe37sUoMoxUhjflmgzNRN2eHDmMsCfPc
3qMDfTdUqruQzAoB88ZKdyUs8krn4g1viHTbQ6FSumuU1Jx1U5eNrAcR98/VGwtc
GD5Q7uBNwj5wOIEQ7txHhV+ubbynR6QIFZnpLG9HWNXlwXxJqVWXMuKsCe0fLjkN
e928fTZ6xRDqjEz+E386d79tiqIxNNt4sRXSNsHo4ez+vPSVV55lXv+GGWnpSgWN
UFBSZzuTgTnGraQLGV4cPf/ZjfeAUUdLGm8PY8a7HVapg9XZTb2Yrl3Yr9NMuU7A
5bk7q4hU+NTqgZ9/tZoBQbnm5x2HCLIYSwpFOvD5jx9TSa6VlsPD1E/DKg3t9Hk1
eT8qr4izkUsk+x8jlfT5L67rv2LUDo2w3PURI671clj4FWr5AE87cUpzg3xnae+E
gxW3Tm4Q+BaXmC7MYgpliKjIZ+eJhVpwGGVKG05lnS+KC7mF4xbv5S6Bailv1o6Y
2qxcbtS7dByVLMfKN68MuYVLsKTrHIFAWZIbSNNvhvNXeyKLxqXs+qWvErJBTrt2
lnqPsvzCQVgCwHqXiMByhoCCqA6qWrdDiYAaRU+SGVPRBvgydGcuYgG09BhWZDA9
qG4RErpQw+cU04j56N/hTAdmjZRKGSy57vxsOkauFqDmnU6q8k3e4wH1BzwPlXBJ
RtTEZUxHvG6YDoPd9wHFybj2+qWddFZoi7zJOlznl5uA6qFLlIkSYNudX46TqTDU
CFkAvssiH1vl0nLXQpb3qqj+/ENq1YHlsIigHrb0TA3aomomXpaSAhQbuiwjX4M4
2hRMBfmFliGpSRsLwf49lnQFaSca9elIwypSW2i/f0t/urGBQk2SRSvTBLYimv6l
mCvSPs2L7kgXqujUgif2gFylHvsGZuFcmzxEFaV/fcqbSYg2HO+fLXe3rvQtQUhg
pVtkCtdhc9ujRUbh8Jm5Zb5YuULziaEhZdVufByJaQoJWYVF6XXJrZzKIxXcXPGT
RON4rdwkhYoCxzbFnbX2t3xKXdTbGIkjYdL+tv+66RME5oXq++ABHZXHxr8j8Xk4
`pragma protect end_protected
