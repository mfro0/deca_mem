// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XYmR5iHrAtDfePTXO24y20wQkJJl51GmPnZdWh+VdlZVulCnZP4QLUmiGVYCyAq2
YGswX98QiZjeZLBBAdNTolZvfnEnulga2YUxt2hJTpIQZ3Jb+tM+qQAF6atxb33e
lwidhn33ulBCzMWdfJNeYRUeKRSeLaMQ53t0AOKB3pg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5824)
058ay53WJuYWeEoe6ur9CCfXLfo8Rqo9wVqrpzP80SlAiNu7L43evMDVhqU3FPW7
DmueI9mlR6KPJXLY+c1PsSbGh1J+gDO3y3K5umgd4thv3noqxMx9ZuLUmVZYpY+M
wpFVg5zopcyvuDQhKxxd0rIfq2dpWx09S9LArqxQ6d+o05idRbrNFsvKjI39IBf1
foHcltL3frziAtWZ1IiPB+BpY3zkSq6YEvnVb7KgIFAstOKHOcUH4C0H4KRXayeL
rexOUJm0PJeURzRElAs0wUw0q58dMz0wWmVZC66rgGAi9Vixs3ChvCP4sI36mfgX
VOrcZCBzHkBg80PfnXXYGJWQv5WdV+bUt2hzl+H1tUz+DQvIVVXHldtr+zaaMcRw
VO18483OZVHlNk0fCJaW+MGrsLma0AtlseIKCKv2tCiqOE15Z2PBRvGIoKPshbnz
uv1jvvLU0T1YeXj+uzTKdbkpPcKg09ZB97agx1WtsH7+iOZPZAuKjxKUfbJDjxbn
JQIgyKjOUaQGdqiFtSvLtGElXy9vHyQdZ+nv0ue3dnAqBmAbPvaDnUyo1ILAK6s7
bY4RLJR3BGMrQjanWsN2+kEE0P8u5NRu5iNUJexnWanpAeSgBY7DYpuLpFa7Pke9
RP7PXiCenhdjpPTS2P5KcJRclJyHF2MUBP7M/OADrdV89uINgEBr/CVOql5VwZI8
DYkk3Kvsi3eTIMDdo3u2DHWDPGW6c7TQJOW2jbsed7xXVfO3D9TQQ/rqo5oL/wLn
FQiXA+6csOcmhd+bpK4UEycS39wP3RMLojC+NOZx3TiZOOr5iyI+g8hRKYgN6Ekm
riHmw5dqpV3RqB7Qm3qXZ4eqdigf7dVlZVyq6g94wAZndFvz5r2olC9KHj32RT7c
qIMWOc4ZOEhq9iRCXLezeWUTyPY/ABXPhGw50+DWUS6nZ6+Ql9+7NIZk47+lBKB4
jk8L2Pz5yFiyaxRd6c0Cs+jn/mWTqNma5ubdldcIaeYmDaRyJEMisbccgHHPQOek
lP7e0zVp/tK7vlHFGI/rCqGEReRmKPo1k/QTVE28ozYMzHo9LHAr3d+zIq9Xqmqn
1A3rVIssjFe3CjTfCBQgMAqFpD8AnYkrmIYgazbOTLl4wZZVsl3RKNyrhyl4Lflv
2PQA9dDrbSUb8HkEBQM2wTEosnr9vnUZ8F8S9v929fAEBktEJ1IketNa4HsyAI5d
5yC2ErElnp2Vuz2tlly5Z0q86CtPe6ZFO8cTdZnDuyJ1PHX+SYTZDXGErunb0iEg
pRTs7A780NpNF/VHglzPDZkR1oBS221XWWGqHwGxtv+Oub/nbBACcgGSz/oDvZSq
NgaESgEOkih0iWioNoc7GbdzSbpPvGhSFwlwdnpFowvrVrL+nLeK0Mt1atJGMZti
zp82g8no0Nv+0dWl9UpTFCxWUXejJ9jbVvvFvmsSmPsVQkryusiMZkMFIUTOev0V
l3Z8+ZAZyoSkv4xvDIlHwoy7cT/knWVksL7oCHucZ/542OmrPY2bWKcSxzrwiyQT
oEc2xD5LtF369KtuTiJQRin0UY/Hbia1gsd9BHz3zQSVpnTfD+l5g1tM5O50h1mH
3neDGJVLlqIJJEQheLBZk69wRFu3WoXuMdG5rSfUNPC+Pdl6JNAF/TnF6HLclB6D
RrgZV/3zILuhVz/HRAoZVnEYY0C66Ib7uXejDelCwe6r8MvZAQ9YtN1i+QugF6CL
Xns7rn07mU4C6z7ult/d6MH3+67PUGEfXuyYS5Pb/MuSSpxLRZZwKXB9AncYXiJB
0YIjTaVFfIPIvly5/crvi/ZKbCM2ZUfp293TbVh/gR9AP8R0+b9AcNHUjd6B3jEs
h9kcSboT+lvBj9dnmph518CCH2NzwFOzThdjxAmuj6r2UZvhYbkCuiyEAxJUBJKL
tTJ8YwjlyIo7PcWbUmhjNuFNCXb+926SByYCoA/GTdyn2l6IQYa2Mi9NsThrDHGr
rgQvCMpxoiGIbWODxNbH9X2snulg/NaTuzXeZ6Mkwfbd6AsIvApXNUfPd7k4cPom
J+0Ugo2nkBcqcfxHiTsfeNHfEbDga3a5Fkz5FGBopmYiVgRNOpXNaQeI8A8pKFTT
FFrXKuOLWbjwcrjG5ET+wnBOPBGk9bVc/kAhS6HalqYRbj6OvGwrLtna8vv4ENi2
oubCXlPxAlima73mHRxz7mE+4J18DajWeBKc+1diAIU1mAf24sOF+TkMnGToR6Ez
visy1UNDVA02BzR5XqWrKmMxzmgJMlkfGehxFTUMKiMc70kfBdao+wkQ5U0I1Nd8
+/mOiTxF+EO09kIEXwYoMuCquWbb95FxKKRhGhLo4CrsNSPeMPKLATh1yBGV/zff
m6U1W0bQg/p3zkr0g9XO+m7FgHh9xZB4sgxVNomSJNnyqbYGyb5deQJiN4CzkUaD
jWuR1PDJYYYF5DSrLGfh3Q1R3yHO812HEYcsMb0DHMIF3etF6/srrr1+DF3qLzbG
ynGwqZWkKZJvd0PCVxP8GKk3V4G3ZFpkjdtBLkYW1F9fIlJ5mmMPqlKQU1AR6oIC
f/ssSvpp46zV5Z5/p96BlcaLlk/1YRrD+e7jaWzl3hLrUj/f7dsHjjt0bTTCuMjA
z6SjBk8rS6MjaGIIhc/moL0bUvs3vED2nTgAKzeJbU/s+TyxzF88JCiSgIUzDg7j
sVnEIehTVFcpLXEUczzt/WUsqyzFtwETIWqPTTM4PwzSuqZKzf10TcX/BEaHeBhR
5i+EDvagk7n9j4RzoTg3OBRolRbNMZbt3mC5+G4n3JcYcGSLD92K9uC4IKpODJ3r
S5duSwyP1m8cWMBA3psBkyI1Lg8veXiisTAoN+28jiq1SQd+jdeGExS0vLP9GY0x
PcPQmcSs7Ifa8nhHeeYb2Q1H9YaxV+mDIB4ahjPlj60bPWFAk37N6pYqsb6eT+xb
7BRAKEST+by65Bc/IuNEhsO/qNpxLk0VecHt0x8fkklSSqO/8PFZYoGyHq1tMJfT
0YDTjECglQhzwu8ZypYhbw1PinZQuoPqrDZ1Rwm5fZzO8kEb1mHNVVpYWz3csZx/
8AOZ+4TZaLfMRmP1ZhPAWXREBTsvgwJwQ3Mn/X8WGyv9XBRwKPeq6VvtKe66hl8j
sD9Md/zK7t6fyUcav1CNX+rEhQdS8VBOsnJP4WwO0d4IVAwC516zlX3EB+ApFVYs
kerE1LExin/8n2u3uUbUeZZBPbrBXMczRW240WmhrMIHU1NwPGzPdHPySJOvuN2g
yGMmpcs89brPIDcB7EOCuqkanYBRSAW2OSIQJ7AB2dNbgIG8RZhVklRpIqzvNWpD
GRNpHG61O9ejQ5Z7tu5dGAtAMLvnD8DKK0j+8ZiUbNEDeImMaaoO85MzmDuXKyts
aRyRpmDM87yNH5RKIDVmT0neuyU/uJiYr/sq+0mgQFcsnbTVj2lxz0TAVviBBmqv
SF5+18DySjVoJMAdDxKEWKRS3Dd1F0X53/1JG9cOm0aX8/d4Rha+VlwgBMFBRir6
jdYwBIrew6mhaWWAESfsm9c+N4bYGorq/CgiQtcYDK2PhQggKaodREKP1LrED40l
Saz5LL7bZRixqlFcxV11qJE5stq4F5VjUQR5KrcQ3lvqNAyFWv3eIkElFq114+Rg
DiOT0xeK0F9eDeos/ibkCYcFkjFBg/5YFugIJsy76eVGvOr/cLa3Z9J/HkWqLjMU
/yDierxa7HBluNHnZWwK5ckpiQQo3CkAztIGiOHozl03Mv2pXFEias0/Uv7hS54k
GLod2FjEbWr/fQ77C8LEVpNFbPtTQLlck6xr/e48anivrfugJON0t9TfHC+uro8Y
9lvcL9+fmI20kt6OfUrFIWMzPfJtqA3J44JZ+fGdrs+RPGgI/XQB7hqJL6jOMMPe
+5eF5AUSXX47IbRDN/8OTxoopum867JcShDY79FeUO8YOxCUTTcfFb5Hn9hBmFWr
fPHe2s8c+a41dLM+n3eNMdHGbfR50X2GPFsoBq0lRyN7gfa4/yYZ/OmM1cPr9J2I
K+RU8oElkXoEUArbYITHBQIopJFc3ewTTBxMqlxwXW6JBdHDmd4CqibmoVnjJea4
6uepuU0ZJnDoEINiK+k2W3Wp5KF5yPDBCFsa5p8s1P7pJpAjUMjDOeQOYZlpczF9
gEmA7OYalxYEFv6GSCgh4tjd8REekfj2WVmGKzHx/jWgR2ZCP1mTlLtm7ZN+L7C2
vgd3V2k4qf051Ih8ah3TFrvlUXEiR6yXFFZwZFuSrCqgDs9KgPclv2K5Jv6oRzaz
q5g97VcKJ62mpbq8erKBgduLHg8uUKiPZ8hDm9JqXLX1aDnhVwIutheq7Y6C6K8v
PY+M1cveEbdZHLNmsrL/WRinx1V2ktTRv+TvBYqmE8lk9ap9N7dZtlqq3gFDVSH8
eC6PRoq4q9zjLcz2/cW36TyCxFPA8EEJqvvn4sUBic6pCN5UWi1tzPaC98UAEVm1
647MmgSPaCxqPb4vYgPIky0G9462HE4bENlagEcp0MddSjT9Qf5XSDj8L7kpmoFK
eHOjUSVc5pizWWucKnvLjo35c+bguuIjku9KAxWzwlE+nOUh+tfvLuICfF3FJj9L
hMG8KqOj7dMlMvXF5LkN2x/otUBECIcQT7tjRmUZXAwGYWCjmyLFn9DShyMVYVo5
ZqKQS36McooRLR0xJH5G5hxsww3HnayaSOKrF5C0wFhJJ+QQMc9+daHbu2Hwom7D
oIDM/7F0WrlhCZeJZnR+MEv5ZhMC/Pg9dxStdVE6UmUqU0inpX+E3r6IPJ3ulz0+
TvSwpzMe1dyR4LseQkFrd4ArOoaUbC2IdU6A8vu/N1l71ODYJkeZjtcS+IGAAfFi
52ogKhhZMQV+al7qAC+0NB98oJbUcZwEVs5ZyDcOPDPBegMRbcG746Cz5+ENWDOO
reLrfFAmzzGFtP7TAURkjF9uJnTlT2MTRZQwpFj0SDKVkPBgm17AP6Jol5nh4x9W
httAt0UeRfAgjFkBDiG7E3WuvjlVSJkZbzNFdTAmbIk4fO3pa37X6Sys47yPK5Oq
2XOYmHWiB/W8Mm45+xW4jjS+DqPRJc+IclkeDuuTfYM4HLcsvxKdlEKTc3EhFTKk
gcfoPlZ+Aozlu+9OpfFmFWl21knCbgnrgh5AbEqI4O+mrSHhKwZLw72VYhHsUr50
UWwdB0TLz3Ak0mYGLdDkdOKbj11GyCXBQXg2HYKw6DNg4bNBefXNNBbqMDNnwuEz
orz0Hamw/ckGsQFJjUTvOjGU20aFiFKAGzvw2Z6W6WhoNxQq4GMyp1amyryoK2lY
MAetO5W7ZJHIWaX/fDXFFTfCwzEOYaPBUfitisaxR/fNUjrHE6VFjVWm9jYFWnlh
albpvOkth+8BMQP16UorMtSb3I1Ah339zy9wsZ8tHenzxNq41hXr5vmRLT2yStLQ
DP8cdJUDT9Dik0GmMj/HLuodYFXWVtqHSjyoI3jAaWKWYW+zVlMJ0CR+tX5N4uMO
+15Mr2qkFjDtVdXBmXFF0DWM0Rn/rN7luE5CfUbtUWUuTZNqeeJHI37U2EsbETbg
UjH35tyqHUJeNJinGEzZVAGRYjLVI+/VQbnVIWSplo/HJ33m84STrt76tCOySEiz
oS1jj8g43tKmTBm27SJxjzPLlInGddICUF6ddZ3ZXD/4Yc8jZZ5/V+utzCliB+ix
3c8ZHMW/4whRcfpG6jkrxQ8n6KbJ3fxDCNQ7QcZA05FnIagDxRcSaeio1LCZ2Bri
2uXn4Dx6q1hzuaKYJJHlnnqr30/GEo8VTY9QqhCy1Rq3VPjZhntWfHCRubDzxTQb
BdyPrtahKK1XerWDraEy7u15i1cFzDp/EeXzQCrWULukKlx3Gu45TfRGBu8vUrB/
EGmXsJNU5W0ZBTiF/02DGd37JpJ9FQgyblAvV28faaj1teIXQnPUFFYhx6WFoZNJ
sXXPb3V9AZaaCZXKt+2nR2Yb3vDkuPCNijgdD8QegpI7H0GYhBZyRucwv0hDzRN/
fmS8GVtQCovoZWqyzG4y4EzB5z03e0yRS2Zc7vKIHGIG4rk4Ad4pm9RBegIHj8xy
W/bdYXJMFDVYmeAweBchECrscEnLaSTMIzW/kqNJ6dvesAfn+Dn//503hDoHWD1s
GVUCUMQoUZwmDfjDYMmC2D57MPs2WHB8QO/z6e9EmCk9dJoyxR0OT288t5GgL/Qp
ATbBg4pJg+zn/XBZVPnqIUV6Dh2kfzRrlY1MkJWKU8iVU6VaVhE1uwS5HIlocfMw
VvQEwJvl84XhWkydjHVZusOAicGc1ofFwLb7R7ZopzKPU869KRWZCsBnWUlRWySG
jy0F2Pr/D+hdJb/7j6TRecvvs0EDCZ5u33SPTsSpK2ayJ0hr2rEreuLp6tCQjIVH
NzSIYbpUu0f/l7pMXY7vMF2drMDUEPy7ftEymi6pfpHx1EJvIvipt23eGE8F1kU/
+P68Q8m1wtIqSfoLzCQOPgZiW83bQnFgwKHvHh42o+TxTwaUyY/OcURAcWyxLMm7
TAAEV/mfRL5heFeITdOEuvuBlonJgWFfP2pw2hmb9RvgGlBiL9qCrim9g5ZpeZVH
nTLwbm8oNlAlN3gXoTYMeegIFHzsgKCTgYxNcjhXE3UChyYKmHIypkcRUH5JoOqq
5IkFETr2ceqEdJ8cSUFlqm3IizMgvWvbGdxcvvzcDLI75nUPSIY0NdmwYod1eq0/
w9m8tq5BmJ0qr3XyZFWkFIP6PRLqhkVr0XEBTkzP9Xcgvw6rz5RVIetXwBro76ro
GsYTW+UDPeaL0KjMV2Grezhv2MxgHH26jbx35giAlISbGGs7pvnMpK6hgLwFFeHh
sTnXg5tVTpI1epuZb8I4HRMT3yRXH4YRkEtztfFVfqgPJDVuug8IocXu2Ca3QFDf
Bmdpyy/V7/ZG+Sf2nOougPTVwO2OtXfR7GKoT/XGpkESxnMP3/XMh4UQqq9fL6D1
sX6eP4VhEBJw2CdkYn4i7tBAbs4icB4Rj103CsKgIxt/IN9c5Hv8M3d0zhIZRpia
TTecZDELVHErzOM41GhVfbGBiqEuvQlj4XlXo3/lZp22Rk0opxQidRk8rTp50po2
65PX5qFJXoBOwubVauVo2Gu+r5pEkL95ALYNWonNGDEH1v+Y13owqD9Cp/3cJbdb
e/2FmhX52hP76KGlQCOoF1HjoL6WqoQoxGHgwfS9uwORQ72pOJ0waym3J7SYWXEz
+mKSW5r8BEgbs4AkvE35T+ctxWxrbMDa8zHTs2/gLFmb1i3g3hrj8a8sWAU5GpQD
5hibT6NeMAKWWBAVCzVIFPlL2dp7EMo0oWZ3tzdzti2aNDKiLP7eG0xfDr8PyDDv
wgxYwl5fYxV++GHKP4RaT4dgdRsxaoCeEaq7Ay3+Pjg4OhX9Q92ANMqVZYGO4tC3
RcVqPYIHjRT9NaD89FxyecFfgqmm0z35kSe7Gj3iHOu17axNO336T2poG9z+uUKD
n0ZUpR1wZjt1gjgjDie8+LuHXyWA0+dOCoSTdMjdRN0OlVYJt42UMINGJNxTgZWs
A+/UtMFG1Se/QHOetE88mKltLfauoWio+OEba4rz5spYdp8rXoENo1On937iXZ77
iS1L1ib1E4GF70Zw1+9PEtw9knkqCkFaEOTs8wrZjwuWwnXyOXfcoxLL9+b67m4D
UE37c+O785hrP8BrJqAR+ZyZKNSVrUwhgYdGqgQLMYUAOCDCFTsB/yVEDa/21Smb
HzeBpTO8CIhP4DSiGkQdOQ==
`pragma protect end_protected
