// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
FSZp6TjJ1enlYuzWmHKP+5lGZW5ZaQGLIa2YqNhdQTb02W6Ee4DULQzKWf+r/RRCCvVZDulaoIBm
sSpWDViYjXnglsnm2ymylJDSl/D8LCv0+yWmk8a3XBbnwN3mCSc/IGfNaBuuTJbIm+QGq4CSEgSW
kJujLc/SO5qhxadLw7qzlzJmXXYVDDyKNsbv+yUBYRuA7CfBMhB2a47Vt39qkmaitwpmsASRiPmR
+bbPnw9MGHHF7wtUOaka6Y0kRCAIgzQKGJtlOjwaDM3lrJbBlqA0y/KoK1Litf3LaMx656Ch2yTX
DJSvscINIdqKj+g2K4JBtJdkMiEjQLJLsdMMSg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29408)
QBPIQl5O3IZioojbbEwYN4uTm3PSsTGiD91Q7Ay9+xgX1ztOeiAQidNb/+gPVSAUWIV9U14YptGk
eTxQHVjeKwzMafXJbdu8m5ZGFdu6LoYZ46inr93n30legDG1aa+B/DcEGAPtrAtg2d59TPo9CE/B
F2f6Dhc3GT7P+rPeth1j6f3kt44efWnUVw28cG7POqsQmAJ/F+C00PICm74GN6b4UE9EQ6mF7k8O
/kgChHQa0KBu1lG7+/Yu+RLW1VgmhxuBppGAjmpajDC/AJe3GNNtDEZzTcUQyrgxWxe/5qHMRhdC
JyB/zYs4yXo7FNgd+mbA69xPIVON7y5fE+av4a1nN95mRUtJXSwsf6DzufJTVVZ9AVadwykMUomC
RYmU6WTRQLgderZ1J67C6NbYnq+Ys2Sc/sfiAC87xXCHT3KKvjO9gwTh4zJ6erTCMc3iNHkfUfDd
xDhPiaia7kcVo8BKntrm+i8L/1V/89lXGU7dezx7sj76lBP1GdDM8SsRWVC5cVrTFEXLfuw4XNZc
xXt/bYBebitOrxANbFtT5otwukmScBFBgFiFIu7DwtWALNZbdIp/rQM9vaUYbjc9ILnoxhRXCbTP
eZ/FTMqHKNgMvV55VIobfzgOKyJLZ4btAPcFDsBoX671wTRYvsAyIeJ4LXa0kAVWn238GZTezOPL
TAXwMmKUVxS5jpkfDLtZjguMXNXM+JTVksT2jWYFttXKTZFQghBCp/Xn91tZW4nQl2h0c3jplyTB
lod5UOFEVVFEpgNftNICkoO0JOlI6QOn5qIZftAzECXzui6KNb2RExPTQlD1KRhQsQdJH8Dxlvyq
GxZrIkXziIABnh/1GPHVVU0okj5FDSjWLKwUDT8LeED+FcdG+uw7JQuE4V0yCrfTD0ph2iWxDodh
RufmYfeXNVVJCg7sjrq9V/Axp05z/mlFgujBsUvcZpuC+2H3fHaBiwgWAdNvF2S1XlFNURwcga/G
iRF1ww6mrPCT4PUrRZE7T27guqDbf5SrTrF4Rk1f8HQUe2/ENRM6O9gY+ALU4zKi3OejUTswhty5
EkGyYUo7sGab2ImC+11oX6GiAHFavX25w61zbBQlJUjURyQgWfFI8FHwuuxClTiIKfa4HEP7RQ39
s776Faa8For+J4pzadvcgdhWqqD9Q6AUE9maH2Qn8CNuCQJbm2XKe5+kRce6uLjUg/ZmyUTO6tRG
z5Zoc1fywjW4clYVw+9KD0fhnjKl2ZaBJRJYLuimnWq+sKsa8pU0Ve1Blwp4oEEwnFpQBYLf950u
0j73/Kv3oSi0rECVfvYPTpxj7LpApVUxfGBLjGKrZDx4Xt7mXABcngHydBVWyV+lxyFpTq01QyNB
rXjYwlZluBGliynfE3xS/AWeRsVz1TsxeSVy7mHvjVyzteeg+UQwmCTlh0gnV4DUqAJpcl943Lyn
ZI0CvVPI+xxaQAn1vkR5vpef1L2s3b9wfVNF7wTmSvGIVOmLRp+TLeIawoXbcc4RyBEHnpCJq+Oh
7H0tXaQzQaISDWkpbherk1hMwNo7eY1AUcxzERSnDwo0cO/R0qdgNoDXiXzp/yCLvMjOn+DZe/PT
onWRsT+xpK2DW6B6WiSkSkvuuYq2DrPUSk/UHnpf738mF5l7kjveWtuuTXPXp608PEyVuk0lIMGw
oVynR8xy7sADaZx/A+nCQe4xK+WISwkg4yE6gG5OvrJi/RolDH0GRIN5udMhDnW3uZSvUOYWr/dE
DUfheTsZhIQJN80RE3qgvqlBqP7NTu2gTrA67BNQXOxp3TYkyKZhqDoGY27/fo8+54Y6pVJrJGd0
tHpisyz2bDfeymmJhzY3JCia9Eemb87GfG1lXxU2tVFrlLGztthALGXSljHRpvkMyHBCzNSpNkcv
/c84lYR/gu3BTxUWvavi6pBhGxOlY2gZtbW5iMRCQx6J1S0e7Nm1gMZIE5F1qYhi7cDN6/xBXgC4
awj8aFrjo9tWtQES/C2IESKLvpItzn2e6v0D7pyd5rPbM2PJBj8iLHF4/HMA7GTSBiwbP6C3Ipv5
lP1QvIPBVf5JneqfCcZdzw1GH52IgAhOToUKxk+IHOLxkPAVLnSuf7ZyPPkkZi4Sj5ITL8Nlo7YM
5jUXgQAZHPPoyULDcHvU78jI4hRxasT2rQnJA1PeiqlCIAfOq9gC2uvsPqUkXQi8P5yW+YYyJNak
AsCci0ID/1zDVgf2BK7eFcrkWFGlI96bo0QuOCbiYz1C4pPFycuhGq3Od8mVtwsnr6Zy9gEsPROm
VqQYaaeKF58RhfJq4GxirQZSEZGYwyh4k7CgVAHu1zr2zGHXDCyhD6FjFND0U9VNe16lajewSj/v
of4oMLUUTJZcpiSR0XyievJCLmbnDPXam8+yj4sJuM8hsj14hgN56kwO1crUgUJSN0znZOJ7Hvyw
N0Ah6JwZGCr2BfZ8gRLc9srtSPiIQiNixQIUTMSU8nA2DBp/p9XWFvOibMdsKQSRzkaSPBt1PYL3
3xXvTfT+89oM0dSWl2xcJhQ939btLGdWYvFJwGyAAU0zCmi+VuhCt52+bcaGc1PEOSf8pbg9UTz3
1LXOfIDZvnbCvbQiO2ugo7jq2aRZ7xg6TYTKveSf3CH4nu1dM2Rc4af7oS+voKKrlBrvDx0JypcZ
4nZBn8wuC+DURJMd8Vx+jqGaeTJJHySBJJEsGKggcVAsNvuPYONI9G/G/RYnXU+xRwyv0oQAMde0
BcjKVebIeUp8hhOYA06ieQJW9P4rcKJUyeMxFqY9p16ZkZ4V5jWeJjPh4zLNKax0e+YFc6nCkZl6
8P080LwngGP8UoJM7E6KKY/W15d7HF+6OZ9F8Zxk7aI8BkZBW5sI3qPIuqo/W6BwW/SnSg0kAHQp
yjVN2D8CDRgXgYSNSA8SmcXeEmV4nOzaxKTrnKBDl4W1Ja5l1h9YTOkR8ObcdJIgugbWehranDa5
lT69f6RRZZGYx8K/AC15tpZyOTuvz0caME6f/xhvfCZJnCSYZ1GU1JMhtXmcsajY4oym8DG1YCFX
xR+CdkfqWNd6xzgafbXSvgdWPEE0hLyzgJzPIbu/fNm9PV2kobnfMuHuXKi4YI39OlDm366VGDkt
sgT5IbRV+Bs0MXzeQZ7gKdFZg/xN8yQMNZffM8tWYjb+Zy1ljwzypYZo/IsYdkcc5sc+IJI+qO9+
F21fwweVBWOjxD0WpZjQtSR1kOZgqo0u3YBUy1XPT7RBBeNOxNy+Pu+SUmk9pCe70bednMB6lL/G
MExwahXYd14INcw8/XFRILMpr+a2m+RcC34KRYUmttdxtD1OzHzykCMFgktg6Y8FmWmy6TcAdKSc
YVxAG/pgFBvCHffboHGh/EOxjR/N0CRGNJi+8+j80D+hR+tLDDGSaFuvdXCjIimrVHlqNeHbo8nD
0nWfgWHsXU3qmp8qohBid/3iCBsnFRJk8Q8uvJaPJnr0iauCI6n7dYUoOE3C530/umFcathx6U7e
vLWecr5xn4CBuPMKeSArvSbmVZP34yO22YIDZWf/yzIx2u8A08yQTX2n9/tJcUpgLSi+fUaRIDht
ybCS/yGrNyWrLtgxqE3PRl0vxilpx21q6zSZWdnmc60vdKUWrX07fihvJEp2m6Ep5gThZ4F/gzlT
V0EnRWIPHHsOsAdHC36du/pQhPK9bGBkwI2SRkRTuAXLfuxqUIl1Q2Ybfe2vX9BEOUx6OcrDez84
jyndIpeEIGwWwqO9UZ46Wx/8lZMYK588nEuP8YbpkPUhNHA+OXmv2GUyEdreVxhfAqnHHr4dAXjL
RKH/Qgh+BXHu4q5f7uYbSqOq08ngh3nPQbAENFPvckpfgZNhec127cdLtbFSN0tmGxZQT5ZilthX
by4Oa0zRmvnEkabJ5rPoTT3RzHOwu45tZ3aYf12iXWqTsySqMj0zjV2sPWfoQp00EQPe/szD9Ux5
CNPNTagHYWQokB3iiuEBOZpoaHJ+CZEsFaeNF5iZWPiF4mkpQc2rS/H3de7pR/h9Dnz5vBqVzHA6
maK9JADjzEP2gvRBusxHL82SlPlsYfmusGh26Y/i9MA7YuuhnH/uz1wG1zSMaEyNmJapCsvTcZP5
PX8iRWBXcbk/Gyas1Jr67H0m6Uv3yeZrmSWXCKQWd6RKBjRb88iotMSnk5zr5jVltnZONgpN7Y4V
rtXCkW5foABnxJPzzo1fk/wDfSBMHXkK91AiuT+G4ltHd5y/2lE7rLg/2QqPIeVz5tmKSok/Bj4l
2z/rFSVswPVsrlmyxl/FQQNZpuIwG83E5A0CDzMUAiG2jKsn4r2lzkd5mwFcAP8J3mAXrMxUVC0v
cwSL1OWQb9YHuUO/VPKsssW+TcyShNgUZG6Yv9m/EoZK50MKJgRxHtpq5/oLmeacyOLrvf1DzC6Q
IdeWJVsTaEranJrg06jWOX8JhlUjzDS4vy8t6dtSY4tHBDgmPSnna3D1zkfSTKhoRPf8kgxH+HLk
lNBuoUMGB3gFiUgEJUc7nGUv/y2GvdOn6XYCa5wmhT8RNQ2m6+Hm1u3IGsjleoCSB89v6kgfS9xc
xRu73qJtmpMleZhTKAcRL1k1hXT4wzO1DUy8Ow5x8GXgsjq1L4jQqT6MpKMiYxM4GCNUHZ2f62Pn
J65iZx3C/6Pr2UoTX4CZB9eJFo/CUIqX3mmUu6QsBU4K3ZQl3L6toE1GUHAdNXsT091zsv7Mk5F3
tAXXsm5YTxGzOmYTb2dHqFzpbzc8nQgkAYqtdv1fzgTy/4DtyXXd7SvCBmS0YXeo0jSnKzdLmj5J
zBwUt6VjGiLMgKDi4qaRgFwYXMPQeev4Z04y6mUbsxIJYbGBqgGxR390ZmVToVdku4kuoVgsNZ0h
2YKEKr5tRU7aHeWuTcGkAj47D0VEcMb6/6uxeSrlYSUfiIIB2FA9FtClTK0AhjuI6xqbR66Qh7Tg
eASAKU2jp7HmnWutcAgNvmty6tRlBVG8Ed+3ksd5ybs+gBkfYzd3w/rsX8T5ya596f/tK1U0PW7E
epK7STzXeUZVf1ZwdoCkG8VjiHKFNwPthpxa9AiITCddHgXtqRv4xnXYpADE6y0Cu/P+upnL9Hc8
0/tV7HH6vuvvFkqi5Y1pRGgiXMAmEeR3EAmB1IxHoZkFNjUSL6Zw9sDv4hI0kqbcEP2TJ6o2J5uZ
9wv6PhPQuJ9ChPNZQ92Q0tPsvzbb3XoTD2KXmgjuH8tkSz0tpzjXmqgPCn3unRtuXuNCg2y9nKoM
YFHLUbCi2xw928nua5SF3U2Ypro3yLvA4ifrSRCxvSYWKPOSIWhwpJZYLNI8mK3Hb5MbU5w6T6zT
t16Xi2OHHxNmRX2FUZi40crvDRDV3jUkthruObhxXiwfpdv37GQS2OznV6YAbLhixhYTnn8hQ48B
n3u/GVm2kYOSW4hG+n/0mgRKQvkXu78BipkWesLB7PzyAbwOFWqgs53R9hJ3L7pyK8leXjiLAZ+0
0KWgabi5KC5twyYPmNe+Le1minEe4kuJ+dGT7bL0WvlLCcExpm4+nkmuHSb5nQQYGhL3Jb7ZRfIt
gT+Ya/7tfPT/aMHmlUqxBN+JUpeD+DJx387I6iDKo7sQlU6jhlSUiepFNhAckQJniiM1KNvQ69e7
XcAhRIQY/sia3Wn1dmXrKkmzTjPTHLhmsI1+9VEctJCYqM1i6DQzif+/RxW+4mUFjQuWWDF22c5T
t7o61S8dkNTMaRB3bgtQ3OPIzKq7+gJb0C6FIRp4f7pZ/qmclnmx5uOtTM815flhvExmhwowKZUp
+YxP2mtO+dsRb5rNpy3c0PyvybdeBedu7a2vWVuJWCH6lWZyUOGDmRtb//aIIwbVwEcNISaRGfpm
7NXOKY4tw/Ca6iCEZSRN7IvRRA46gcmIWgIqTBqx8vRqH6JLLqLktWcImt1ZqH+ph3jQRUSdxu9o
GI7ETA2K2l3eZpGOqcAXjJDmzcUwGIOpg5PJz+cxLXQvj2xMDq1My5slOqvCrsiz9s9x5iJEYFm5
e6RQv7wwut9FsCpRVMRI+ffhRy910DMTbLmMAsEgp/xSHbaC5RrWDk3ztn/Bhuv4dTRGO5zUFqTr
87jdl5wf1p3AWnO80Wy4CMW9Mh+TYrrybTiZ+h0O04hzm2iTuPIiH2JDQxT7TTp8Bw7OwqHMu6aY
sqdCxef91Zm9sXVpwYRWg07C4EzCXqfCO1H4Bs+rfC538jDY+y5G63mfSq9ycGyeNzgrEkfHcBdT
BwBxPr5/Fl5rBNrWSGwvwS2n/3CvVRZXJWfFS0VQQbx9x21G78uDDdvLovcm51KhPrlCalCpJZ/C
g1lTMKGmZeRY7HJc+8icFvJbtlNd+DtwPIBNNQncajuo5OWRuQEsPIiTCIXw2ISuMr69Ttst2u/a
NBVH6KSrANiIlAEtU+HusC2bRIPU5PcSLcpqcaCIXxk59Neo963g0zebo7Vhk8KLot0w2SDPODcc
gEIEOL4Yr5nxjBpyN6P8In3DnH4LEIKq07eTH7ZeLgSHyKqfxDkZXvkE99aO+lFF9D2pxC5+FC5d
ESZcpBkG9lnXIt+ALniDEO8EamebR5pD7xXUXP1IrWBxEIZm9ElOiYrbkjdaQdwfbdhwHvxeEGbR
am/Len8/LVqzbT5mzg5ElboH84Uv/gio69Kkd7LEae6RQnhb9rM5WeKqU2nfCHntdYVaH0UbcRP/
FKSGhZKWOdGv76tyZgQ6sDbow/ZwYk4lebxpAfjQGjQ0cQK4pUql3xxuQ7IIA+mMHP9zYLW86YmH
GfX0VIpv0+K+a6gfXlHzu0kC4shyMOLnP7ZjCJuV2dP9zrd6MJFc0VoLG3Djq8H+JabeztFbKaW+
Ah2jfsY9BxW4zBCftr6RyQFBTccGZjRGOjgGTqc8rAQkQSUYkk7StuGYFcYar7CzxRL/U+vNnIQR
Rr8loJ2hwnlK9On8CsCDyU3u+MHwfoP7uNarz9aPKVQ5uVuncxHGE7UG1zGwnTHy6W432e4P9C1v
n9CNwk6axZFYeawX9H7H6Vq1dLUuoTcfyap8m6198dnjl9rjuGdWQWiXtNb1w6LnlQf2kRnfkIcj
zu1SO9c84eMXwwZKjVBZoRU1qZjMMeOfxcPLUqcmNQBDfOR3iX/j2RyWlhVK9aQM8kwait43orZk
lesVw9WfcbRif478cu8IS0LT0YMB8vgLW3etyc1EUnEPhVmEXZrFbJfKIKsSOXMtGOQPd655bpMd
Sv5N4JD0ogKuOPO6dbxvtBwnwxRRs5Zb2mBH1Brl232gkuW1jE8fgwVFcGJk61iFp8pjcXV1uSbm
3jAvnWlXqU8dNzWhIhKJ4nQSxigA4CSrST9wz+TXesRXyf/7qHZrE57M4ekM/dZsZ7omuJD2VVgx
NmgspVY7fWxSJ2VVgZlgkkW8Kko2mxBLlEdBKTQzulG1TmeX3j6ekUsfwPTE9dn6yhELkCOXuEaC
FZU0lWqCu4a4gYQrYzyUaO3JVlOwRdJRbiftymAXGom6I2E3z8CPk685hwyLcw1t3+VVZX3xlcu/
dsUzijS+4CJSPSonWV6TotUC3VbEbHTIcdLsuqDm6I0LjGRkVpDgKlPsnlrX8M45F1USiaxABrLU
uvbXLLWo/n05ld7CD21IPa3hbfmycAUHFn6p3nm2nkBaXWaJEoFb++Z97BfWfri8leM3hCLLDDhB
1CUOzrBEusjHVg24a27g+m4Vj/nFJpRMilHQd9d00Bj4w74DAZGx4jWy9GIcaUDJwEgpCbx8XUkk
VfbrkFIStkXJ0H/c6V3AdzEudYR0Y5EO4+Gl26Z4lXDRXN8n5rQhywR/Eqczt0d1o9V1SaJsu9F+
S5UQulSEcXbp6qfv4+wqeuaUCci+GL1miUQ9BZUVXpEWUrIU2u8AyNHUO3biB6EJIc1S2xRfp+Pn
6LuEUgv4RtLy7HC9ohnnEGwPe6s+utOClSSz/2L27/mn0EC3BCQb5BhkUMT4OhQMQxcQ+MlSMO4C
rWowqg7x7gvFZcqSnhf0Yk1uvrByGuwx3v+ABpYP2o3EohiHUlRFGQhFfjGKYtaid+UPP6OHYi0f
QUqFXKtU5vWcetwHIJKGNDVbA8RvmrUaOyAK7Vr+ujfI+zJ9erxZ+xL1tu6AEsOKaHHXZ3pMFnVr
HVwhTzZE50wAvDwt6Z3ZZXZUDDplYkFsbOYcH38FTAuoOFLgbfWCa8xGD+zliOUSd9WA9HhLAm/V
eOOiOhFIP7IlNcBxjIjwNIp/0WDDFlD3xrpyqBRqu3asCrLEHv0Oy+549am5oSNmoD/scMVbGh2Q
gLLeyquVtZs+uVSroTLV4idATFxmbqkQQC9DhXEVaMztDhWIMLrx4VHrOgMpsGu/JDUubr73kW1k
TqSlRJudW2hn07QNRgt6kBmILenBxGMOYWpdNGWDVROA6933CLRqaxfNMeVKPuQt/nekjhy+7tFz
DCvXiena3JJpAZRgn1fYRX0f6sBCmyZ1EEo86ATyBIUTDQ4c4tqjiGHXQE7+P12FCBVfO/zN5Z84
6md+nxvuAV14IsobvAS2Olzs4nKZQwt5vvoUbZroh9/C0pCCm9+DwZF/hZcJvQTC3c/IFv5xgauq
JYuvu+TlEJcwmaieuwA4qk82I+1RWTWeW1v/QTY6rNqXQPlkVhNGHwxiYUdAZy9CNknPSP9yZHXp
GZQoCcGVqXapfBNJr6kxha6cr4EZoBb6bsnyxDJ1KUEmUlnItzVfeTApg2052ruVZG2A/tPuyg3N
EGkcuBzYnnm3axxlYZme7ahAKl4UU5U6L47332d7XNLk+omx84a7VYOl4xSmD5xmThSrfgKxQmiH
Ro2mqwbSgFPApNjBmq05bZT3bfn9WVmZk0O9qX3jJVObaYx9paSt+o3gXRid2q91pXce1Xbs521q
Zveu1oQ1SNenhSsLr4zmgTx03t7ccs6yH5PPtiYZSlaRGU9StZcMVTYCFiyrk7Pl4SBM9nNLxmXZ
0T/HUEYlRmdV75tHXaMRYlXpLao5DYrQvgpC8rHOYpcuK9mkU1LANCWqbOCsYWEXk+cbu4Jn6sde
rWWqDycLsPKuIFTMp4ZZGxmBLu8kqKGgG/SuqWzrOGFN58gl52pOuWpv0bVXQ8JjNwmhFo4fY4Ca
U8Z1PxUA5ekQy16mnkBZFX16NUZAZM47Of88L6pheQBhH9z5kybNIrrLdB5ZbNxqFsO7OBi5ljqN
4IatiVPTNnM7IR49jLBsd5aF0zxnXxxwcGf6WVQvkWdDsnDLXxRuHPp9ShBxkWg2JnknNjCL1UBj
NTOqa1ExrqTXb9oPEe9iBI5iV4gCty2nYyuXNtPkWJH5DENome8+yRUzV/XTNLjut+c/j40xAbTp
LYvMMpmpWN5kHVQ2uGiNeGn/7uxxR8nydH8gu6zEOyhATd6wP4iEl34bAp0VB9PhFgucvQtzGff+
+2K5N3+DPDcQ52dFYDZ3ElcEXZ883GYG8TxymZTroq5KlpuhgBedCZhiwJAWAs0JfsMn5UP+F8HH
tvRGU4VfSISZG6T6/59n/h+bjFzeCBdkDpkTrZ7R1DpCjmQXMYnYVqReKww/cica5+Ltx+r1MTpn
nNvFESxoUoFePhuf0TcAwbJH35ErczaFImspFq+nySf6vZH3YVQcIKbKoBvkiHjpH1w74tpV1/Vs
5lDrEidsgSr+jvc66Mxu5xGjwDNRK2fuIOZVfw1S3p4mMwsNvYHc53913RU7CQ/++LZuGjURZmOq
BQiSuKAuTlQZZaMXQpbMOfMPEqedzzFgWLR5PUoBxu1j/xRROz+M6chZwMi9U/ThfEJ5GB15Kk7y
bQLKpDzXk04zVFpMyPYM+W1+YC9If14orDTd09/xUb2vXTj9/NyTn6psTzfxNRDqO4hEPGW/C9Ez
KRlAZyCIG1/Kma0LrnNwWAtjBDn7Vl8n37vQSpBAHvYiKd00zGaAriQOdPUNbAN7VGiAM8IYzQ+y
3KPZ70qmHlv00IQmMgEA7AP+7X4Qg8dLaoZtU742cXNSlyUiN86XvU8esbnqft9WAB730CNdedwA
F8cFezQKV76gfl/R0rDXHbICSDdYBDbKvtFuIMFTa7k8lIByAifZkaIKdnYacys1+XUu3PfHI8Mh
moAT9KnfcWb2uN8nU6JovAJWe/qGuRj18wHiJL5sJqluQ/62DjUGyWyj8Kqak/UZtpTW7TRiBTT7
s+EMhwt9qwUtXgxewpPYdgsuS3q81vE6uPWLjM3HePUBEXjkcnAUH7l6xoo2oO5tEhIfvM2BJ/BB
RZXpXfOWoakoejsg4tapU6a38Wq7L/4K0lGl3SL/9I68c2otydTPUy3kn4dIXqeJRUD2TSaFVlaq
DaJNZMye/Y4o4LNLiKf2DUIF/qBzoplbZtGUPJt0jNZpiFcinsbSO8BDXTLL+A+LWisKCj/McwPc
VSQlGIKJbaRywKNuNDd5C84GSx/31jfMsjS0vFv8F86TIlB/w2EhN4RwO7XXwBhxYTEe7NdcibHT
cKmc38bvIiQfV9jK3OYDy2IS43rLSE+0wSp1Kg8NPV65/3tNoPWEo54a10cIWTtjwfrpDtndAUQR
QGTRXK9G/gAxsS4aHnRZKynIbWj0Wfq2OLcA+jgo0LuTvHAQr0jXpT517guG3VsDRv9icnkbb25q
LwWm2NbyEXPdo64UHNVbbtJOlQzXsMVcx5If4ei8rdDR4iAO1fAARWboyBjZPikkSfleldxN5k2h
TqJblpVm17i8epqhN5nnupc1T4sSxvL39oFJUfgLBwk2PEY3hwBpUTj1GU60duVh9A05oc42nD9a
DAw/j8gOgNAFpoc0goYlDxGT/NVEiDmkC9/3F2K42p+hIuXT2RIvJqF8m4nt2DgqmdXSb8OyojtB
qXdKXp2Fo0UCEfxFUlwvliMLNPa87Tq28YkQOxHf0Zrft0kenFGf5o+1nvWLI+4FEwjpzCF1+5+L
2feYICMKdhCXuxG3j4wjWzaeTfz5m3otGu4mCbIQJOR5pfG7mvlFWQTPx00rxZbMtJfPU1RAOkJi
Q+cWmLfTiAQ1bESwg+0zKNRfSsjm7WpJQJf83abg2C62ATCdtgRlOqFke96SmO5EwIH4o5B1oSYm
c+dxSelMZVn8Xpl69TMLO6NiuQ8PnGNYoI/YIaSa0XUnMjQ/+tQFzmLawkr7o7x0KXD1SYTsdiLJ
mMxV4D7+9h+onBd55jy3R3oAFPmeobxZa8BCYuJWFCdwzJoKG0hPgjmygdPsdwOCU2i0XOamvTzl
f4JxFtqOqEq1Qr21eyDA+B/65yZBmlqNCDgzB/aMoJSe6CW2t2XetOb+EO1V9oZroUvwInKQKXj+
DdmbgP7sGGjmEdM8HdCB6h7tYnpaGr2Vg1G0jVNJudscfzziDvGzjPlOjzaOJ85EEdkDvMCz7adY
s36Z9zPyXMqGCWt/ZYzwL5xZvr3P7GhlrJqeX8IsOtjgjBhBN/L3AoEUO/pONukThUTkG7yfkUi6
+1iZ5mIxHtD++JViImWSZHQxAzMJ7zfTuRit7hOSg64gBc6JQ01Pe4k8R5dxPWGDnFUpKTyvC5ub
7t41EeUhKwW8S2+v4i6uaRj4leGfJLIiD9BXGakGahFQebNaWGax38WS46/8kBzASghBNBDfGElr
UFXhyXLTwNoiMcAMuUikcFlJw+uLnqHQPMuana6NAdCZznEzfBsJqEz2u/yul0+iUrTnddPA4wRA
LmNRU/O3ad0muJ5T4o0cFKi1uGUkq3ZVzLvzUPH3by7R+/vlY6ecufMbp9HazIfaGltotex7TcxA
cokCWVRk1nS05aauNdM80aFcrWbJRNx5lwQHEX/PKD/QJBwmpPAMWv8YXSfRoWRWQcmubPeAgTy2
Oh1ucR8RUnAmx2EE6Zxik+YYW4kQFdy4pkNSLNfVqtoRiFZxIzRlN4r4Yv56NTYEkYLB8iNJbHcS
AEKYDh0ZqSIK+VBMdicHQCUg3XLNVz6MywtZJAYZb2DOoD3BXOpcDqiYo9D54vxiTCmPUdpX036q
5oaxVSvcRYoB2CDO/DXze7rWbN1yJOBw4LtipHewQW/48MAJC+tKMMUlITsaeHnQOjFQjFFI4AY3
YTcrHxPParRNl+aAOycZNaEDOZdaLO0fOg7BOdwRZ9gJCuPiMngO2LizyCXe+vB6cmODvvtYL0KO
ujgFhKfXhgfK6FWTifaCoOHMWz/3NUX04draDgRrVxYF+iy+dxEVuo7fykBPq8BXgFYUNLEiaF3E
9Us2WMPm4b9JnSdxMYZCSkxF8JyCwkOogLX9dCgnBoa0E1wK/ZaBLT67NBlOcsL2v6sZSMjmRNmN
WqZ7t0VWoApWoZK3bj0J4Kiu6iEk2hBlGaWu/j0byS1OQI8rAB7F8TAPVcR/QdHSeq4X7OKybrKc
N6vNworgHo3WMGHIsfcTptjrvvollXMtZjrw8vFWseFMWhuCYcLn4MXp9TeJFADaHBBnmmhAERhH
eqRDwJOZhZO4GWXeVnWplAc3/UVwfgj/SpCA0dADGBeGj81B4f+3XBh0JRkdyVf312z2HwOvwFKl
+VIbpSPaXVQQH6jxguVoal45Enz2ymtrQ/eMaIILfsTKyUJjRSZgkl68dngTEBQOoLFvwsdmEhCl
0m9WO+E+tywX87VX/VU6b+TkOFPf8PrfpQ6GKJ/0BypOTCG4tnWlppD7n++7TK/L60PksAP8t//5
TeQR5YV3xRicMFqRPARoc867KYfuXdUROip5tqPy4X2vWVgB9DztHRWAN3no/072g+7oEjczWjr4
BnRXE+5XrgHBUMTNnOCYOmz3+p1CP9o2UQqDUZyevmRF7qdBQQJ9iM4KCsfVvvlR2Ua1MqskM+hs
JRW1AID8zruEbD8hok+fHhfhxlYvxnv+axedmpmjOnavAj5835ynCTH7MfTxZBlXJMXYK0PYj4io
pD9jPOuPwJ7lY6GkMldttWqTxyFLN+/yzNAglPv2siPZfWBVNqa/VOYnQi5+NcoolakuwxtpRbDG
v1Tme1jEXQiL86K34rRZ82cz/dMaiZBOAGM8Dxu5UTfLKGTKc1RzmRRqlM87QGsyzi6/03VeucN+
+TtX3iBRkKpAqQg2UpG7V9BbgcIBNta8mVXU6BW5r5POsRwZwuwrL0GG7tpgG/sIgw2AauFiTJdu
2Ie93vkRh61FHGYIu2kP99at8Iza0zOb2J6eiHLY7jkfZ5G9wFfTeLIvvBcTjnCAeVzFv1ReY+TS
QNosba8w6Q20fktMA76iEt0RLmUPukajT0T1QkJsDqnQm+crFG+8oFzKDQ4HZxCcpHuAHqQOvYRk
/V2OtPnobUgyIYZkw6c58Dw3M7U2E/sn/pQIRbiCie7zfvotx23ST6ZujcEeukWvcZ9Ch+BjyMef
RIKZne1terWORr17gm2X2vOrbvnjaeFemzYejJkdLVfIT7HQc3A5yDc124jv9so/IV4zbOlSfIZA
NyRSwGbZFxUrFzRhBpglXX0IH55Wwfzu8k61hveHhVo/oOhe+zpZ21sPUE38G0CRKkdN4TWPfVmZ
CjBHtC0uVpyVuScZPKylu0SfsgmwHid33fii7wK0M/v1xXtc7vnMa/FQiOsTuIuUdrQ9YVSZAt88
G7IK6mTlhKryJ6vE46mCegy+DZzdFJa9VSSNs7bAOXahChYq6j6WoTfrSL1YY/G8oQyQu7AoZr6U
5ng86xFEZHHyPrJmWH4YOTNLyq9l1dXImp8jh8+lrDQHInCEngBIh4GOHvlP/0Bd3ob+Ak4RLO0K
JT3g4/o9OqZXW7G62QSZ7LW9qcbQ5tCTs2c6MqkiI5Jumt3JLn5kfv3PNf1P4YCTAyp+G5G2RXqH
58V6UV5IdOHv5NBhrWn6bBI6Du2IG4QAUmZ306YzQB/x8dkDde5/XiPir3aikFIpaR/omKJ/rqKu
qGeEjIVNnNUuvq3l7w06MlhnsE+BnQNNgll0J79hHJEoIUZgCTCThqTm3+S0dCyr8vmt/GDgjjAx
9g3K9ANggz1QHjx7hcs+vroEr5dsbbWzE/Wtvkk29P9vZbzY01nWQ3ep8/Q0vcNGPfS3RiIaxy2o
k474bSHpzJPiCq+O0REfufUOXOwTcjGwMkT9xyPgj/ZWpzw8gsOdWmgjCLj54ZjQwV9QOS9FawJ1
hyuLSe8hmd+zazJBTQzWHr0qtF8/4rwYOT6wSfFUOSNmbHBOJHQWY7WUUyHD9nOKHEJOs3yvbU7K
8A00WTEP/hGknVNTjYeI3NKlI90PompvrLKgXxOsp9N4T7as4Oy2oDzPPbghZho9ZcnMrmTf1GLg
lJKG/fabxRNURmvxxaBxmBtpDXf4Ous/sCwgeoFgTkuU61mhtME5UGhpPwWa8H4TQe2AdbkdXToJ
OpAKvjg6yF8y0BCLe8xwkT/p/iTWKHyaHGMeLvF7/H6dX737cVFmLtNYLln1Nj85cnpNNaAwdzWq
66u4YJ3MKABtlMn2+Z07jexCKaAt49mLYIpb672vqg4QA6g6JiOKPxQ32bVfKfpdVTCrpGnQERiC
0m6GRyXEp6NuUR8P0AftRuSONfn4YJw0b0SyCVzxcyi7Ap5uoaGprn/ENCrNjVz1BZwtp9pI2GPV
XSKcP4kjd7j2az5w18A640KdqNoTCiQL11spQ53P/ZegCZdlyX4sfWiuXBAdqcMBLeIeOrk5mTQ8
JXPwuX5wsPwm/L91JyUxw/7P8tWmAlUaPXEMh3Kfz8FKfOqftpFeILGYRSpgt9fWN51rSEIr82tW
sTqkfQSTU2kyaOKpyhmVYiC4ElX3oIyXq59Nal1INVxKbeAzCwgLEYHdvbp83/iZ3yA13DGgq+/x
V1VxVdljZ7t2ZXsOl/MzYQdvuVrQ4YXil1+Q2N/6UPlydtWRuaFSIUcyc+4U5rzo2XkfwiyBpLlr
SoH9nudCBQLuyIEFi0ARg37kHchjELlQzeLiovZOPs3ikuAgarNdCYwNVnicSvG90NG/3ThiSEmc
J2TiQhlzhu8EIfN8Z3PTHQyG8+6d2aCcJ5Lbju8wKMnsAjhUnZDdHW+eV1hNoIrXHOzo4STWETGk
9Tx4WQ8bSsGffAjRSU9EwgE/MqRVQe6BT3loZSMlxmisuz8JheKjGUzYbdV1aKZUUwYXbWG+DWu/
FelkYb+QhmB87aYVAU9PT+OL3bk8WybC2TW70Xvt9l3wFgfagrLPOR5Bay72VS7K2sKwkODEPf+M
bAW+wJsgDOmRRqluFcLC8+f2odJstsOBpuGiBDb0mB29hsNFCl9rAkoVvFt5TBWfHHQM6m/m7SYJ
f6lNaHD1WzdYL1s1Dm4mqSpLfMjjCS7VG21IosPXSi15+g0fNXSHKm4bxT5ho5aiP3IUZtWENb9G
t47Dz97nvJVl4/H8FUcB0to/msRJ/Lq80OUUjMLxjiD21igViFqaT7H9XhricKk5WSq65Ho0FPgd
I/cuqymejjYRmAjFq57gCEWOEeFLIMeGZ4iS69VWwfDFo1hG0qy3MBTcIxz5FHEPdII2eHAfExjh
3vGJrXkafVKpyeaLmiuuYixh+t6LHDoMcDF31EwhLwjyDnlTUNVL++sYhfClb7FSfmm+vr+rhL5x
9E0QQElsAD0ubu+AFNsAgLSRZa/Ij2Vz6FtqKc8j4e6WN9KrLae2XwYjcPV80E51Qbe2G9jgWRcz
odB7+CqqTZVLdxFSRteMUEMYv5BvRSH/vkLe9vAThIFfy1eUs6TVLEUzu2IJ3Cp9o2MNtrm4B+NY
4jSJQLnfKvz3UkuIf1Bn4ORkU7L571z+X8mRK1r+EOC2LOAUBpIm9FaX8aG4vqMm2hdMEh3HYdnW
Sqli8EScj8fcxx1sg8brzPg7zPXNY9PW7iWs0t5jfCHodvCzVcb+PkyDX+VMpgvwTRo57IFVjBvh
K1u+BmLjOZRmtaXMs7GXtYHriTFbCZgUgnyJH04yvZhlu1ZU/3wWSHy37eDaZ00bxCobf7mE+9WF
L3VwvsrWrkCAey18jCGX6zaojrt9HYRR/WxJ5uUHd7iqljCph0mQYgqg2y6kgT/VsTX3gGsm8h72
rUKX61CkGwNlNZ2uiRU/RtWFm1VbYtMThOeqfhNbw3XJoQLNS0nA+zeFyiSrSs3c+rV3+h+svMJ9
/153Io/YwuAIFeSt9taKDQrCLY08LJBZoKD13PpAEfDCju5OWHZPw28jk+7QUcdfe7kc5a9FuoFb
lZsxMCdSJuu5fX7oF+CZrYEg1Wog4W1fkT2HHTQuV32LuRekLGGOf0WIFmeoE3PEVU/KdLgA/Utw
yWxmzVU45Ay0QsIwh0Mu+tL6fANlItd71XZAY/dMeKhxAyk09QcHOtngElHlJN5b9PfYhbZ/AsMM
+LHB1WhREBST0tqVEHYMjTVkmnm/ieSkonaBMTQxzfrqSWGyqOF4hszcnr/RN4R6m42GKNIWnsTp
m5D1JjUn5nfG6eAeq2XPwowVSRoJtbWP1XaWXsixidF/h7HtbaZoSLiCo0Thz8OgjSKQf7OmrP2r
Zz2EuNTQNP5yiqhgM7Ogdj+CjjfA1NjJH1ElYryrAvFnm5BwI6e6WrTydZzdsmFhwYbtRplW7qWV
HSMUz9Mps1kofesDPLb06ut8VVZSFbhOUnSzUB6L+6qbDvuWv+Tq16TiYxBoXjjKxdAXwBdNtMjH
WaHpmFkJnjhoZiULsaGGP030P2KUMaViQSk6MQCyzZipTJ/GwaRd5oZCcBi/fUAXezinMBdWfSm9
pPeJIjfm0uzzQJ+ip/ou6LDFtaCxb4GmM1ttM2gSlHnd36L9nbWG15KJ2CVxUq0pkIoV3LDs7XJg
XX52DeZYSinmiVrPPqtdoU/4ScWlE2wz/IXgWz+Kd0ApUNSlixRyYECCb82YUwZbVqg7UIpbZGB0
E246MrClXsYVaJjynTPSrw5BGDeUIUvZhJ5WbY/bHoUoOE1pcyS2LhWUBInd9L4v0Tw9MJbHpHuc
E+mlpUeMvkqfpf/GLr3dZ4Pk92M9vfQ272jzPX5yvNLpnVVxDEC1SEx5pbVo34CWuouNroJqCo0h
0kE/6yNgy0KDaVF0bJlj8cUdEDyt3Q9+w4XIbepEoQ8e3z8MI/j7M9hOQlgwluwUpbGf32mJ7mL3
ioPBju2Y4PE0QMrdo3t67ZamJnvyubYoLVu9eGHR/T6qY5pi6qNMzR30E/Vzeyu9AE+/DyHAr63e
y9WgAPhQp1hYZk97Ol4KgogDtsU2vSbEaEcP6JFVwnunGTQl9BcvQ5QmOko59CTepUczmZIQ36B+
lgDn148zbVWyOMB3cYeWbAT4X1g3QyHl2uPMIZk0wFn8AO/S/QIpQZkDMl1FW5W6FGclMIPp20OG
7vUpK6p4F7sPEl+5ODSDq0OhkOaPWaIbGHTonJyQFxxQS1w/YGp+APDlxshtN3XcQgJP6byhywrh
qEFc3W7iTMir9mG9fIz7WykX74Q1m0h57T4gTcRKiKuRaqkr+36RtYewnMkSpgkfFZPwsBkCExGt
i3ZqTJNFec2E1ft+gIjNsSg82zzRbPYZQc6RYMt1jSJa6U0e0GDw8TTCV+nkqVTLxhyeRQROZeIF
uCiHOZOCxt3GE2n+kURanEYFPNR84W3QcWfNT8NBpbp1E26K5I/LLbncfGuZYjDBJFdmY2zZlksF
5FgGm+C0k14Al7C1oH1AH4+0K2R7zkFrc9tVea0SBDeZe5yi1ahJkwXw8cX3SKMfDUsabBG1OlQv
2S9AMqwRHdug410qSJSzxEllnQhkPlWrBTvWzqEi0FLqNBpx6Zqo5TN7KftXAUe4hLnCw/uGIBUI
h65LGWbld4/wDfqjbMRnGtDH71jjqP3j7vgR296jCeNyRK1dYaIMau8I83aXCF/RIgGuvTHfqFYm
dqgUB9Q+l33nOy6RvIy3ejbKE8l1D6iChT958sxGuxwU09PBI951QpcFXeDqMZCogCACNpxeXq98
zoqnG+QTMgLAJex0e4fv0KTbzqCgTKE3+EdPYo+QgkGexObM2cHVUMbFf/ina6RnloeNp55FRaCM
WVySfZ4A306k3jmq5Mwd/fHHzKzx9CxvarRiPSwJ3/LOkJOlT/UEY2Xoz8k/nuZqFELca9jQZob0
pJRikPwKqG282wHGpic2mIHqqXoCJU7b8uZRzAiTJVUaQTnE7EPm40e7M7FuHAUOWmNhJdIJwrBk
f+3gQDmwLB10110w5eeEIC6vx84pc9DOFc2643hiZom6Hzag3n+DWaykpy7VstkhGKEMXc9YkNOn
zYZNUhA0SyvGwJ4YKiTANpucxqcjt4ZIuCZ+Cj3iHxCRGuaHxZqAwuDfwR5oF8Zz+o+OvF9IuEWq
Nleyy0fVnUG2AHTMHgW5xNYMlMITB89t1aLWsMf85ap/qc63ztOzu6ZT/qK+sXKxItPP715GZbj+
sMsyjW0a3rLbNQRwcLfVHcdRqZ/G888VYW8LgBsxVeHYjXhm1FZfHwOcy/U23+y21+aowe6U2n2J
YqSSDp+2tHrEEIK1Q6guPG7CUzQqMz49RmFIkQuKaeHliYUVWdnTWhnRbVHpqqVDjP5m6NGR0/fD
cLDwH+Sz/MZ1dgl6xECCEe8MxTC6ge1257o7/s9EAQSDaqYFHBhW4MXMzz9tfOevdt7vmabCAkV/
duujCtKgHla9tRRB4jXeaYrL+PuK9aHI3XKCv53Muj619XwGjRb77UY5CXL1zdPNUKV0eOzyCK8N
NYcQTvnYUOt6s5DVcbf/NMwmSk55zXCVffejIu1aYd1y+vHD2OMS6ugy2MSREXI1dhtd98jxPRzS
i512WB+SKvXGM2fWtmVewp9akA3TaN1W5zYrzIlgUKczEV6uORYN8ediWGE3Y1NdfMeVvZl+TVCA
/c9EjpawN9lCCuS040rzk/11/NPvnPMBv84mjMp39cKWCprCc7RygfLhn5i8oP9OIo0uVD5ewlCO
G0KDivoS4MsclCEs6nn0OLE4npE4A0pn2mUwCixnYCju4mlW+oS00N9PPeGFRPcXO2/wYPEw9g+K
t9+H/j9+Obsy5kV82OR7s5Wm+0JaCwJaq7xcR3c0nrE6msMTC7VcyffaVLMZXjNQwNtu2CUtCMlL
0LFXuAPFNpg0zFQMk4pWn3O+A5dlqdma/I7HrXyWeMWZWg4Um8jNsmuHJg3sjV8ATbf2Jpb+wGss
MgBF8ohvf8755r+Mz3j2yO16P3Tqq6tckns8RZz4fBK0N6Cqtd0HmLS3V0M6R9e9ToJC8C6EXK3c
HlyROqeBX6RxbeEZinb/dzJrDtnmgLV3lt4WfXIce2cR4/PyUxkcnH0fAI1Hl9QvfMh5v57CFp7/
HRyVQoBCXmBvf0CKJuoa5nZ8T2+ssMs0BJXWFZDodSvZnadQ5AuD+dBkroRMN3cl0pZgr5QR4NvB
FdWY+vUkFe/hYZofnnqa6X6GTEzjVsitYvYZA1LeS3NPihLE5Dpt+EfwyxlIl1uo5xY/DZjUuZhk
dER0iLc7fIMrkpRIMf8Qeuo7Yb8ZS0OjiAoliqvzyD7ntz3kFnJtnrJCPQBNo97Aum7Vzql8yyf3
c2oabWoJZVT4zH48032B2SC9sNsh+kXTtMf5gIH+WqDKaFwAPzGzcT8K63+UbSHFOt8RILgaEoDY
MrJKRPzfVcfO7fn5ouSWeXfahGcB2eyaonOzDdYDnHAWtH1pELvkGQhSl60tAtV4ZwePn/iGJtL/
Op3ChX+K7gnpevJQNSteIrpYThBAWSCxROfzY4wN9EGE0wimeP/AsYrxeyRdm2jvMi0uXGB43OqL
Zp8d3+BRcWxy+oKFkyuxFxREHBBCuTrZsjp4jHVG8vgav9dLiVK1thouGLXRjTujTi+DS8J87SyL
yWFZwWoVJ4zPb041KBmm7RdoGqD0vVZEYoxEn6slSAiPH1ievQRvxYluOUAEeDpf7o3nXYmT3aF0
O6LJzVYFgMr8IAq093mV6vzJjfwWAsiUqBZ6a6vglK+M4sAEqXDbsPWWbRrnBwwuylkQcGUSOPzb
BET+XTMjlQMQvoOtsuLPOwE7tkRNxBTxOxfrKhwuoNX7GbeDr8HwnGRH75Xns5JlKx8YjIeD9kTk
iZHbKc0EfmR1RwNhVfjZAAarir0EnU6D5r6DH7y11wr69Ts/xDeB600lTYKiAvCKpdBo3xxTYso7
Kns7wkL2Db+MOgAetvD25HQZMZF7YvIFnpI2yvDamoAk1QYZw9zV3Ov40xh9JUG9ThNw+1wJ8/15
M3rPHKmsgobDKUALa6oEsV5X3WwO1mjavwUdA2KCocFhr1HbFJdoofOD3hMpVigxh+VFvoMqVZb+
rphAxP+4EtJETUi1uNaTHeFnDhCM8BjBCrqpvR+mStIyXwB5Vm7lbCBCc+DKQnNla6MUBNcFGUXQ
IlPT+f33Aayr1CPi3BlHK0oxFof/wVnuZEiNoA1m4nr+L1oHk5c3oZBzhXU6+sJjh26NijLFePxW
/eFD8LecKlQuKHTcyO2mjI6WllD7ILqrZfpMSX4L0uPEhBH/GcfUgcocIOq79sLnpvH5JPYoOfpy
lwL6ZmsjqX9Ovu2bN3E/pkO1fjIANXAQI2ARqCV9viCU05KQP8GCyOl7Nih1Xsti0uYSc57HKH8E
O1cks8bloVs598jW6oAiuinqBGkhJovlRwq9FfrGnDt/acqFEdq7o+BeIgJe27b6S8sM6N0cJd3x
yGYzaIaBcbz/K+rHKESRBliUvq9FQvBNCjRAHnJrWbny7NmTVBw7ElVaDPlN5jchoS4KVrL3m6ap
Te+RTAV6DG3tCfJHDAZOo63oRuFj909eRfhHYhx3hJqngilFve9i4rs4/LouL4hvpk2o919uMV0B
6EJuDRwfbn+Y6mDVVpMgVZrrQTy/jU3WFi3Yr9JS4CdgMgE2BhIOVhKNgc2Vr8goGE8hZPGQr6Ei
oA8TAitciuZQ5yvp99ajPUadrEk6KMUsdQ0zfi2GWn5mdYVDXsozpUismbkBIbYZ2XjV8nUgX+oL
h3O0kGJsRYbjvDH/68z+axnqN5LjPbU3ZvI1arHn7PhhkAVKqER4bWSrDfDdgGty+hWZR1AhS8dO
VoY+xtCKbWOjm5b/qq7bpQXHTSeaoGxmqZfrIm5DZGfVPzVprBrJHGNWDrxoFmwZEGpRAhxfBus0
iCBrhcQc2ZWB6y/lI9l1srbLp1iGs1hJDHr1G8f8RczShv9k/PmeZ0vzLrQ8DV9w4FSsDzNKS3yF
tFIQOvPKnIuaUMq+95S08Z96zO1YaWmEPe0vzWjj1ifrNEqezdDcShUEhEjTpAiyk2bVaGJW48jm
SwsIpx8IQlGj2r1YixIwzKTq3XrWPYPAeND7NvXpNSZnKbcnoEvpS34IJrPV1ERaZnY6DYs6TFYe
dwGxPn2sSuWDQQpOTT7QHCKvnPXBvQa3IGGfECQmWyk0sSVgKIf0tA86axrP2m8eYj1xSb/IoX0s
ffMburQQJSzcXViXZawv6GMK+HMtllCm5meH3tu27RKU5/rwza6mPAHA7U1Gi4UflYHVKlxU5kmN
vSc4G8P/kkJJEB4uhzKnD09GcPiAlQ2++bXPBumBAr18VL79ON/DCU6Sm3aYeuOLcy7Eao5MXNhB
zOFOq47V03ZgZAJvGQT+1kCyMuvb/dpXHQfJNw8qHnpd9yT3G89F6YjVK8slsBLgD8HMjYmHzLvJ
EqNp25Vl0LIAx/jd7ntFCLjHP3Zs7gl3Nxr8knMrSvDqPlwuy4iKMp4kd1DiSXB4U5J9iMoiz0z1
uhlKsQ0E8GtfX9177Che7FQw68hPaL6yTQkfqJ03X8WQ2dlkwJfmQ9tTBpv1fETqENhbCILjC4T1
4X6tHv1na3rxoTR6fGz89O+jsEoVnQhBOPq6X4T1cmi0EEKPGW3x/EDu8265+m4uN3TJsPdRwUtE
lAsvGA6kRyhy7RvDpVL4FsYeawo18zpvOLBNaZ0kLvKU3UprnrWaL2uLIzbGpm6wGlfbFOPVe3tz
BASlbdZ2fcCJS9JaWyrrYZxaulE2KfQ+CqWnc4qT6MoAjeRBZ79SgzNZ++VNlqLFUCpNXYWj6I/5
87OXVJd85VnkZAI7iT+/gZlhm5o+f9sTuZMx22lzlfptCgrHh8vgQYsv4P3c0U+mLw7GoGgauu5V
AjtqVOLBW7QAnXAc1BeJ3vlJztPGREgmRLjbwuCamsUuKROoZ8kpcXWHrEjrObSBpELa7YCqJQIX
Jjiof2lTidYB0i3Eq29Ztpg91BbMeZmsUL5PrvYzHQ7d7m6nDjHM0OQkgfPHteYCFRdd3G+4hfF9
bBnCpdtYVP81YhdhDHGT9jtf5zQ+8aflKFYTK6nvV6p0lBq+WhX+of7lpaGrr3nfcKKpVqJVeJiz
756iktvgqidCVRB4PyhEA/6W52tzCphZCp86hXRzDn9COprFcwX3pWWT5tQZA6mWUUFGD0Uw3Eu5
gvekNOaQdmyEHaO1VR3GouxSzpUhZq5DztLn/csL25ldChd3gHSjOU1j6jA3SnZLQ6nIxJOsSCv/
1OqThLjrp9LQXoLMUQhIVuYy8tRVSQlYld4jE2o922a2UaUihkpm8d+ToLfcFMSG8p2012Fui7S3
hfJXo65c81oRsMe0P8J11WsO/eCI2M36mGuHL+CKS0ZB61nhY2MO3EPCGhDgcI6ovEqubI31TgDU
ey91GbsU6KLCTGto4e5AemKTg3lv+aGV/A8dmshj7twEOH/RWJ0N5FGFw7kyE5RjT+cYW3RaMMeI
lZ6AnHVsx359sRriz1cxfoljDVJwUVMCGQe0JvANR9u21Apfq4uBtJhDKu6s4I/tBijqBKPsnlKk
aGmAGsqYG6pAPTdvqsiKJ1tOU3Up6dxnfocHBBmzcWThO2Jw2hymlz7DnOb+x20dWkZKp1vM0rQJ
DLU+hv5iDTiYSzVnpvYGPaVP9psOBm6bBPCwcu4S73osEvdishhZc1r8ZVC93glZ9iJfqngoqT0w
d8nPg4mwIdFOQwXAEdYomXtdjvmAqLWNMrBVvAwuV+ouCqjAhUjP166AbAH/tqaxhJ4TRODLuI03
HiMx7RJVfUBDI+OqlKycLvP4jXG9XOhSSW8DXRowEpk5naQ43TVH2SPNqofZZA2gPsSBWm7O3SDY
6G49PWh2HMEbQE5l/R2wVULx7YeXclz84V55Ac6wOUrUktWWjvMvR0Jxo6pp5Tb7aZeMyA27kzBm
sJj0OnsC9XDRt9jPGBwN7Y77kwJZJOrRKb4K8L1BP+RMjSAD723GYGoe4ABzKBA6R5hHYfQBLwl3
6vFaQMTNRDHYbJi61f2cR7m32NkcYdz03Ylfir4PRADuJNVsbIBL8XmNPD44KIXjjkilcIO9DAY8
a5UZPjXZM3O3wzJQ7CFq35dt73vleKMhQffpWYu/OSxzdGQ7lxW8ChpKXkwdeaeY5Bv1d6Wvtfv8
q9Zn3vQfhUGDeli+DiQYMZNpxyEk//zbWX6xpK8JKUR5RJmGz8K/2TmviPVKIFFvrfHkPcVS696G
n2vkdaX+xAVOBNuuutgr5b1rIXEIY4D1EeUUz0B70eT3OJFgVYA8p2v6ObeFu4mTmdik9pk/XJ3i
sCqWQhM5fy66AtZjTKctjquKWIRJmDdKPHfn2N0hvoeqyWgoscaxULRBBf/tDeQ/j6uxPEH5ih8y
CP++nYeQvEc61UE4g0qSLFG3J2duDLG5g9HiKWR+jpXm0GOKxiddPMfk3vMvQ3eUEGBpxknqwYbC
IZqWOLrV4HT3dHjdANHMi//Hkk2S8U2abA4lFR7XJcgwC+OwHIu05OJ4CTACGnq7WABFNvJrianq
iP1IedVCPLUgSJ6ye3ikA7+kpoGgEujW62Da/hnnJXo5YrfvEJqmJl0MVHiTHBi48T4g/E/6dSw7
DKaQBDqJqh8/1Hyi4nROdx+1qlyW1dWCvZrW6gqFOdfuo3HyDdB9NBP6LU24F3Kz2smSdG14SGNq
kQp0LYbqNpvYlFyglvdEesNlhFECX1o+f5/Pbimy/4fmkW5ddx9DnYgAH1JezuL+hfCKjy9iZQGG
C9H7elsQTAxGlv3qbKThw49vI/ZvN06HW9kgDgnruH9SPdtMECXHy2AHQ2X4vyqsAsAXbMhZMlar
vnruy5+8xx3Zv2JbFs4Zz9tALrIVKyE9/KiaD3L9gCwsNsR41vV/Ciy9HbFggjjPk2Qp2V7K1lfv
6cWE1oeFNjys+iFwSJauRZZnhyoDKXsYw61xOqkh5K3tupJSaFDaGFMgh6ij6EpaVF9xljggJ8Wb
vI6RD1gjRMc2OvE/ITwDYBB4MRt35H+LnYAZp8vFDGgDd4m5pZPv3YVG0OGzwVi2Zt1GYzVO3SL/
2GoFRZD8u9A/qLV4ImZz5g57/QRmPQlM58RZc3S0QUo5jFTUu5VsTIdE95/8R6wqVf/WgQ2CEZhC
TbuF7qcloDt13MQbAsddXX5qjxqpxthHHsGqHXJBjJuwvKuY6IVAIxJxJ1yn4VJS2iovbfBRn+0U
3PPbuA9FUCVgHUThruBFEegIleaxLJNq5wfH4kIsbgk1vZzVIFVqtae0t6UWYkQuw6o37oeTCGgi
mjgwqqyAFKcAJhVZ4+a/JlxJ1LSo9T+WXOZXt0Liq4zT7InV2y3ATlZYoj3+MO4K3hCCEIzyhHnt
bLYhRR6BvelAS5nZx9+cT1ZZ+l5DG4Q8M9bJRbG21y4HNtfhgTBOQbHSqTaFvGa/cnosrXW7oM1C
lA6jrU2orM7R7o2/C9bhicGH0Y3YBuV8LnqbLshKoaIF1Q/Z0h9ANYEKSSDrCSFuU5JDcgYoGpx/
7V8hGQP6bIWhzW9zjvIqGuAWU1EVKumXqMA3Xh1slieWqh/vzn08Pa/+7vG8dVOFt1rnqtMvF6lG
k+RAJfwgkpNU0v9RrPWci32CrRLl2lXJHWTdvFZaowimGhYUyIDdktFxLi+sqVBxjEdO1mHDjzfB
KVMs3ZwebWIlhBvYA4eFRI37ebk3TAwZ5i4Tl2rjGYsOmcrQUDS/kflM5HcgmP24SkYwR6rIqFFO
zplqWGYQysjpngoP5MfgTaFu2dBDCW/Qp8pNtiMQtXfwhWYonQK2YgXGBqNt+64fKeeipbOq5cQY
vJ4GPMNNh54DDlKfjk4s7Mw/9dXkIoCNasF6dCqEUUm42R8pnaR9/G7VG1p2tcj9jR8Fkhft2trZ
91KeKRtAF/ftMAK6eR85B++poxNudgihehzq7UCJLigppZyb9CHULLGDcWQJrFF/Rzjee+v/CZkF
ECcWszdNcn5A3uXFMZ50W4Fv8QhlRRJPXJL3i3Xd6MNlPUee+o45Y4wrIRKa6/g2XcH4g0ZnCHgx
NIpX+hETiqTFVQCmvAArj7fT74+DhTJSX6DgfY/A00DV84wubHOwSL7Fl5AFwo+5HskbnHpLSlGq
8r4SaLONqRZQQt8KF8zg4z/RNX0iW3y6zNqnlYRtW4mdX2rs16+laokygpVro1Rd40oWi8DHe5OC
O/68YaqKCZULcBN+vDL8QAQSFsP/wMzQemvvZz+5euK1Zm0+WYKbMKNSgvQCXHP+bUlna8kyXuy4
3cuMK41c3HKtmR36rND+oR18oobQ66O6Nay7i1zH/twgysABXKx6lg/3DCPWr08tMHQ/qVF9nhHz
KwlsPtjarmKIaUhIzncyAoOrw1N9O3y+FCD6YsU9z4LBAUUjrGmpRCFkC6Qa6rgF7MKWl9ma74UW
IRGlLu9LHLsOXG5pLhwE5iOr9mteH3XKmP++5s6QhBlPw1a9xI06/82ZfoJ14M5O34WCIyAD/eu7
CFVwiSM4tw089SfMEGxf/q7+4J9PTZASIYkln0a6mIaRdNV5wZguheYoFtX81uHgOs7GGQJ2EHm5
+dIQidMAPKaqpCL929ztnYE1l38Jsx/KTTGAQr2BIv2j1zfy+IEmfMGOIsiJvugTCmE4xW7nz5Fr
B8DKTzmdpVlbBp21yMFjPfD7qit0LUCBTXgKs7Z7D/lLz4YlkoNzmko5k3zuieh8of2jBfxMmKba
j5mDBKaPAqEJNarrmKeSZzlIU3xs0M9ZjVxC0MRkyi/0OFbxMuxjmn7x1f+RKEj/zk/YNuDJ1/1H
9OJEfMo4dYMaVLgVtyUJMI93hFyUQ4SgOLJk1vVtzbTcepfL1we2Zoy8sdt+6PukmVtA7AWiD6aL
Lc+QNwxHi/MnfY3ocJ6iFwwYWomP+DNTWSVo41QzHb2bYHTr87GNzuQ6F583r/HkL6MDcyJ/ouRU
Gl8QWjg8FXa/vLCA9pxY4crUeA4Hf5UANkLhsAk6hh2aw1yAgRrVkfku+CkSIg9SafU+lD7KLY2a
Nf4V6TActGBAK9NamloDqw+P9IyQsz9DT5J4oQK8La4CbYxJpgWx0MpZMscNDmPl+e9fjSmRoCIs
sbLuki7Kb9i6H6dDNxH4G10yN7OnZ1eIQUDGvgvzqXQYt2AW22gd9tlBlA/yPFgxI5diLBdmsRL7
V1NfHJtNnscO1R+3RF0XEWYe4ZaF59hhr56xzQoqLYbAr7N+VpG3FtpEGf/koFJ5Wd2EjfuR4Zik
Q/mHvEDlbkAUJ5GNmw8NPVUnep/MUa1UffvIjHkGbmB2d2S3I0UUsoQemoWy/FwUHtksP+3aPfCp
XX57TCiKLaCZaWD1pljsZWY2xDWY0uN46awesVh8mez8N5pGjLi7Sr4rlXoOpJeRbkQI5IJPOY4U
SJde+tuFhQkOZ+3XkumwlRZbDtYZ8syvYB3zwGdzL8tmQAH6C0sorvfDVoK2knPSAL75bjEj9A58
Y1jW+a4fRVoRb76jXtk44Y7Z0DdJYFIVoUOBFS6/zw2x3wNG5y9eYahuI8sR/ww3c3T9uOr4o/mG
g4zGP/hrYGVY2WXdw8vvERsFbfG/hQVcBDzTA5HDNQBIUQkZaDHJqKmG2oSyb9rULMk3J9/SkWMA
oVXQAlJlGvAddjRx0prgaMvOqiywbcBKcKm9KNJrC3l/U/c6cBZYB1aYsDjAr1WDtTbA/HikwPWv
r4FM1g2ol2ufT86751TKj8O2wfEcVOFH/o+N8pGGvfCIGt3kynsCGA3InpDPgvapk/l3I8e6g6al
spdCL+lyNZ648flEqMp4x1VNJcYqSYqJK+Suy/aFvXmllZm8XE/Us94SlpTGn1Da2Gdwb2QHRZN5
9qvG0AeHTbOwooKnoYsFe3nRRR1LEtidnYYnCxXhjv5UWZ3gOocrl+S3n2+EUBznlyGFGt4FMMzI
RoCqc4uis5gnpt+6wceobuMfymckWIHhHv3m48bIQK/WhEzizcsYHxSEvqOoG9LcO1Tg7BBolpu4
+juV0s4nYcRwC5daHjmz47okdSai4Zjczo9X4ZHEXU9ogZgkZqX82ioGdLoQ/eVJEFwYZs1uKkMs
m1MyvDVNtDyfsKhDG0n1ze811SuD7M8ReAbUrKzAQ85zQeLkcb6DalvUzNA7iRPMAKp4OcN5IIJE
oTN/GeoS+VSgqglO3guuOi4s0KtbefUnywGyVizZlMEaZkI6PjXAilMAWrHoU0tDGpXHehAlSOik
2hQBJVcrVspgdpwZbXGOZef6+LCNAX+0sBEu5eVoiTFFfVEJswC4D9sVeYbWWJlJMrtcXaT3VyPC
opJPQNvTP1PL9uvW65cMXD7jdhd/es0M2CgKKwEjmG8VesxvKCpMXei9QPvj8mMbR3H79tTjvXL9
QEZ/tVJ8ILFLrITr0J7Kr49y7E2L31ILMSIU/Rhu/fK5Y7iGrB9Xi6mfL8dZhHV8LOrDTg9t4kQ8
1JPh8nK737QY5kiAId/rAS+WEaZgWA4/2cDDbDBE9gH5G+eFgEXKCoZvtz5vkTDnsV6EonzsGDHu
K1fS+JY7YdMhDmwk2OIEF1P8Pgvmw9I2dMjwUAErkPc98So5eD58IiMSuLQTAPXamHB6/Bjuef4f
gb1NDuniX7z6boRbx1fQutjN8N34WI3PZvO3a1xzpS8kB63MHif6BQ5tzNrkzBbpmJ8XRI/rnvJC
Tr9sT/8RHkHVgsta3gF9YKd30XdLApxc05O+McisvAnRgumyUWFfq2cheTuFc6/6sR5Srw+/dd5b
fcuLZ5kO3WIzE6jlzSr6oHp7hgofVG2ObjDd6MpWpWjiD4C1BfLnwMaK87iQ3aR5vhIZxOfHxQpJ
EfLNAwRD+sW5jRU35HxfB3R77G/qZx0q84x7YFfRaJQearP1prpSqkF6jxBIKQv9BGeeO45R8wLa
x4OkaQpJVCrUp2oI5+/qI49/hAYsW5ZvcA3fy82RIydg9nYNtQZQPmYy2psVQngvfmNzucYoJPb+
NLAhJIK7ljQIi5pIxp0W5QWJJuE9kVpVdwDME/mbAnOiiARZgo18rtNvWVBxLPT5FnTgii5e2JA5
rwpakeTmW/olcZM/ZPpmqbchj45EBwB6+fXucqP4IFG1gOMpK6CmaeoetE5WrjJd0R1//GeRJChf
7oMfZSECd5DXl/aE3E0QC2yqGWV6au2CgagK+KdwnD4Hky8nhmt4v30aALmjV9qoh0ji0m9Zt12G
0lCROUpqoRgI8V3YHOTy1e3E8mcpqNQ2OPSZYyKLKtEWAHJ8EvAucUPm6xKq5rXJhWk8ph3qc0TE
Ya7Y8rp2aCfl3OJGZBddUM2xKpxIXS37vAbsknnApS5ezQM+Vx40rv3/mA6nhlddWfMKsCwzyRS0
SLtknvGm6hbrRqqL2p0wtXCZbQAcP5AVUQKbC+iVXQX4wgHMKM1bTYRBN5BJ9DN20oLh/VcKRYew
kqE4QmWDgXPp59LDE6VgdUZxpkc64KqPzpCnn82pXMjmKQ7j0Ij7va64pnwjdMz2doClC7MdVkau
9UdXTshW9xufs00NzVYHQsl72/IeIsfP8vf+087CqQHNO9mx/TzFCw0NtZ0hcQFXFRpP9BZJooRD
2F6IdYnrn3iygMxFVpT/kz33tmWtgoObF2Oin/gAH8m5cynnDCnXn46d8ig6b2k6Ts8sDwAQ1cK7
P+yTgsJ2UwND8RLyPdHf89mIBFfnT3Sg1WP/PFt+XJzMpWeZpoZzeORXrMuWLNjFfK16B+TPRllj
xBtZXGFHQsJ2DYhQNQFJaLuoBcN0dyggQKEvRl9wod0Mq1bri+gYzOSo1o4ywuzGz8PNqMmcphyJ
q3Jn39YRtmKRzGlfxzCw8TBN7FpbL1GyZoAbKKt5a2cO6ftDIDWB5haopf88sjdJyHdpmI6F+Wjz
+vFnzb3M9nUPnykmkp9USULFi1GYw2IcFGB1NJk2XPFB1ju/uIBfuwc07XzrxlBErTmgxevikKEE
0TQyY5VyM2zuRvK1ExSD9NphgbEaNpywcJzRMAkfl34QnGkoJFj2ORHW/mDaLr1kHposOTMFv6Or
4w+39tK4r+vFsr+/g0kt629n02QRfHXGWAzunwY++agbDQFw0+s22+5OrwRjvtnwu5yORTgSO4i4
2koOp/+9+KEUWXZM4fQ+KJZU1pF2g829nZvT4l0YwmtlGaUVSjfSOu33pI9AbidUibyV2AXkSHGn
DnWT9m27sJGx1qIhU75onH5FfSKtrrZPtQmoq4TMUqlM+4csmoKaa1X+qQqX7HARqqkasGfc7Sdz
+EPxRmMBjdxdAxcaodFWcAhuNKNXiCkXytByXIUOSBUGV+5wABt0lez3SSpwmMyIOqQre7/4wJV/
VmmJ46Yu7KO+7GdS+6D7BycQHlz1Qp8hlo7dRCiAA2AXUOZ6OGS5OerGk8WNt5A5Tl/it2gRD0ap
CMgce2CGfhGxPo+AAI8+zFhHkkO4xOtIqnoeODvbYEkQ4sILh/jPXstB1Ua3PUxtgDRtKzVIxJat
iMTtpou/i27zHb3pRunhHHi30NDJEM1xbVTw80aNtUSd7Vf8NLn/DN2R20nPXCIauyNmbOMwiBow
Q5THpfW/nP2reObRBHc5aAudPeuiRuFnEfiFDQqkP8BsT31KxBirOR/bfwS0X4v4zcNR3pboDxvF
NPkiheG20k/adkcAcPSbzHiqm/gLGURarRuKm+Kbv2kSoxWuYtNwrJDtp6c0km9Bi953n+mln2hP
6jktWvB6VCOFmnUGZ2xdpE5ng55z96+jhiogemFnhnN2G87hQmyr5B+tkmm+euLpJ0QmugJuwHPd
HMKn9WYfryL0QMqajcaxC0IEiU6LORIXjTTYixKdGNC+HbafIVNYOlirqgsu7cfTjHYO4xtfEIWm
MZxfuKfORM1vSkYE7EiF2yMJyvKfcLY4EaQXuMKl7EU+KS+by1uRc6CfsPfsBfmI5ybQ8OaLg26u
UNzF5Z1I03mCoa4stqzBt/wihM6R/BYaeO9JtyCAAHgXWnUxi/4R6v3UMX+gnkhgJBygZGvULC+o
1g++H29KrphKdYt4cvSHHqf3Pms/ENTEr+4/OqM6+lpJ3gknIABlxDrY9Sjlc6vZv7SZgO1/3KRQ
sLT+NjaSEswUM7x7uQrdbAXypy/48HQrpSOW3HzJJy6bSE0N9JTzy82mv8YG1lGle9aCsAf1jVlc
j9/FS/1pYhp9GXnZTk9yqxp2+IncWWNooYQ6IVElRBrd+pcbMzttg4SyNbJz57nFUDW7kkaqDfdy
cE3sD62l38mftDMFYT6yycym/Z1uUQSBpoRAQ4gotEFsMw+UA6cQFS2p5C9SUHk0eMFendcRrvAI
7qyOQjxrGpXE16u22+pMnAnIGPpcU8OnY30ZoBfPYTV0EKeGGmujXrlFo9BDur4DOc5c2J0B3EBi
xK36pYeejD9oSncLfxSCLxSNkZ+kaJ1QYXm3vmgxJ5gsBZ9Za8STPcLhvw37aCnYc4hw0VCUoHwI
oF71FTG+CzgqL45YuE3fZPaPY7pj0oOLKtzLnQUqCnS333JUY7yu8twA3GZENh04uzAe8HQAx9Jd
wb4KUP2WJpsyFf9Edm4eSyfd/0PWEEBGk+z/AvmYVCvTLglWHphMoByJInJZOUyEMsbKHfb6G8QJ
9vtBqSjkV7qBVXRWLpO47lx7fES97xf2QwJIP0/ibq+mTxl/G/bD+YCagKWiB3BdjSRVKGPWewn/
Al/3ZqDS9RpEMC2MRu6yhYhVteAEP3Vpi0PUXhoCab+Cte862jPg00gtpMVprKz9zKMRqyunOCec
Kc2HLCdpwqmKfMif+bBPDGJvfCyI7k1At9U5OgWyKvhNjjiLAzSLKWjaNBqSJVDuIemiSqol2w3T
yRs60iIe03vYjNYhHo6OHejU+HdC2oJc52Ryqicam1RWKGT/Do5Wq9etx2rlDiQPwy/KNwnE8HFX
jnJaTmb8fHzCR/dk0IbE6tSKtCkppkhsZJKSdKKX9bQZSD3AMrr8OX885ie++whqZ4ITFWdzc30B
ml3iPXmhD4IAgQsYAZ1Kals8hRHwBF3YElZdO9UETGe0138OJJEf+7IzPzOa3Dt4dgEqBWmNAfK2
GKaS8CNyvWTOzAYxKMzuSkknEgW2QG+V6vImD8gww3E13cEW+9olAz2TMz2K8RPRWMnVEbttVlKM
LMA35yrn8fWVmMRrlKeY37UCaJgDqo4URr3i9KVhNIsOE9juiQrllefZVUklQdtTfB/lH8oTOqLv
4WhnTtVOf8fAwHrkUxfjCNjbmakphR1XT1v9+YxvBC5ewCmykc0gUGw0R8zlUjioBYYyZqm7bg3E
j1cHk1tYLoMs9q0cSMDxSMMNowcol0H86PBx4XEki2jmfxMzvFF96uf4HaZYuyUNkC8ekU3it5Gq
k0oqED+9hAdrd9exKc+8DERkZyAoc52nnHE9vecDbFeynIXAf52Jdh9Q3Z1rTYYASxc6jdyb+Meo
DEj0TiKkvYUQ1ULc9F3CE8thSbhEj5f/FmldyGdT2xBuB8+Ml1lMZSTLJt7nG5BBYnX4mNsi05Kz
iqTV4gqERG+0khNSTZ92wz+ZggmrhkHpIby2Po6tq+744Z9w7zD88D3F64CeR1pQfqLNkdwdU4Bn
sa9row4npm7CuLkiAc9qrJAeRnSSP8OXFillWVTeuwpyyEQGqa+BkE8suQ0yk5urI+BQ5bfcnAgj
Yg3W5Xdhg0A/tSc18QvHmRHpcsibpd/lzoK/RIDD+sWiIo+qKNzcdKOzokWrkuEwcy3PRNX8b4+2
aGj3JINWTV2tY+Ca372vSoH6FmjoDN5Z3AcotJAdcFlqurYGbk40V19pUKhYJvh5iKSFkeV/u+Ws
PW/aUqAbu9uglA9CwSY3tVPfydXSi0rllCooCWI1+5jwZB2L7Pko6U/eb5G0BMPwjRYWbUUqrZOS
TTbiSWfo7oYTcUK/xY9UqzIINX5ITRbLOrEGOcxtqIZPP0FdlRXwGD//cZLU2WUTtgMRPz8TCaWi
aW6vyaa1irlyFd93sImw6u0AJ5PD8/ZASrfbIxd5c+6433D/2DZAUT7u/bKW4WNapFETKOgIohTt
tpbyTzAYTlFMBmYZWFU4NBjQ+NzvIw1a1XsUq0kQ1+/vyAy7So8w8m49B/zF2Vcv47H0cRRv1n9Q
zOs7FG2m7sGTCev1nhJNkI4B2qSm1CtZOisp35iFWIRo270JHOC9286k78CO1lVTgoi3e0ofmpid
xWDinavM6ouyThxK2ONI7GFtxrKbs/uHMGkBNnrQpA2FaI9uo0R8Q4jx8+jHBlZO54dlA85qfEog
Zg+3b6HBy1hofixrZ1+p3PFVxsKh/3kG9JjWwy6UN1yzLg5T/YbSk11No2ZD1rwbK0wQJNzdnplu
frAU0QQExDjBRdEr/TXpvCo/mZSpRkhpiGiOod9Y0UHiXz5orE9JrCLvwG+pmYqpCsHFae9e2BaW
PXmcMIEaZMPvjcPPaJgPF1GS6pzV1ixxMwtr87zTRbgPPVsHe3F9C3jDkXg17tZNynwjNBUO55ne
+9APqT/JA6dMbJvSK0VhD94cn63EXznOVRx94qAQAkevKAVTRrktQN1NhBGNd/6UtTiZykmABnU+
XH/VRSoHLfskei8jYMQfGQTtKxP5S/Png1rQToG6BYqN74UgulmQO4szMAw0wy8V1OtxsmuUiciL
tMgJCxt2a/IpUbT9l1JF5Dt2VWAJkz04F1a9RJduDFlF6cs2KLzd3AK7l2d4CT3oro8P66OZRz7Y
RGllHQ+AfINBGZiA+kOwWtymp0ZIcG12an8azTRJiLWCcsO03yaRtYcDgHsjzAxdKTR5mhAaOcA4
pXyPsmZYkQwQjq9R4PpokBJaBumBiR5F3xZbOQUuADLi+2OwwbpTJoxJlHPI+J0cNxTDXhJxfknx
tq02tM9QH7NzSy7vKSOZnkzGMNXD6b1O58rcwv006Zw1IyG35GqgFfX3VIy3L2NZ0byjTobCP+t8
NU2aMzKRLaT2wEOdIcV6b4uZluX7ecnv7iVa5XZk2LAczcysw4K/NwwrPtKaPKKqTkWDKdr0CLo8
64fteZPQSj3w+9JoaP1/uN6X773ro1KMRa/k53Dfe5Q27ZkxrU2WqVnpyG05B9TfEQsVKWUbv0IU
/PH9dx0/r0qsU3wa2WXvAb6OzA2Pn8VCX6hiB/1mffe9ui/FPmJwo0HqEtro0mrbxEH+6IDbTLKF
jbDgLulv7Xeuiy8HVeuByS9AQGI6Y8FSCL7hQc7rtyGZoRzM8W0WPF0xXnsHZgKs778f5kwFydv9
bNeAmn6VIKlrH4jMj9Y3yOQh2Wq3Lr/2ZGjnACLa/V+d+GC45DQppOmIFNv9mWpIvG/2KUAhNj0S
1r6j5sErm+QC3GYIKZBlfnkTwocjp3U0zldEnwsG/9dJgOn4ngJRQ4UZptTArctwPRj0qYubqvOD
YZmKuauxBy5A9HoF400/1P8TeK1GgKPAkD2q023ZRBcFByqLxgpIj9Ox56G5T5z043lJPlzNYBfl
9jdYlcme2bu9FT2U7KC9xTPvB5oS+yuw+cBHJ0YFgANzOfWUpwl6sHZ7nghkPdEUmBAjwDeEYEGq
mZUFKUi+YxBwYQaKj6N4eT3AENkFyXaK2GGKmWwIn59tZEgQP8ikcrDNe3fiVQIkkOQOcPRS2EXd
ZbNXcnJc1EHHxTQMRov963QwGgccwzoFw7Iw5vY5nezJ5pJycDuhyQhx6lo6ukFwPIZikdmusoYC
HVOaewBcNkft3SLhrmiUCWMIIvttqx0gAE70l2ZieghZzrro5gYJxeUwrFx2K6bd7Q/w/b72G2RU
Y8XP3HVPz8fjHlDFO5yNsOxwUJ8cN97R1OkDcsnfjUuXwyuF5eXjdXDpcY2shcokPYxyzSlW+92C
04Dw5iz2ZGrY3CqhgIw+eTaDjQyEywdjS+NPiTnB6/dZFCiCu3ikr0HM+ZvIFRfg3jOSsl38gEXW
BFcYDa9mlCm6fWmXDzzKYgDtb1zOTjLvVWv1jFnyzSDegWY1cFr246E57la+t6I7+lFuuZS0jyX0
5NLvuxxTWJ7y68EBAWQvxcheGuK0qVCVAZbrd5ili+EWEYA5nlbN3wA8qJb3tt2GvC9Bj16he8Cb
TUDa+LwhGit3thBe/sEF27UHon4flDcHWxSRrLuk/w4p54nIX+fevWNwl5SmDQpblCO4bXvMM/tw
teHCn/ybYPIS3elb06R85Coi7EcO679fiE4acmWc6M95v6mnW2hL6Kc36dkk2EQeN9mncfoMOk2d
iffhayRbLl4ijb1anHvYGYe9b8NRI8Mb22ezjxTRsBXE8LYzXul7kYyfs5hKWzdYQb5Pt45HjQS3
KntulK/1OsfXSwaC9R8NwE1l6QDInHvtNyTJpI28j8DcYa72+ymfbrtIJ3C90pehLnATeJpOUNHQ
yMEd6jpkMbLebTzUkkh5W93sBvHFDVBhYHl+jX/XIZvGpOeRDvmigQ01ORsVXlxUq1MmwhKFrKCE
CDY5x7Clcm8U3QH080jXA7oxQb1zmCUxMO9e4sEZb50ptrls1LPpLVtqo9Keb9+JcqNkWVi8ZS7j
Utw98k1bjOvQQxMF+Wdzei3yVou3LSoIVeU0ZUvvMjFKNPBOkU8gqryGszdL5kBd1tOmI3gqw6rU
hm4NT//V3YBBFlT4syDJ3/sJ90AgCFxPZ87Ut/rnxpzb9a7JdMqQkEqs5uFLRNzi63q4FSzKmT1A
Ic3vTO/Cw19gNxRoUUKY5dPOuE/zYkDYKJ5Kupze4oqJ+1DhMG/sgpLVAtBO7JMZK+c7Zj/CVcpT
u68+mbOJDl5WYUKfjB9y2w9W8df/8oDZLzAcfiMh9mk3EFh8hNYKkXR7oIRuX2sYkatUKbf1w9d4
anICIGlHQbgO0UpeBDR1MuXditLvzVpoQTTXAzPO7ceAY1dOiC/TsXlaCzYo0Y2fNy9sqZIjp6pA
KzFj0f8XurpXPXsDIbty/Rn8JUyxRuslwk6GHmuz52jqbIoNEY9zWB/5ai4v7rjKL35+b4MZYkpJ
/QMwBsLKUP6Xwph0mxWteRC7HPa+613gGfpswicbBA0DCAYBaSfuKmUQSRtfxVriNYuwzhxdGyqn
J8W9naUxr8glR25JwhxkeR4zUt6mxDeNwqWhNDF9ls1BsykxbXBRJiLqgfimvr2da51PwJJ7gXAQ
Otmlnxe8oCSSKbLbk3DfrUegIzRjR+mukFxDfBpq51dWVWZwYYJLBu2xMUJPXQP8qOJsN+wQfUu6
/x5Wk7kcMIeWJ+pPuFP1NMdOqNKc37B1lwaNFUUGpZoe/LtzIb8uKIM+Q1nVo/7Vl2upSfPXUhz2
veizHRByTO5zgTrhsIXYYWIAtG5hIBk5+qIZejt8J6OpbDsy/XiXM5EG0/H8KOa25ItxQRuiNRU8
aNreC63JEStOJg15A1Sgq1KjHpLSb002UgPfxAbdbdVrGzPiBe5zKzIR9RBJYE/Ea72vvQ/tLEcJ
4dJ8m2ugD0fz7QPl30MHTDJW7viX0rBk5k1POQN+SOSiLHhyLFj3OrXY68/X0GXDjHt5nssrCUiF
rH1SQy48T7DcLCLbCi9OGvMpyIQ0VtQ+g9Z+x06CYxw9jcvxgO1qX81LSXhtf7InwV4PqF/q9uvK
acSara2eekwkhtYo59ZMH4SGk+KFlLxsBr5oCS8wCvT2I9f/G0KCSO6W5oZz0Ax/Y4HkIAKVAjG+
wxOyI1x293uYmxzT8iSCcE/NZ55qBtCQ6TfEB0Og7ZAsv1Hebyd9Kt+coHFNxmBg+Rw05kTSIFd6
Wmoao7YspvSUHW7m5A7nAMgAm/Z17Rd0yx+WLiRSDb9lYa/Bq0GiuJQiqbnl0tdzm+L+ccjk/m9y
FNO8vLUTDhbc74pXVaAcyiroSATIbdqc9Mqwnmnva/ZO9GlvNXZPqXGbQflP6TH+9HbXbBnfl/hg
jrcutRkewH9JmQHG5Totez13+Ol24PMMhHkdNOUnGkHWdq7c+381S4KDaxzc5f0knYIXHqcKwwc8
pDaPaUdiESjOCZESUlwAFGaf5eQgsthNu5oJghfev/R0/DUNsJasSViFT+OK2QbT3zuFN1/F1TtJ
HcxCIZyZwwQ0KiHZ/SPMpsdMKfNcINRncnScuNLJkD38jI5SsjzdU+UFep6JLkViR+6yr4r+gXEC
Hz1KAxv9NIIJ4w/DVAH3c8M7DubvxISXfdKnENt7fiU9JM2iGW8OSeCdT/xKwztVLnVLM4hQZ1xD
SZZ+bT9YNlKIh3m4EPLVbvCwplRn8B1cqL3THau3dDFJXotztKAKV9xGs63Ig4Fw3YnGBWjTJTAb
bZq5lfIaYU0DgzHreKpp/W471p8IQxqyQo92QNhOhEB4InnsKItvblSf00AfaRJnCT0WjUolelJ1
ssglKDlPVto8nCrnaQwGPtZtGvzMpVUTyUT3wUUUaQRNkoh3W8rp4md6Sp+UZKziZHyPLLDakF4d
fCA1c8+SgRMAYlgLZcR0m35oWPyjSVBlnTVnmP4nWQOY+kl6b+IJcndlHkJM3O7yeg9ikPs5btN0
P441c/qTdl2buQzjuXG7rnZsy9YpK4MBpqllyLHAz+Mm7v28za2IgyHJBN7fc7+4jOurydALND7W
z2pTI+1/s8bhGu6TnbvMuI7Jq+ANw1gVjXLB5d1XnsnO+FOJnNMbpfW+zREQwIHTq1+IVABY/bBS
inVCJk+CcHWbuBL+qWxxoL+KHPHalNHYfS0ekGATZ2HdiljEWadh1xRT+jepDFnxzK9G1HA3stpK
WzWslstZQLf1rOMUke7SsbKNlyDxp6+z6E9e+Nv8uzG4BDnVrx+p9UsVl324EDKU12Rr45H3K3Mn
xens0OWDMQXTkseG3CfbfxmF6ObEb/lAUAWUkc7PUWqkRhMQnx82diDNSgvYIbH8jrn3cTP71OnO
oma5XsSN6eMQHQatrxUSIf7CJNrl2P1yAizg+aaYqWVaIupjDiEMA5vabbtfKPkj4CThTF/5wXq9
BaOO4mznvKoyZm8ArE83AjN3uIkE28SjzLtVi7DYtmCpkNPuXyfqQuMXEnVQBQKvxKy/DkbhwRbA
xCU74sHGDFJHnqZBz5T4cULLNOZcmZC2Dn2ykMh3/owdakIrQTKjBmE+UBXgsIfEIO1rLNp9zKbl
BzCaDX8Gpmwxz4lih1SWJw0ZM9vevyyYD8xrj0h9Nbi5+laTbuKsca9NPV38P3QYfv905D6tHHvJ
ig6bOPn6vxoC/24A8opuz93XFofF2baeKb1+yBHhG+s0S9rQmufiW7AXFL9NjP5/TI6QdsnPUfRj
lo2c4rxd0ELNkGfuUq6yDwob5JZNUtRn9rltXTJmBoiuE0ToPvbxpLHumAJDoAL+qTvGArL+T2s8
C3azxYLcn6PeRCCM2hIRz5w/9tr3a+WQtukLmXmcoqYEfnqsM9iCTBbd9V/h1VQ6KLTEd93hsK9Y
HIOJ/Z1+FEqtbRYimg+yy5uQKdyLHE+1dpAv7Z/UgfYqGyvYAOmGzYldrAlhv4jxVDACHjnKlRem
ZVODLTV831eOxtZJxSHg2vJpgawK8HL3dejtnDCddZGAl3XBazHz2chKWfLwov02J7Jc5YiGh176
QqeGIAPGB0qdt2k6cLPW/WLRZ+vIGY6CW/ifLvOSvpLkj85tOBr/DIGbdd/kVn/d0t8D50mztvOs
OfZnVxAaIf+mi1PnC7NnEGOWfYKkzpIR9pciGMksQn1s1QfVzbtwEWnVPRTH8deD5IKZ1/BHSXiH
eYeNmWscxxq5X9rYH5zCemMPcJ2YMPF9LiS3GM+dx4nJP1MFFXJhyxK3t/UFfF186G8sZaIhhKRF
JG1N7seB8VoI2Pl+l8fcC9TOROnJmGtP8Bcks+ROh86nFY43STPqPGu7p9X7pPhDWp8dreYrgSRC
Y4io7CoOL3yor/zfHC71ukKVeQMKh3NR20hlPsVsrYiqA80AB3Jtcr51tZj59lPPBQk/Zl+n64GN
Re0/352t3kkEPP1LoblLX0Cv6JTk6SLrd8T+e8SjN1PQvWRnhQ28Yly2HBH5r7S9/PlzjuVS6TPl
flomlrO3cD45vnYhEAUhchp1otHmAbmzlvfl35/Sj7Kyjb3iTG6/ssjzPQVXnLzjOXVxBKutjMkM
fDU3ran6tlbE8zttZs5SUi2+2+zkNy2DQl65kMAs0h1WnGgmTKg6UpmoBykepKq7vkQ0Mis5Ty/U
7FC4/ufwBv7GCJvp1S6rOZP53hwrxGCbxgXSsBbUaxiT7dGsX4CCVwArg0P2AjmO+UHBCp66nAvQ
el0Akfn9oxl0D8bHEMKdsSVckQMtYyOSB5VIEPYf//NjCUh57NBY3Kc7dlgj/aIdV6xBvGu9U7D4
rkbOAi6AD6hfaTCItPSmaG1F/cf1hn5V1ej5FZmRlplzgsNMVK9fS1D3iAqIM+TUKHVu73Cxr6qv
itibSlwLKtTvdksKxkglJ/zOeROyggHvHmuIvQ9b9gZUIAAdde8ezAAJPcqTnxddJTpJGXNZNmQY
HY69EKiQNi6VlOtW8KAHSH+TY0cqBLtdL8LnLJprXVP0yJ2kq2YmZST2vN9LtraYGuT5W4wz/P4n
juswtmFQ69ChX39ek2fhy/HqN7NRUfypKLZzSsf9aXqbB1vGH5tax70vRCREZ7zRySFXBrDrXzIW
Z0gc+qX9i0kttsrd9JawxnbLDDAEtKVtD6T8D/T0CbvxtA/XvCSY34Xh57jglV8ppNAKWxTh/ltw
Upujrk7QSUtyIh0fVQU8jR/5f+xq/m6jD8oVrCEHwgr+1OGqzrOIaNxiBbPn1UU9ELPStENl9NUc
kLe0RN7Zrw868hFVdiUwKL9+uCQ6i/xrV6JoThVlFUAJMldb63JYMdfLE/nzuJ9N8RCT+90=
`pragma protect end_protected
