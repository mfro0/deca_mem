// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
q1wN5umv1d9d2g3LoeZ9CCg9i5us+Hkzg8QnBhBfaRLJ1bE0jplsNdVJywKZIIUH
Vp1Nk15v+17l0DnEuJeGQ+pvfAWHi19S3FCIbTRhJujYkbv2GqnRyC4j+72Ikw8e
/340dmZsMohqtKD1agJ2/HQc7u4TeNjVUjI8UfmIg4UmfbsUO5HFnA==
//pragma protect end_key_block
//pragma protect digest_block
PEvJV/qjus91n59a/4+dVovITYk=
//pragma protect end_digest_block
//pragma protect data_block
PPb4aNBXjTuF1qwiSgKtugpg3ilKR5NKpdPGh5gqJ41x9E78UNAyDUpeMMAsf7Fv
6kRlMGncrxHzGaBcTJOOHZ3jVjigrzaozH/6j6uR8xxPcox0dQhkM8nKZm1lEOwX
GpVzMZsxXklrwpQ60KbgXQhb18f/4HCu17zgJjDDfS1vhkbE88PQGnHXoMw/6Avi
UH79gjCd0xgOL6K0zSjuPZxo+WFu2mUX3330Fm6FxpjaoYM4adaVFiJJM7RlUE3a
WSY0iU7HpA+ZT2fxXnxirJlBKAAI2eBJsGoRx6SOpzvJKAVR9Bik5eTd7kAC4XhW
SCyrwXxUEI489qOd8dDORU5tZuHN+B8o6BB6zRlB05UlUjEv1DO3CvsJ1hCTlNg6
hhF8/aV4I60bQUDE6s6PFrTeZIOBJGgQxWR+1O1Mkc6nDbmpq7A4SZ1yoKxdPC8/
0pyztxud+8E+l5qLpToE/a3qqQj0fkWkUP6OO+oUwIKUXTK0SDYx+52UtXoCLTtP
stVFYpcEFOiSAS+4xSpDWzzEWeGEVZPUOaZMaAS2GHPs2jIKcx8oz3K9Fb9aXqX2
fT3GihYHLs3uDEVJ0JuGDAzft6p3tTGHOkw4bjydMdTDDdxHMJWLsZ9tmuNBPiNW
PQw/AfL4ISGBnXkw3TpG9iOVJdBAvUKaJvfMwkTrsOTT7VvG1xWbLDMlvYt3I75R
UN5PcBWE2epi0gAmCYuoDdSfjezM7brSacj+oTDn6NEaftl53KPK/q//z77zSMrR
LGrSdZhB88T2AV43ztVQs5dKSWwO2DFxZoxbk0s8E0UfcyJAF2vVbrH3Y0Rsz/nm
PBFDnYHAC8vG4IiC/lm0of6bhpko+R30w8dEbv+rqBsD+ASeQ4T1XRvnGwAw/DR+
4YUG/ALZz2J4707N5HS12UWfWWaGLHEQV5Ih0U1iF0XJUwQY7poC6gINgS8JeJIQ
5V+zqIFa/cegziM+cN1n+hSP9aXAfIe4H5jvJ975p2HtuLlb/nquHHo7S3f4qReY
UyfCRkNDsbY2hTXCZvkWOkzWrEj9vGEqWmX34/3O2HSHGi0DgoTtXc1eActA53ht
VYwuwguKDJwVditdbSc2jSRN1mPNx4uWthhLWes8XZMIFpfd6wW/r80m4s6EQ/w9
gE7CvOrWTggLNMlNUKpB7cvwE45+aakEjz5Qa4SihCao0AHQY4dXhp2sBFJJPrJN
ZrmHSeKQfN3Id7mbrUU+d1Sf0HkzTiUQgpwE7HJs9qEftfMd85CzI+8U368jvtjS
TaXmOj/KPehLoonuYXKUIESUERktKuEzPhIWpsIGFap4XJ/jnP+NsmLJsrdZswzP
Sqz4bTxGIQKXnHNbtmE9sRLMIJxJmU4tEght6KKHp1HslPI+JaIH53G4AUyZUck5
TIyTDWtS7vThfajc+cBNnFiH9yCzLOVal9RKDOhkkys9m0aovPT+bMETOmGc7BYl
eN8oDSADl7elzsvFPgdOgRE6SiADkG7NCadON4CLJlcu/jw2qFHjQJ4H7Pjz4qZq
i37Uckuk5em/rsFRHzxgP3mqKLEbi0Xsxb4hMAv5H7r/zzjrsjjVZtpm7MShDZG/
R4RzKsLpWSNFH79NeS5Te/uq37RDgxWH28azTQq4k9K6mB3bip3VitAMTgaZ3xe/
yt4D9JjqzotDawrelx81hY2Oqke8vdJzWTEbrx/9oa5oMtIoqoZI5kBu+fJzvo2s
Yv2mXEAKO0VbSbXSKVTvXd3Ji2AycL4HwuNpMVP/vAtMYKs8f4NyxrZqs14OiOVb
gPa0bKQJKC4W7ky2+RHFdHzcc/qdEfdsdjp+O149FV1ahRYAgN3r9SeCS7yk/nvc
iVznGz1aL9Si4Z0xHCidTaXNZPTOxHHteC1GPuRjmqXdNb0WNt3lkYhsL3I6O3SF
NvcZZ3i8/1xt50P280qPWL+CfL8Sh5Wsy6TAUnwrD8DCVU/m6Q8041cyFQYYxT0m
8ahW6X/K5a2rP3G0ZvCgb87PTlk72rNo+XxuY9+hHqDzEKECP7RTVx+Ut3fB+EcC
xhrK/VPYz/84tN5fe2wyHAd9mGTjSJYSWpAiAzFBOhL/70qH5FXBqQqjdf+LKGIO
UqzyEEU51dE5sdK4yNsNT6NCpixwvkxpWi6wxAXwew8seVOlFGYSiBQQ+nRupikE
mdTavGYeDvQAIBi1imv1WdMLmmp6942ELuBq95N8YprIRmsjrOzLjYaWGNSjHCI8
Bw3Ox7phatTmwvRKoMnkuwfoysrKD0DK4oncc3MKaH2Y1dg2mnTHMBkb6CvYgGkl
PWfKPDMijTDMd0y1BwsfKvn5jEZOW0lAPYJHel15Nt1USmrAxvXnFI0kjAE+rPyL
/IOyCL7yDktmSISaL21oGBjKXZDfkrKgdNDAMFOyQCGNUy4Jfez/gPaTSa9turd5
Fv5Nc0E73uygnbTfogkeBFobV/+kruCAKmroCp5mw+v7B0ibL6Y972Uh/mTRbclR
DncoDwK/iYC3yF3Ut5zEDLTlIc37dYmOdOUIBY460XxLzZtxyNY8LkmsX7LtOq1A
jPW/CS4PQCgXyKeSVhWm5fzneI/wx9CoDGp3bL1qkbmcgqjkk5WLTlR2tsHzqxu/
aADXStOA4iGjH+gevdvJWB+FavEpL8XIDb8+SESE3nUIj34ceqrzvwVyLI1rxYiV
EPd1Lg7xb4CGRez11SYxeMgkUDXSir8u1kaQnMNeJ4XpHNcOYk0tjZ7F/VS9msRv
IB6wN1P1dpTb3NhJBn1D2F/NRYsNlJMcPkoTfETv4a92BeDVFRRjeK1OSxGb7mOX
qPN7vVa5v10ZWVXhZwL2e8s8QqZm6Z/8GjUan5A+zrW1bnnsC05Zaye68af9ZyfH
ardkFlmreCYUsehRtNV/45c2+5odzedoyQB5oapE9iIdr5DLOvDfwnLVKlGpRynD
NoVX1rkWN5sjgB7tHQTtZCNAQYWXpmI03GMXc7X/xRo0fH6MEWGNVsDnEAJAljes
JO83eLeAuMwy+MZXhkZm8DyAszVStOJATOyTQfEbVWbbdaQRMRYP2Fsehc/a5Qh6
nuyS95gLIh6Vu4LpQ7/GqKTOMqkdqveIO96xHuEY55lRHXtElABP+sVv6nloFh0a
UfMA0Z2xIe2T/Ixtz9bSPR/3QbVedAykYDI/MedXDWXCDifEM1jv1MP91MM7oyDc
7fVtu4IvwHk01e5zQUpanBLz2RlaMeqTpsGnIg5O+euglJ7QPkCVCTEuP9ShDPqX
iMHhQmzSqJj8ywbQOT2nfM0qBXJHN094F3cbWht2c6OBCcj69e3dZ0fRYrkmWoDi
4VZ6lVxnx+ds4eCm1+9vHR7ljA93Xf6ao1NmdKIebXKowkZ8JpXyQ7H4gkUvyLRs
UE/D2RdGYpZAyCNkVjC2PGHD/ohGIKkpXjj0qVtFSNhnhB0tPJHBUTn5T0DwLRIW
ilGmtk1+omyb7tfaJMtLeTAIARgANAK5J4BYqnpNk2gXKh9g8lzCGQdCnkWZURFd
GH9DcDbfoctMJey4bee+sBByApsz/5u2wAl+LoPejj0LNMs5Fky9YuvA+uNnCGIE
2uVBxIwsDrBoS7zSYX/rFpaMt1sPd9203TPyrxBIJPazGiXA9CaJl/me8nUOrX9s
2TyO83pCo5YQLhNSCw9P1H7N70P5HHf+72lI43PMncc+dnHAk4h6JPajxZacS4Gk
Ixyi7vU50zGsPjk0vRH6zwkVFjds32D5QYakdZdY4i72igOBlaqrPmwXgglxZo5r
9jMXJFI7/OUnEMg0WQvX4HHsNGfp78PdxhbFvetkm43DvG7FUR9evhwoPC4IgG8I
uQmF75f/9KkQOGaTjA/PpDZw33DUHYPmj1ymuDSke8tafPTHx2VwcIUIdqW+kMHc
hWXYJZwP5Szhmlxmsx2WycrRxhiJnvCJIW2FDjGnZJbdQao4KmNl1DAmurZBUJ28
Acq4A0yQzz620X1vzutqMiAapf5JWgt7Wa1j1LlGZXY1IVVZSG4yD0zezr5JJYsp
PW9+yGxkYQHVS8o7xWKqbhieaV9kAj0w7ZWO2azho9BKWzxSC6C0jqi0bOHGGDIs
iiAePVYmUwnHNwqt1v/ks26qOFbdHPJU/K+3uVzIB6t2/Bog4vIaYH8kYYfOqyJg
qWqo2u+odrWWcVG4BmUKmqOnvb5sr4iwZRYSzvCAbKqDEqlFHuF5OYb5VNkeB0SX
fH59bxL3Z1kgMO+lZSUJmoWg3BP9YoQpLp3YxyESfCQRu0p9OrqSPQI6bMhuIhhS
jxETQOfqdh4/djBDD/ZGkF8WBn4jXDQUfgywHrmAotoR/ZRLmarzON20lg8gvn7S
69+teD4XhAaMDsk7Ta0QaOgu7R4d/aWK9SIoCwRb6nAg8vVcuxCx2uTJ6vAKjkWZ
MZrk+901idVnoRlcdHhH/91xTgnVROQcEsKKQMK6qlYb8klT9YcjMQ9Mqt6C7Qti
ndE4lZ5XDSwAEhEoyVyzCCVQQ+ofPRw+t8eZWTktCw7sETy4U25kFYXMiJfGFpdD
o3wf8cC1YTUu/RIkBa3yLmdTlwx5I3NiqWgqne+iUZ/9rE1qby9RbHi/14ovkI9j
bjy18OGVcz/5a0jFhHrAHpROxyK5w2hHlNObbqgGUsKN/EmOYqMMeE5WfUWLe19P
C4hEAKVccDwla0nzyvcQ9BWMehOKu/jLa7/qvrwXhh8mQZaJGX2MAUL+vlA8/KXP
Z0y1prKgIfRQ/BKaBrn6e9SdxApRjIg4poWmwrZHKi2Kl3q3DoHoHPDquDVrQ9PX
OnOcwT+ElyIcICpW57ed2ZZJX/K+vr89oav8dvgacbxRGPTaV/MBSBPswpbflzuC
75xRQRPYgaezE8lRc5aDE9zC1osev0p+I+TeBAXBZ2vrJeXHgIQwigAXzQC+KXNd
dS3Drp4EmCD7H2YBqZwQl6lkiszraxP08uFdzeWJBzMgK8hJQOt7l3R4NMyb3P02
5nLxslq/gsqztnrBTQjknTHwu8ZqrBs5e2CWoPaLjdKKu6xacNUIvLjGn+K66+Z9
NrOp/jVOkVpu8lUXdaUA/1MatLxKOzG1JC5drfmhB9gDLeMvJu275rXHkG1WVxCH
Q5fucwYqBDO+xtWylnGoID21JA7VO0SAuWy6Zva7WLGd7nhBKp19wMPq6Qgr5hil
bsV6irJIlCjLvHoY0ARuHQvcGRd5CoZZ4LENLpbiMEe08FKCp/sYVH4QthsDjH1O
JGnXgTtNN5nAbsDZGSeQP0SgrunwvC53k7jHVyfifZbRmP2dC++BoR08uIDv95rT
SNLHeC3y0D15Ogb21TJFq0JEQmDoxrbBDrh50y2N4IUGpJX1ptboA9z3iCIg+Brm
KSrDv2+bUeGupH7kJ5pCKC1hjZO60BSTo1cOsQjG89s7SjqbV4YGACkCYJuqUE50
jcGTgTIGy/N70eClSkVksjS4Issq7+V/deEzN9xykaVuQ6HL9nb4UpqsSBd4Teqk
gVKW68ucKYtunpFevG4vVqwMd8GsVRtnJE+YsqnyqMyN9OS2+r0IonoJPWmhXCZ3
yzw1+3gxA7vXVOhEQf4HWdO0NO2g8R2lETlwKYi9Cinlq0VwFlxS/KvZyFoufzOP
/Is+GXnseVQvsFbbLzL7qwcBKo5jAlgC4jCszKJpnsXW9z6qRhebWMdHPdQD7eDK
auj4rta/CEpT9rp6hCfx8RbRbtQM/EoJVjOFq+cXQswkenXZ/ccsVKPz1qZ7rY0o
qFGL53ZvHrt1M6mWMXy9+4iutVZl1S2bI0vCldJSYMP099PQl5lmdXM9/OO5IvYm
LLM/luc4FM/bZBwE2IeBD5wssQGu+toTt1gU7YD0ijy6VPbEsq9+egpEb9t8urKN
Zxq+2Lk5ik2q2LU+IibfdjxzAT4CfUjfnLWK26BfZbJ255SQ8IEuEIrCK7F0h1jD
cXFTw04qjyqIhCvkpb6+IV/KDAAzkAbFahDsU+pTCg48hx6Q+fLadSYBxKBsWC3i
Ppm7SMfcvww/NKMCNdeOWPeIU7nn8ZyHW6qdbEGTDV+9KmAyNA28RB3uIugpo0Pp
R9MTrZV4jpw/z0Z18s+mKRIK8ZRNFnfVRu/nKFn8cLRcxPeyvkAEnm0DS4Dpvc7T
9zJYyxjNMmitw68Pj/rqIPbv/jcCAiyQFHcVCLJyKVMSM56kF4yjm/38eMKXtTQO
io3ra8BX+1yu5NJ9CdK2lGYY6WEOKHa5ZiN2wkh6DmfmNRlbHtIivsNwHaSn9spX
LLd05cu3FcYhSfv/Ph+V0GFVVews+U0qDFBrIyCTZgrJNw/L8IxjYwraw99jgX7/
j51jFkis3M7dJFJJMU9WzUKAphqR9yYHh8gd0l5hWCPZe0z3peaBvp0VSmwN192l
8CMnC/2imZZMmOLUaRSSi7kKaEJfkdI8xy0tlv4za2IGGyAOSzezdEcSlUWhTNJo
tN0h3FBqtLvSyJyTsKdwwRjdNL6iH8LwmZt9wR9Z4e78U34bMsV9tMiVk4PSJ1mf
UB5i1lKKpIQdpwwO5U3/nWOeE32B6sGpKJp08ZHclsoaK7sRhN+L09IsGF6bBcO4
nOhqtq3cO4qvxtfoO4z9UXJfMy6PP4Wprfl7x8PlWyKC+XkCkH1ux8T62Cq84gqn
MyzP/nou1N1p6Tmv09CGg8eAzY7hBvYYP4dgGQmFGa4/bISFj/6XDZJi+T07elYE
dP9pMzxi7zZAek4mosPNyZTRKIAOCjWic99O49FAtnOxhtjdfkc2AdXOGpRPT0LV
1Ffx6IlwCDdG1WRkR2bD+ADPSkIsdR9NXtWnl8clDpjid9T69Rz04adq4t5hgoyF
pXhTVUkor6H5my+MarP0DEmWD7zKKOkqNYwVjrIfHfAS/cQvZ9lM58avyV6HNKJ9
CrOPAfyrKT87loco7ocyX2yyCfF6O2vqwGhgjIsxtTOMTulVLWTuq8dILoromF0+
jo2bBkP9OLUfGqAEp5dvpUJVIkF6ZqUC0fETU3/QdRmkWlsvUf/UEPCYubxeDcLo
UPmnxWkJVElXel/8Q2mzKzaBncNX1KC8zzVaGcszI0kTYoG057XWIEBKOa7/3w7f
QO3LHH8la2QoDQIqHVHKLQikkc73o/20ltNIrabhMMpVP3UeKmdEl250LDFiTltk
kYxTd3eKQyFIiM0LPEQnJzT0MNdFi+2k+dA2p7jP2M+6tGsFTmyc98paKSwnHLoc
z9XyQFhPHHwXE5VBw/rpqbnsOCMPcwlmjENBv2Ft4VzNz6T4vEQP2lGuXWgucR6T
3Z/Gcc2s+10GMGFaiG586e3lBnkpywYAaIxYaRHZKppsj9muf3Afw9JEoCJtjTK6
PMVyPJilYASlrsj7mE1P97N99E0joXuln5DX7xXH50nPNomit4DaFw8Xf2TO3gjp
V4f1AMECpwWmHFUoilY12ui2wSgP8/IvPtzI9mzUoT/pqqxUvkg+vBEp1gGUZGQi
3mHcwTntVsx+4v69odtQKAj07M3Snv9QG0G5mf7/Cn/tt4e0pLq5+QF1WEIYXZ0x
nGWD7J2b++nxpiMYccgUYL0hjeHMnQ3P6vuxaxPE63y82cPzIJiFVNgLIK0DN6IU
ZzMvC+aUHgU0VFAR2ow7ySD5pTVLeEAXqt+wo+sVKDwd6us46VIcMWKOY3K/1xhW
AeUuID79DrP23UdScM42hVxse3PF52EWC27YiWiBlJo3H+lKof+WNt4tvqQMrXU1
TEunucPWSolxl+NfHcGKnkGaHmKU8TnU+Mnr18h+Uo5kRqwIo4FSnF13qohQZyGq
CdzswluZ5kskbayuSfEPdr+DXTeZRCO2NxUtxQmqXglT/hXm7DwpzgcJlCt3iDCR
49vcsIrSRNKqVKV9JewoxxESuW6bB14XoXiDddAeFXm9Qj2w15YhdzPsD8YBLcI5
pM0Q1XHAYx2VKZuuxTNqxRJV6Ia2Yc3+rLV+0q78q7gfXTvfWJgjv1sLDT5eNFF2
FHX85acKoPLLjvheghbQ8h8oaIiKdM7sb7X+rqAFkJfOXfsEK1S2ktx2a7YKoqje
2zN6oQlJHOo5qu8njLXMoBu+GtJXj5tio9pYkRdsPgqvjTSCJKpphkztO4NARhFZ
HcW4gxKwRjvrdsJud9vJ0fP2DIFByDC1/3qWFoUwSQLw8ZhXGM03+xn+lG94gls2
oVroHmw3aTrVfnVa2umon0L3PEcaL+PzaZhCW90lMZgxi5w8uApKJ874bfk8Y62E
42xka2V3/h3CBd/G25wzNjjTqRzJrBeExSXSBtvAehxLQ2rQkifT/Hip1xnperzb
xYCh+MmrGFDYwBhPGy1KeZPCgLdg3wPlPhOFz2RCw4NeDc+lVruyJp5aK/3GqeqT
Yv3E/u+eELOCgMIVHI4pselOnvosCE57entRj4Rzntqj8aU7Ut0KVCUJUvvgriig
rgkq8UfNzMDjVRaderS0gBMjeIqmHRNWgb5lEwLSjTRI3uuOhTdRu3s/w5YMHbYG
df/Gpi9Pe3JMxx/O/sNGqAhI1yZvLTi7sekPzSp498jI0rqw3uDwUCGn9ghpgMUC
5wJTYotCdZAFZam4s31n9/8rU4f62CEGczKRyeyZUA+h/MjijwK+WI1uLk5yQ8jL
12DhD7VdjdXH/jyOX0UK4u41z3889K8AohaSXObscU0vmgLKGoyktnhyGzZX0rA8
IHo0BhXeIFEC4485y6uhZRuvfyLM64Vuxp080tu1Jl0t3GfiNa3gswos5cL9UkEn
prx/fAwiNo/mQ0zEkeIKcmsVCurr9Z+kbonk2oHPRNYRCU1U2zarXr8LdQpWaUPh
MLyKnSJKyVzw76FaORxqI7gSD1ZX+9qmMo3GN9dUrc2Zkcpa4qN6ENwNcSMg2Ylg
lQ7f8FRSFyIi0IWRKo1z8s2v3TCKLZBFQJyAN2xPagxAEF+ygD63CGkCjXzu02Wi
XdlpIt8JtvFqnQt6FgJkTDNbe8poqdQ5buCDYyaexzdQvwH7TDTWDI9mnhV9jvFk
XdTvhTyXf6vFs8YRgFAjo/oKVpgfa+L7jjD7bfKFShueLrgwJgvUguG4jLfsoLzx
jirjkm5V0nTMUgnFp4wK4q3vHRMnWmVO5UP7SBoC152o8uohIDBtTYpFBm4lY0kr
pXETtxGRZIbS75JbI9ZXK3cIwoNjGZUybOHPAi+vhUlQE/k8EkVuREOQ9VGNUNnB
CQJlyuJt9i49YYdqaGjqLk3cMnK5sfov/pMuEM58oRSJRZBBmV/opLfIHy0zxVvq
1zifH/e3jREgPutIpifmJ+M/yEyf50uslZa4/2iazfvOpDVQcNePTome0w5tlcoV
UDkxlIXrYKmxvEk5c6RDQXOHLonAaZTDsGam6cIh0jQ7cmlazQmlzjMSh8XFEQ3l
RYlkPWcO42KUvhHAZ6Me9jPWXv/f1i/FSPYnO8OysB/SG0QoSGyQitDPRJJG/zUj
AQXsJZzbM9XN28VR0/MIy6gaEsNFsUu44Aifu5p8mmFrr2KCuXyK7o2nq2XAf0/I
+pNbzZ8jHcz24/Fe8sZTAypiNI32qSR+FpWCVD4Qg37V/66PA174ri4UoMwTwLwW
BIWdfBb8JkasPVsM8dP3r+ZVfz6XDpJoGk31tHq8Qie8Z5QvuUooxQH+s2NXNGLo
6b0H++jtW0m/jlUMIZAU16Lwa139iYGKymPQTMRMeIlL6n1Uct2o8TRgKk/dnGLx
fOwSOgyUvl2RTer9uuMsm/GbrDapYWpfWkG2bxdbMIMjlGt5Or9OOvCBpdHeA/+3
rzR85LkqxZD5j2lP218eo/y0vvlqc/VGETLN0XSAJHxQHUMFuqgMG4j2e5Z3I0Ri
/d9cAPYWOIqkLBCIb5IX/UkGVlzrnvksAjuaP5iiGLtkuX13nRa50uVx5Oc06e5Z
EtZDrCW2gcz08E6jMEmIsiSCCHk79ZgRkycczAmrCdNGGE8zvR3mS/0yr0fanbqi
Dm342TjmlViYuOCQ8J1DgVNJ3sX8yjUlGXGZKRBF+kOm/oCJY+Mcb5eYsolgJHp3
MOk0yKxm9nygL6KlDwXtM0qbxHKFoDSf1WC2OhzQZISkiTaULz17ndooBMWf8a0j
5pSQKaa+SnlXmzZOgN8eFfSfifx9hiImw+n+L5iKLQkXKdkEBi68MRZrPVsEtvUi
dGRDI8p7epvW5o2Iq2eQW+K15cIZ8/vvuoAsqsBq+CSo6jWBJmoEzY/EC5Emohst
xnLqPBFY3nAuyLwpH4+vePAzgQldP2VGGZGFAGCmu6R3lHTacXWhhPx2Zc6WG6TW
YcCZ9A+15m89dOFqheEDc1pQ2BHi8sNHELCvi6SaKNqiFm63tf7A56dNRe3uIlht
DxhGPAx7xbnV2PGmSZZi8ghFPNNi+Cgb4QNeIMq4xi0nG/JALUPpxOebZSsz24oC
m5qN06mPYkNwiDxq2b3SM1bE5BIfx5hG/62lsTZP5jMFALWngXms1wJuKZyBgtd2
xNGq7btjwJKWGl9sbCIBgg07YDCwHJGFiOEjtLubpvsFN/R1wzJXnOF9jF3Yuqby
JgUzVNS9raUKWJAmbydsClb43Mo6KHBbTdeG7GrNIUjTdFZVjGpWD4urFD5baiDW
5j7y6Ab/BLXIK4nXV6o41Yuhqqf1nBpG+rGQFUTKG4eDwFVokUr33xs63fVUg1jH
VeTNSp/61HWLoD1wvMAHnlFW3BMGJhbPePmANYmhAG0HlJR+6yEc6jca1CSaxPbM
K7l1RIoAHRe4XLLC7zbHsXL54gE/GLirPXQvaD96ffUwAlRUCjFe2sCbjzNYB4CF
2Gxy+qHIh+nMOg7Ien6PCMDZS4N4fyk4aWpal8t9S4D+9rBYAHyiYUlCKJcZpS5A
9UKy3/nxj2zvRytGZn0kBt6aGtt68/yyu3JjiBLkP83H22I5D4vBsCPXOGLJDEO9
c9KNnY9wZlp7RRbzoqRQN/sAxaq+rw2HMQe66On25Hm0x/+xwGs+t3BfsQUwcRN6
IV3JfAq2edLxITH7OhcJuK/1e48qrDNIqIPtW21dP5p1xqR+bCuRrLBGV2JF231F
Tf80sAAG0szwv3N/KACmVxRLdv2kFhmUPRm10nKvnuCZLE4e0k7Jk7bBbkt4VYzz
jJhcJGtHcKOKaLMfpn5yHXxxk9RQoe2YmEfGHnkBxsIQuPP8uopRbZnQ29sn+o9k
Jhh/5nWNKxMTo39pVp4sprEym5th0d/oZf0HTfQ9Pz+4pOxfRVfyN4PmSO9/blO7
DxiQ46qVeP/I7bB8ZGGr08kcXcAC3EDamqCLjFCKJncav9DTJpeQCAM7ISwfnEn0
WDiavoWXvzxM2Zm4zTm9zlemCvDzP/+t9rOssyRVP4pELKmkXWbEK04/W/dhPEPo
KmNz228NF5y6mUdlWVHFHx7L/r8wiU0zZ0PuZqfKFTQq2y7vTy8aOJgLUsZcILUm
yCLXIKQJIbxvV6TIhy8xtBm6aYroa4cCpF1E2FE0W0eAp1sItoGvr9gt55NMuJHN
ssQhykjE3xqmo16tPl0csZAZ7VlGuBgmVsfUYBZN8cGn/O4ifmnAzFibgJqi5cxf
4BYdehUM70juJ6/numljfps7k6nHkOLrYSguSUnQuzSSZd0L2tXqj6OYDq+Kyk7Y
kTCZ8gQiK5/8BA38DbLLKD7SD6cB4II/K8LP10XXO35IM813E3+4CLMqTWz5mTvJ
hPxFMYPJgFpWJQjaMqLS24fpF+mW4mjiCLVtwNNFns9SkBOzh1kVxvi3dh8qNGia
fm0Mg1z2S3H5EMhNneTz0XHKx8kbAyUQg6nMpJRBd6zMHliBKtVKo/3mrr/+KA9T
lp6zwFJmneMF3DaRMyBltlPnI4DheLLw+HyK+v0oI60/yRHD4pgxc0iZr1Qp2gvp
wdqg49BhVefOkFVCDt9fMig9IE3idKYPON17jGTZz7KuONm9JGzj1LqmRHTmdzHN
o/EMVpabM2/x1P7qHPdCxlxS6KB+8UG6+24s0KYpoQxDuQOJhM393GuIUUAZog9a
312fJGsmJ9m6XHCtlaIwQ3udd9ppDcw9b4hRb7poMsG1/OVh4kNPgEw4KErHooKz
WvkiKVck4ThNsOfNm2QyVSJnv+p4IjP10HMNccqAGCtzTxXf3FohWX1LtBUHTosI
IFr7yetv819msO8WPFrFTChbty4/y4UaMkdd9ozgDkKYgLmvUGyScl1PkHxtV93q
741EWzQEyDr8xmq6ulz9pyZVa4M7zwYfYt+c7JEI5uQ8n3+cxWSF6VCcnJnY3zbE
jRmJKMHbFphKnbewoqKUAMx9AWyK+S4FjLW9xKel6oU1lc5N4mOtoKBbwdv7IjbF
Q1XgLZoX+MNcgUds4P7pxhXMN5XNPj+6jiaVogJa+yywYJxTYGRR+rx9gl/BCRKS
7WY77yAl6zoiTIVBxu13GtOF0nSTQiTMzmby068bn4Y3CBKyRZAWsOSH52ovV7d5
uHnL0p0Puo15CTUr1kCtgim/JQNE2ypG5OuXyj4iMM5MJCnoZmDaPNsX87mv4Bxi
/GTgwwot+C+OyoQ6CLg3vYnOm+qW6L9HYPrAXuLXMBVlhuYpX2CDfYz64/W42s42
JMAvwEnVmQM2nkfuyepPCkrxOyC0s7S7Jj6/4qkAObBXgT8TP9er4TIZE5WBG+mk
WMuhEWzS/QHtHUMrHpVPTjnJrePJtn+aLyr/zuNVMF4sg62RgAhP5AONZkJf51K0
pUbMZjSksDJVQyLoFgZV5iwTOIojFTV0ZfqzQ2e0h6HdRGGh4FAP7nzQXjkCTKda
WNE/2jcNaoj5uyz2a4OfiD74SxdFDvVeYoTFnwhYY48PRXQ71Zy7Zrw7fol/9d4J
FieLBpe580zc9fiNiU0Xwqu5HYOAl4L/7nV2AuKzqO7YwWhjlMhxZVM+bzg8vWTl
8avAK3NVmjylKIWIZGLj6faUMZz9K4VFmE8FWpzAyFaxZmr+o/5KX5xEpd5fwiIG
wzdcNvPGiSiGl2XSLguhj3tAbx1vzHzsY8IIJI+3kMWx5XYnF8T3ezzAM0bxK5Jx
n3FtbcUl5a9rU9uWzPSLazHBpMdkiA4yl3sqBUUlHYPUVeQgVONqFQUD0IZS2oH1
8dFmRJco4h7qoslrzxI1Y0w1a/u/O+o6rOWgC6cEcYgtRnm3vPpIeOCf70pc/79a
IdgjM2WPtyUyLdqMhOMUOBGKpUQcPZVTP3NFq2HIUre1HmhNe/LAta3DKXflEvJB
XXBW81uWeBFsts+TBs1Sl8l42087sAIE/BDp6DVWdnQyxOqdnE3ed0uwn7Awu3Wq
TvzenDJAxYKAnh3rk36sTlYOzVgvv9NPR20Mm4VUuwpmJFNah7MkKtX47sAkKT4Y
RwV2gsSl6OjiWkLqwd473v1VBaIJyblwDM5o3EDlC1a8P2w9arzQsGDNEoEAR1wR
g0fZIKR/LyBsoyT/N93QWhUVisCZY8nScCzx9XdfGQ+lDGrbidXsNu7YMUBzt0kg
1N3GetN6BnSteyQkSlRsqGqZqTTe8tE0mHuL5ZQ9jUtc46dA/0gYZmEjjbsLcvxU
Wy8EvYFOG7ab0HsvpmOFr4Kryb93nzl7G3b88rnCQzo/eOcO7fIOcptwKoDAPSLz
fKG6Jmm8vTvDOfS4rqQ6GgLc6DVptebEP7X7Eo8XkXgZQjXVcnXk339Mxuo2MnZe
RoR0U5etHYGLaWujNWFYFY6fvXsCX7BBgIRWHMnT5D2fSJr5f3/2b5gyW/HgIhYi
yET6WuQ6D0X6eONv4TUdpquHZnfnfCTRJyBptWbMKtKMnznlrOdYAsLNxI10BC5d
QkxcQgHSYGx3cGbHjO01fCBjp7q80eSaMaUygfv9+XyN0rwUINgC77tbplTukZ/e
ZAY8nRj72cYjJaxje7i+lmzIJrq8hcImuk1Nu9MUtHV13IJCIjeg+GFNUnul61bj
28l2GBP5+4M/JPztv09+tlxt62FEUYrMy1WkMGL27SALZ//yNVz3dU9PasTkRhfI
4R0vQdchGjKf7J1g+UcoZktXJSMqPkcLzP7tZ5orJm3XxI2qIMsoBHiM+ZY4Nbk/
ZvQxQUaze9hrfzfUclXLN7l086ygIXD/36uD2aNPs/KPpx9SM1uHrPCV/5Z65oN5
9PMPf2kqhqGIL/nmIeiUzXej3PMMGpz/QWCfgI66Lgwr7bOwE8/fFSPcc3r23wlA
otFr4PLldFwYQXv9czRTETYTyUocHWce7TThONHkAJciTCuqCQkGVBFr1Qerf2k7
88/SAaH2PT7oDbnnULJS0ejIeVwWMFsI2J0H4ywcfkyvCZjAjukW0qCIUPzsaVDN
hmykbxaB72+ArV1EQRsSDUCzCAMzF3RQzafkfzXeJka/edoiv/ZEGzR+Swk8HtVu
5RvxWqByMt8WYSLb5wTxFjtCq6apSvv8fOHPQ2PmgoXgFprfLh74nPXtLMn416ZH
ScVTy2M1fT4yQWErs61ff6NkW3cSS+31MdXIt4Tfe29xAOq8XyrJ7bYju2vRE2ak
Yr26Z1XVb9f/6PN1OP6YGjWRTcJty8jBgEtrQTceUo02m1W9YvsGtTNWe/IW37GQ
J+RdcxqxBdaI5TnRpxAxjXzxrT81ekHbCQHoIaNUUqtLKJIucOsMiRitm0bAkd4s
mj1HrTUvjmtsn83DzmgFLkFGqZscZ3ZAz08RjqxyDSDbvQdGtzGOkP/k049215pj
vhnNxWMxdBYzUHXV/wzJS741E+WCK+SGlo7kDmNP+7tOLgLgly7HjqxLKvRHGGOT
+a1pwcApwc+GtvRpTSHC+dJQ6ZUWfGON6P8t3A3Uh9/Wk0V9jr+os9xN8NcB8qI/
sVjLDiBJwwmmJWTNZlf5ts8ScwBuM7SNqAPB1Hx+OhJj44zS0bNbueJShark3+yD
6l6XUTB50cLmBYTcEsf9vq+RHB1/1ErQfw/n6AxqNJFZKUh1MSlB85jD9Ehaao0q
Hu8d7/I7AF5NbWxcXTfel5Rz7egq6dHhWXvcKZkU7pStbRD0osn3Z6Ifl3HH8t2H
H+Pdw6B98i70fnXzc4vhnKNX+dcZKkzdZ+qpMlL4Vna7yGDKXEBvFncdWISnzP4k

//pragma protect end_data_block
//pragma protect digest_block
FfVQkzWpK+i6QV+sqhs4ds2APaQ=
//pragma protect end_digest_block
//pragma protect end_protected
