// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:45:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d0AW+gOjxaxyh8HeA4yHMG4bPJWmT+g6L0QTgEG5JDFIcQvCBq1s3sUrmGjgBt2b
8eUYpOefq5XZ/77n2kOMfi+766Eg/LejoN4QaAMv1HJHsfTB2az/Lp/ETlYIJygW
1R+0v1oo6ra6Qdrx5Fw29icXqFJumIGpTfbsVdTF9H8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
uvscfwZJEQxMse5aZP1TRBxuX7T4WAKsrB+0fGR3CgJTSU2xy+m7Of+HwoN8ISb5
ytz8UCEIb2RpPmIz5W/1UzNGOPRzP0sjSalDBGXI3tD3t0c6PS8wW/NvCsvbKjfC
hYrxpxxmPSsrMYnk/dgKBjbnvOWyaQhTz0klSGp1QiDpLuFIIE1F7WbHfrCSFOIP
dstLEG4OMsz/v+aJusaSDZVFUgyTLpRRzFBpZeGC5v3zK6V/BlDIeVAb3JR1V2E2
cY7cWXUg0pNQ6LmLWyShDB8XgQjTFbwKDHQNfQtm2FjDS+F9YWSTUdi07RLx596p
f8VVeGGff8wxnfQvKhHCuBayjsgOHjnNoxyW/BxYhj+r6xaoAVl/eU0rl6dWoWi7
PaBlWhQl83Eh9YfDXPrD4uKIjP5p5ko2QWa/DN361PWs/WPSiaue3Bdhg7HQAGxq
yp8lbPm5M/LZqoUY+S+7qC6vAuPNuSGQTrJ23O0T3U9QshUBuMpbGM3GI5MdVrjL
wLh6sj41DZCHvvfngq+KPnHsvSDZilOXWiGG+kk63873W88GT1frpZy7ECXUtX1q
Rbv2zwKolxW4uYWg6z9gS/fVIY/ndWtt2U5Z7sfNaVfblO/s8pwHGXH4BrLjVsJu
nUWiaze5XW0tB7VX4vaZdcG7GfS/iB4MHHhCqQQNvlNWTYKo0uQXH17kSKy0GX8O
WAIT2rXoJUZoq9fBsTE96UKgUByTYJW8ZTgv+xDJ66O608JzYMJzxi2NsQfWPryO
Lj3rgBYwn7p//IVhzYZxeENrWbtolgzbXAMMUOHgWVkHcEW6qGWV94Hl87egs0aK
N5hvp1OQ+nji4V7sMXhWLgY9wFgndFNYljiLWM7EqWOhL+2u7v/Rr+x4ZLXQZF2m
A7saQfp7yddb0f3yA9jlqLRtNbSasXOlPv5+/0fmXQaSSJXT3fuUXi2HN6CNT5Yw
MS6CLcCBD+QI0OkXT3MoC5GfkynYrKXqSSNvkGDeDyD+zUpgSvMr+886lefNu4G9
sJwl73SELsR90k4kehmrxTuoXZ/3SZMJh0fT8l/tGJUndj/2En0LUR4FE8vrVnUs
b3oF+HikZrrwrAKuYTr8m5uMaB6b1+9MKpUQxOVFl229NWpzVXa6dguAadFcVTPB
yjxjyCi1g+XrrQvyUOsK9TcDQiptUfxidZIpv9siQk2dJrz84cwB4GEBT142rvJB
cCsUk6ao63eXOO1kwkfjPrmO7Q3jKcKeCwYdNmtk/Wkv6WaEOqlpLPtsFYojij4/
R+OqKL1PCksDnnZVw4AcGUANK76U3ZIAn7702FK1KljMdSoQoATzHMhSxaSlyAyZ
b1y6YPOeQuLPWMD7H2ni48pcvQWpV+Dw6CKk257k8BGNLmpyDg2eYxK1KnXw/QOw
jNVZEWTroRaVJbLdtaoNCoilJxRRQTKm+ahI79EfXCdr0vuSGP+IWl4qDisD8J3T
XlIz+UMU29ljjZP/JkS5LiMctdMcuRDCRMurdyPIivWWNIca0AMEFypGUxr07Pvm
ZYrVY0wipmXcmRhkypNbATCrqF8fIEKkrCnpRUHVY0FCmdw+jzXryEBL1G90k7vA
7NRAut9glPozMCPVWr+sW2DAVozlF9TQRVZT7cpkCeqYapAR5NB2/PbF/pGan668
6S55jJtbFE+8MQZZs/3OXEvRtJGlSLWA8iRu3LJrLbhi7QA1YnNeew+sPX987GTx
5fDjLGdj/1//ixnodumju1RGQdz+Qoiyl5fXj3TGk/nWHr0bvm7/+CyekvzfxL9b
Bw77+aT6lEXqCaPmiXExJNni9WtlOiw2GRqQJCLmDRsky9tCOuhrn51ptN98zAvP
XE4zLRZFu2robnM2Ss5UaG0N5OxglW1Ey3RMDGIFbrWqXXs547NkLZvfv6wAsTOj
qa65LQ6O2XhCllrG25JsMD/Cz6lEHvqtKbU7L1Q808K/kZwipA/efXHFXu+k8yDa
gU+SILIg/k2K/mKcLoc9C05Lxmo6Piw00pe4igOgbZZgFTXbXvSZ4GVf+GsXiQgN
B51Omu5yPMcvhBXa03ART0WxZ/qjEZat5GnyGjMowtVfD8ajGJEKIj0S2zbVvm5C
c58HCuiRl2wnlnZ7pq/VhMiJ4ksYrJgzBgNh4rLPn4QKcr10CLlbAS+oRe9nED55
XPMK5FdVvjPVmd+0O189tRkWzqtDLCta29ctXQ8Ndc+U2gUiSBZxTZXtfvgf8lOw
HTwJZK8iWi3GdNKHJFOEg/RRfB9uuAt2rSQLXtOUdcoKnZ1sUDMqFLoH8TaI8XXk
c6LiziZKen+0Sof7iR/vizWD4UOhm5gl/YcBqIRykwCQbikEbVc/Y4dyAkETuSC6
9TGMAL0LvwC5XP7/urW17aIH/hI29FeM1Ks5XnURzXBg+Wb48CzmjF+u3oB4+qpv
zeDLCH5J1zFTioDIiAT4Hpz7xcQ74D1tLyJvaCBdR9RiNE9i452kKfmqPNopQHxZ
oyXMlHC1IGVZri576X2OI0AUKK4Lb9O9QcFixc8GUoN1wSBUAQrmP9wX8rE9zdG+
Jjz//VarLp/gcSrvtZhhBXkZxsCmCKMizlbbdovHYUWKGaIpzLEyfk76mOe2xAcS
pVPY4PUTzLac3Rzep9OPtvTwBd1NLQ71u8n32UaM4DYYFs76PAyB+vL1FbjBQ7dd
Laaumj/ptLxTREnhujCw9eCR2kEaQ/lyOt3w6VHS+yBpTPuyh+dJYk/vUTbDr9iB
wQCw09AqNYyk9oKicWshzPzIv95mAZ2djrZItaHQi2MkKGEhubxTbvhRVaNtequ1
xOCrBtpgT9uqr0S8PVtQpk5GsS/PzsEkZ5c2l5OM1kPzB8h9kqYIOsb/JvHLBGUJ
Rn1RYOnH4m5aYErX4dUoZCbi35wB5i8OePIdSKq0cpFBH5m9hYB7i0SIKxw8+G4I
x0iwGemRxJd1mAGlDCiJ5QmuM+9Cifebk4Opc4ZkRmQXJwfl+3+bqZXbvAWuG5fe
XsKajqN+WULDMC52JNc6wjeuDN44RtymZX1l3w0kW0eLeAkVMhjug+TJdcp9BWdo
G9y7GeVt9PDL+h4qIw3bLcj2p3061orMQIVsLTdefmjF5bBUX0Zka8bLSaT6PQBU
ggLhw8QnI1CORbLykzBnybSuACKFHcskYhUv+WYw8WPsF/BnQcU6B8fZdGYyUx2k
aX/Vcs5bz+PcT1r9/XF98gRaNEz2Et368+9hRE3RdX669SnvlWEuu8mpAo3ReJrj
v3QBcc6PKg/ZfVMbNXsNSIcsDoJ468i+ivDhfJ4XVm+gASAGcM6yjxVjdWjKTwOU
2+4vfao7dZZRLmk2BEeYcxsnYgF8UQ06Kp2L/DNpRR5b6RJjfXB7BuSBoZCPXOsy
kUMg1xp3o9q24FrsYHzk4hpAtiJc2/FzJzF4OIwi7KuU29be22lwZi7FAwLwX/UK
sblvFgp20VEOXzAxkHjOjeqte76hYOIiVBPCTVSZFLPTDOvyViZepmfp5P2BR6EK
pORvXcOXyjKSS/vCOswS+CWqU+8jpudDotXuL3F6J8Ir4ezaQy57KhDvCROErARE
0GP83+ZJBHQFCYiuMPtIGzpN6Pfq9HtQ7MoTr3vsGXpKxmaElK2sjK6/5bxnKF9W
sBgqCzpjkYMsZf80omjQQ27KluJ6S9zYzWKeLkeezCd4miufb0QHmgUSdUADcrFi
nHqM68VmaMoIA/V0X/zjg7XmP9kILk49IVXwjluXU7F21knFLh6hFwYs+XKKlZgr
zgsoUZ0eSUC5qddZJSPm4pVLrknV9GlmTL+vTtrEYy8ZcNZfWhQu35q3D15UNyUp
n5Ow6eTnz+G3vms3U2+Ol7Exn/MwId7yMjVZSgpFCBRlICyV/09dXamzbb+OEfUe
X3WhcsST1NhoWr9EGo/nLTJdOABeaMkV+tbO73dS7GOKnm5Iqb4h+NsPYpZlavLC
BX9UgyRg4UeK3nMNEeYFzcbgsCfZJh8L/PAHs2hooTX9DTQJrax7g4LXzHDf2DXs
ZAUpr7sUuvrBU5z/2T2w6gTm0L19Tdraxc2+qtnwUp2jlK0HQdPFmP/DylD7VVe0
LcD/jtkTV9PTiWnAnEwSCA8lAmvsXvfsrCfcGfC5prjRg26yP9AEkXEUcH0XRj8r
83mmjwzS5Bu+gpZb2iS0s/ylk5c2Hj49e3yczjdZFeZI22hkn5BAY4TeRbYpW/Y0
a0P+ZVxrJ1T6Bii5/zCGN++tKMMbNmsTixgL8OH7eBE52gRdoXkyu2Bi/kgXo/Q4
c2RjjnOp2aZixv6PeuzaQXjP9h6+eiCaUC0GCf6RNibVZ3CCcfA5lPwWPNsdpiSk
tKQWiZ/V+D6QjG8I4MrxiQ0Xr5L0yQgHD49mG0QwLzg0m7ghZsvzGfiecSb9311y
GIfCa9PiDbFpoDrqPwye/6OCUFfXoqCf5+KJ2V8C+iAVaLIg+zXTDwy3gF96LTyB
GrLu14a+j2Kzfj7bIHfc0yLYMT3voyW6XWAGlt0zMWECrO7FPhEEvrUuLD/cdn0V
FtkhRAnhKg9gHa847CviTSn16I5JNqOHwCiSehzgc8dg0uZhtKqEIKBsywvw9/Aw
fR0ANey8XCOdrq4MgqaooL81u7nS6QOoCm4QcUrgerjYBAb8NeqH4sS3LTwJ8tZs
klqD230EVWs4nReZEp9D7WS4YsHAxOwBF6ZythZS1Ecx4xqr6V77t8gr2iYxWAnG
ttLN7HdW4F5t53Nnc00ebZXkZTFOTqbVyBTYuGcr92fg4IoXkxaDqDdKKVyDB0bX
eL6Jm++e5FnO03VvKFIvyYeham+CA4Kjoi70rEKi0PhUSiradU1fMHDUzYDy3ErM
hE1t9f43/L/uR4BCUCgy0bowPqV6wDbiZE8yl7i9MDFzm0urg/mm2RDP4pTXdHT9
C0Kv1LYMXOVj1NOuKd2uFkarqbnuLyP61N14tO0XhF6kRpwt/yWdtTnpwiUxv9Ar
2nShApl29MolLyMKJ8a3jbzcw9rSJByf+gBt2zFEX1PwdWcxX1QHoAe+F3b03Kt5
5+B5pHotoOArau03y744l3O79mUYQudwj8vg91oBxWbu6giyNDEACZ9exZO5S8IW
4fWYVOUkQRKayvRoKRCnDNYOJVGhCNvEWjkPXMO6TtMzG6Nv75ymPQj9KEFwxxWf
orY6unwwuPjHDyrzGQpuA7cu2uEKgKhMgXX8ZvQKP/RLMGLfgycxAU9jFYUjHEz1
u3WgItOS0BHmoQGwbTzpxbumfbPYmdoYnpmZiCL718cGhY3QOeLkZyT9Asf6vxhx
dSpn+RXa9/rS/QSX+NJFFGidUZCbDTSHBGvu5+4lHj+X7ZhZRtBWIcn9Vb4Jkgj3
+frjW1zIBZBfVV0IFA8WnZZGafeikrJHy6DeQqJv3joWxQRRCNDz/bBF0Hh3ndvo
lenLe4jrtnGtc7MVgt41H5w+R09/pCWSB8jjjbiBfCSd4V6SLaWXrhIJ4tg4V7tI
OU4qwJ6fYhPvHfUahpUx9Gectu7MZeALUu4X2paKFZbfrxdlGpbu7rFCDHuUE9lW
du42VAt+FIHH1hrEFQ8fRwqOZGSE+2V5dguGQjyk3UduX1bVbbcHtYiy9jNh5r0C
goDJ7uVwn+NROHEHQWG4T2otOxcIrIEm4ynGsVFe+G85ePQDt88CIYDq9/ZhVxTT
iVYGyIIuu2N1DzYjT4iHNoKae7zAD5wejeSQna8kc1pggMUXYUHcGKTM0Gzh1BiG
TheR/ani1OMt8pdOxLMUnqtQZ3+14vuswZEVqBBfIwiTVaojiLw/1oR5Bmi2DMRX
QUpFlJLxvXIUt+JDA2OeFZXPLWJGPpiXCREL5s+X9y3y6emst67ji6oi6xpmYAMV
H2G7KlrpWHSAK6dsAV5WiFPPTv1n0aBenPHv+rLfmma0A6ZOFmFs2kvPQUsi6W7z
D4nrkeTFV7bqLGZuqQVpoJNTM7DbRFVxK70coIkH+qOAKPwmnFL9BmEe3QKQazow
FLYVwzlJI/mUXwRZUmrc6DJn6bGNxUMffe9i2pnPFHDtRLG4r/BGgFAyemAiyo2p
/oDYoN2LJ6HtWLAa6rbT6EOAja/BSEggpkzy8O5zOnMCiGZLebiPj0QUIwu8mtE/
C6v7gdoIhNl+niPdrt+Hd1E9a8fRxshHB/we0B3/kaJIubQQecilU6vgeflnMMdf
tP+O5FQAZhxeWxaCjlnKHIghFSOV1seWSLix+4/4gMqgxmOUmj5R/KZfDDHpKC/A
lfWqHMgGq6xErJkgH46Ulezd9LhldGXNT1NUcHX/SWrJGZdpTvuvxgeu0ho/ctDp
7Yrm6IgytdFU8HQ2DEGyKp9ikIdIVYk/eP19sPnmx6j5UjG6wpwJQ9ecc5qdFy7w
Pu0MvTEWRZ8e0VXRjaaxssigxn0YodMUX4w9PBS7IwlKIQNOoxSUWfxujzS9+J6c
xJcNkdqUM+Y2NxksvC87gmap+BMD8qta1Pvcb7CHvMUm/tnfGGx2nLaylhoG9U9v
opQzQmxps9DIqlZIghdXENm7EYZUsYjj0QvToi3gm1eB7YNIrBVHAgmhXz0p6Jn5
b2YPQF04kOhxGS8Zwp4aZoZVh+OI8Acl/Y5j56eiXVJAzt83A8ikXtXvFxfXUBJk
TaIVy0BNQ4rwc6v2jkqnOvuadAX2sPkaYfKybUPpCt77oYyWteH/aOmL51rJ0hCw
HHrOZKNAwwxENsfZqIgLOSVv4b6CM694U6d1vlwQJyQRFRwllLGCvWEXJTCwqUgJ
kB4TOXHNmeohOE/5EM9MFzCtjoytfKPdTY7DDzE0VGbHMrYamGYHpkqvaUeMOF3J
FA81+s5rSXJ1A+VXzHSv0TSFhuuPloOSY9cQL7SkB41kL/dEGs7/qnn1Cpn2No/g
w499BJiaz1J7l/rTw6Zm87TByKOsESxW9i/jvU4r4vaBDVGNM3Vo1DFih9Ow32yg
M7ehReckGE/wCL4RfsLlMJ6KL1EvimIq5hyYugzpiFhdYVjx2Wypdk4xdxJxIG/k
pmK0dYCeZAUHhl+brxQUGlkQIWFFkoFv0UTG5ZZLvfhVGoPRn1dX+BfwkVB4CP/j
oBSwVrBQnX2gJo1HabPLFW63IokQvQL8dD+H8bf/rljfHic2KE4PvZtV6roOqoua
qSmsNjC+ShGTJDKqdjiJDQ2MyLuKTcpF1XcEVtFy658CL9NEkmjHzuQaRbTMjg/D
HnGzOe8F4e1CY7I9lkv60eCoRzjesr1ttVCZm/cE7tJ4o/yr3WJKdOxkVdr4zIaP
gmW0foZv9T6GFLa7oD+8K3BbKS7PAzuZI/ddC2M3o/5ixxlfjb8d4wI1QY4At+cf
/qCjlFZDQvY+9VcfUx7q+OrOh2kXB9oZ7qK4Y8M88MhurJ9CwNxU05NjxK632Zng
1u6DKv9OtBsQJznIn4N94fo3Z8M+SnADNTEP3JTI7wkX2Y6KyujE1FPkY8MfVbBU
arQZMJJAa44Ld5V6eABD17otle6iBIbNHj6/c6234SD0P9rExDgtODzESJZquwfV
7nQhErihTpTavkK+dQ7SQyvs+zF+foy8V2eowSbxxlSw/FgSEWoI5pvVEr2valIh
CKKR+CRpmIWBlqajsx7JfB8+SNUVGz4DNZ2FrV+ADnxc6hAE8YMQlA9wmdeDe9Xa
q0YxSMXJ1oNitPzpyHZQEu+mSbg0/vATnoW0ZvOYFDlsTylbBGGX9cfj4hSF1Myi
x5Gn9nTNnKKRxXnYw4WOucgf8YP8rAnrvRw/e3375XwxWJ+MK/5bisjVI3x+ZZpI
ynOXNv1SEZ+iuPOAZ+OwPqQebsj0jbfI01wRzxk6m25VYs1I7Z8EEJUGP1xm8skM
5cgOJE1CJkA4KfzPTtULZGUowlF7W58qovuMUAKUzU4EVCjtpb3p2T5n6n0Kl4Z4
mHMhMwlldVGloozM8ky8frPnuAMP8+rSyQY+LrFEfQIoN+tqWTcffmHDJxNkqCio
PLGWENZBxVa4puzdos39TDD31HYz93Emw82rUlnvex5PLdav7vrNTCesOqiAmXam
xyR9LNHWsg4H3CtJV74fvuLevrKCp3BDbIHzLx7krj8ZR0slHA7JuzLdvUr2215S
7lsqpzRhakl2M0sRd0C1j6AGA8FrQyQjsl05dE5SlW4pdE5bv+J6IocIfqySjP3T
xIKBb63zv65eIyl8D9HW64MKYPakwgIo/+WeN+YdS8WpVVnWwxyW2fVYrZ2QtPYU
USRZ0TE7V0nIYEiG1CY9E6uykaGq5pUr2SjmU351lWzV9T6HJwdByq/GMljBxWA9
XxewAV1dqy+10/bBvRe+8SXX4Mf+eaSQ6JZ0tQoPE8gcStgBJWQvOChg6NuS+SQv
ViPa5BD3T9Ttx76enQaKxyKh/PJDylci4A2esGcJ+L+VWFPCO5mPeyVajQcxLeOv
vFdMRIpObrqA33dK/3tdW2gbU720JFfk8i69BC22PXrvBwglZEK32WBpofhdQvS0
kXkSF2Rc+q81eEPa1KHWeyZDyYTmHOPsI58utRmm95hxQjEu7TiZvlLy1VJwo+Rh
K6tfpVeUhPOpflUezx9iQQRp9vDWjfJt49/Al14mED+Tdj7+Jxk4ZMik55LKqKhU
uG91DxquloR5oxRexacZmjKOmFMDx92nA4FUnaXOcdXaoBBMUzLhRm9YwZM7NU2x
3w5GLWLIfFlyKYQlT9wwpqrRB0cUGZM+mTJEfz68RStFSmaIxgW8sLj1GlBSOGFo
OVw5HHTcyRD2x0C94Va2RhY3vY5gAJWX8ynILrVU4zqXOGvWC2702z+wtve9jLPD
upAIxL00FwuoVtY34Hge1IjjPOHanHF8FjUC2ywleG8Be6QA5W+9AV0vM3Adsh8T
Wl4LpYDF+ccS1Z5ADG/Gl7A2TGUOZEb9S0EOWnjwtvf9R7omNFWXRmxIOWQzMO89
yWI2SHMC1h7Ry+beRDHwZ6IfiG4Ke1zvwGmFJQLaPqQC/Em+F4guW67tWlfVNcNU
cF7KCOKMygZzDZjq0n6ftxLurWkAshKlgB40A9FTucoGtqnpY2cfcxeGx3bIUVuD
IUaAr1PDmifbU6prOyC1Bf6IN+xXZ7rgD2zzqM7aWYtzcXfQQ+kC7Ye7E0rWdHWk
pjId8akXYvpMXL/yjFyRjkklVJ0/sjbbgAjfuevE58/CV4i6LxUV6qGr/gFFPvec
bODbej/xfvvS5dVk5gXbfi9/hIoKbxCFVzQRMTQyaxhUsQLbMek2dC8a5N7IiWqv
DAbRpwnY8v3p0d1chWkWo4lEN96+pjF5bjSxzKwS2sl+feqs97dLO349EnY++9aO
JOp0Mehu0xSl+zFiCqK+Amd7vw1jEhkGKRymVST/VhEBNrZZExpnZG5DOiyL+n9a
97j1ZUW6PDR+EohZ1w/X1M/xejqGTYfUoYJLwfZfgxIZewfLy/N8BRy7ZM3fpagW
cXSrO/cMcr+jQiSrm2mYNDI7rlKKuyTzZN+kNX8C5jrXkjKX93VYsGUsRV+ncUhr
xBWxY6Dl9ywqpIfGQuFpKC8CsxX7jbC5Po8oVP15iAvhlCLPzmYKDDb7mC5OE4tf
Grh5nToYP3Cv6yjsvNffD/1erTqV/upwyH42cs592RWn4rbjysqgWtL5MkaEPGDH
kJMTh0ms0yMzsxVfGY2Y1TOel5SK+NDKvsUh+q8N09keJyCXbHdP3aarVWGb1klS
02zzx77jeR1dXxmChzBbscIVvsctrHBRo0MqcxE9cOk2q/pq62TaZ8nx3qN/8Igh
Bf5scTHAiH3OwPgSsF7JnOHbeGJFi7Xwv2nQz5zJBApmk0uXVc46VD2l+WJtn8tF
DL/sKtIZna/z1xo04W8CTGHdKxpoVnV9JhnkddSJMxkyfAK8ZfcI85aY40iX+xRn
jzWTrUe1ZKVT1CAfdOHOhLMYVaGJSY1obUeY9mJV02udrwCAUmbYSIon5ZbNYj9e
9Awf0mnkwK1LM2RV7VPiv36191sb3DNRztvDRFQj5w6Po5YfjQTHN+FAaJy/XHO0
qDjAZPZyzkhUX/TgcTgvCpprZbPf6B8eTRjDrxEaJgJHrrc4tT+MJWPoorgBPJIU
FlBSfYgX6fod26HlRY43mY8puhmwNbZ2eQgkbH+GiAw6aKaH9w+e9WSuyPKI7bGl
JZMsX07Rj4WwdOGqzZA3TjbBOlS+OK9mzDkyx9rXS830T6qSBDvXpG5RoMHJtKh9
rTZWNrvBWP4pHGEpsscBd+lDnCyjZmhxPpDCB2DOYDXIYbJKKA7XZrQ8u4At75Cs
+quC1Gee542mJ4q3l/zkGqXGsCvSUl9aPgUTnelsTVfUJqCiLpHUPd1k2Mg2VbJj
SXyZVWm+BiUBWj+RLC1S1m9wz8UxwhoZzL1CYs3PMdcWFiwXYe9TEVwo1qU90knS
X4RzdsEVgMuDAuH2rCVw6tQHblGn8q5JCRG169BXjvG5I6BzbZhzGoWwI8TGe8H4
e+1fiIg+YD1l3G0FpR76UobreHg45frTbeGtc3xHrCRLXzCmQFHxcoUoVPcQiapS
WAEoGU8Dq0sxfhCYNWGaWOYBVwukS7e2BpPB9Wks7B9nAvNLxo2a14WOjj9rD6p4
V8mkrqNhpP7tPkEVnhxEG8JEC1+pNUFVQxqiYpuJ8J7xJCdIe6wKfhNHnmzQ9RCi
JljttMV/IK01LPtmDdkvxxxMOzwIYMbUD1x0sou8DX/vnPtHPXpQt9emsPNFKqSO
dcMIvge1vpSnSAP7i0XbquFi2c3tXF2nWcSOO8oWqei17x9oqyXJDndv8aV+dJyn
xyt/qk0SrlOgzDSWzz6TMLqKIJROIHGFp5R2xjoabS2ZXnlF6MpwLt8Yu36HxmUT
zY+bSbgO5FSqsEoQH5/1TptNVvQ2Vu0Kynbs7OcMKViMS/M4VycIqi2iRgrbK1bq
PZg9J5FsdyK25QtQzbyQCMT3KL+GUSjStqNXgyjKRti/8d8009nr+XD9nccSv3S6
5uP0MdyutEGsMocY5w84fz5M3KbTDO+TUCDLBWQFnZLXDTQkAo3RrqVK2Ti9Guiv
9eShtNM357xjEOPVmoxXO1i4O/GxjvCCQpAjP7WYu2Zg8QdeFylaunUCVNo40DVl
nuXEQMyn7oDTHxSS5AwDqMnw8oRcJbuVuzNvQsZUW8n4kxUeRsSYqohgw2dLtUtt
vXyE/FS9PIFxO96ePBILEEaR/4aS84ZV8n2FWaQvx8B+jg0Ve2ixXWElQZidWPJq
mAmgW4ohKGEnn3NUDQI+GhFnasi4ThxHA7EQm2SjLkt6JABdQoVIxlLtVqLyL5ad
9uM7bN7wBIyRSYUfOIO34PsEtz9pJUKKuOAR0TfKOK3eKQbt9MIcFTASy2FLX1fL
TParvur+N0PrHOJW0w+iTL+euSCn976is1JzSVCG8MDgrtGZ1ZPB+e3ZBYCvAU3h
GfMdQxnB0tgFYrJsL+akKhKzpiXwbfekSKztMlgaakeLOc8/dKcXwVHg47L8NFAN
tUjAchjAWA9VGnAnOHx5vHoAsUwP+jImrnHXsb90vVbM0tNlkCeEqIN+/7yi5iMw
iG1ZIooPylwOre+mNZO9QwRuPYlu6KS8epeUKIQbzun3WExJEJtCWvpOjABnKj1f
J3JLSAaKh6W5PzQp1koe0kexOfMwzpBl7ueSxZCWBRSn1K3bjh+xagETwJb/k/bT
R0lCBUXaZHKZttAgXb6sI6Wgc3TgdcfpxnqraM1dYb7/hOq/JR8zNzc0xLmhO95m
RVGkbEw5wynTaEOUBqDEXKL2m1XTutrzukRpyyGT+9iWx0ZCttpH+sFEuqYhcLLX
rwwpWWoRsfN/IwGYFP6P6rgx7IZ0bdCGSFpRlKvvoAi+0PGwZJhzc8t+dBz2K9DL
KcDdsLmiESbFCtmRmY+yAC76JAmuA/9oVGjOoauWg6UrwC8fmd/GxX9ID3nufF4A
cTg1wMZERpGYVc6I0N8xJMjmgA62CoZPeEywz/w4OXmAkhoM8H6kp16M8QMsqYUC
aRZY5sjGsmY5WNS34Ww+ErZB7yKfzpqsVRRk2LzdmuimAWdzlNTzBluQYDNC5/qH
EMOoNIl106bVvFpKunCv743HIavSKW8y6UXPAykFzBSFVaw4AvEskDF8H+5QYWu9
SXupnm07gGZ/jnmc5sy0ZiYMLag9TGKix+YfezUBUJMEgnyQ7KeYKrdPu8VA6VrW
+2q6LWxTHVq9Uvl2P2t4lTSEFIwGiwXIjiVww39XVj48K0uwRoo8D7MMtcpRXoQX
oVrEXRz1pcEiMUKgM0AxJqXHRTAAmnzJYwYC/eJZdA05lkLXYOsRNUSMKIiAkH0G
BNGiCh+QQP8wp6fKF1sPvy8ptlfsP8FjfnQ6D6uSGsKuGAPPOZ0BXTXBGf43J1X1
neuixS8Nj+DI2pyJwztWcw6UVQxhbdy3w6TArxJSPle2QMigWFZ5QV616SZfeyI1
gMiE+Orgcn0ZJ5H7WBEDXz6y9ZDeK8Cwi9gnXIbY4IGkShaC8wxcpxBTe6HN4Q52
38erb/oeO0mev2eWW+1PbNclvXukNbDVV4HdHgzUvBQTUyQzftMYVb6EbnO3wRro
EHi0tHdYSA8W3N3YroDaDsfmlGkb1C0R/mlydg+0XFPS4VRCx2Ong8lOilJIrAUg
9Aw8GKS9a7r5lNjTkAr73VeRAWVF5eqsn4BoWnIECPitajvRYvdBI6+wgziAVsNv
9D7ttrphqvRA3BsAxYOehNwmybIMSl2PcL2AV9N4J0ALPNBhdQMGax4Ihq9ChC/j
Yw89dD4brfkRNBNtBJ5fMcolyDO0JY00KtjGDu/4pCFb9uMmzsLoXQiyqyM7E7OR
j07GaDY7BoNAXFND5XLrMgInMYi9SeX2a3o5JUKmCGZmHY5zG7m6yFZ54iAf5mYa
QCNzaon+ZgewSu7rFFMPlHt/+zMdp6ycSXZCKUiEAmAv+MNoavXExN4I82IBNGuY
4FtJ4m0ceS6T3XSM9FruxYRDdk/AR8K0aAfKX6PRs76wau9T/gl92ngT9d+N9y03
+86HpQqmHxuUtxpi5krPkG6oKcomuudROKlyIw63CyU7cjJV37Hey47XoWxZxoSR
q3KVYJiyNuFrMT9isN9llAH+WSfbSDncf+HjZyDtKbRWgAk72F++WdGTtagvM18N
WfiPfGC204pQRZz/GnmudR8ok2ZmqmX/Mf+T5HOrCyHdXDQvTSoc5Dqw7gHzfmjR
4qdYHivh6upTSIUJs7o9LvwHBs5sNy8l2ysocImBkIN6NzVAEvs+yYczyWDNMBVx
Tljllb+vYLsG0l6X5ACMCwRarB8g3jmlJYph4/kp9a8Vo/a8rGydo9jxNCSlyQJQ
At7bgRcDR4jEy8FuBoGr1YUD5MAepz6Ohs4O161ddY1K3OgwXzaVnx3bFoTy1dN2
k5mF5b3xB1VdgzWzl/e8Pqgi14bX1Yi/dehQVIuKc0+Yi8nDPFf5pEuRjZcgm/K5
PN7criS30MeSKKNxqTKsgVev/4EKFWFS99WZxF4be+ANcQum+XZoTW5RZRnz9xuk
bVWfunKtB7x+1eu30X4t2kvfI17IdWIcMuMhmeEFD2PYfiNAjC+cXMuaJyi1apPc
N6c5Dw2RWNSaKDr7kYYgUDz+WpZyUvMFRRGV2aOT+WR2nvFXiluPaQLrIrDogx1U
oEQRcfmtfe1XWc0s2Uu6fXfv+yZtRW4OdKJk8IxjAcDtvRjtby/nc3JilTCg2M1W
DuXkDFcVVlwNkPwj11/HI5TFnJL6OE8tnvrLKkfBVZ4rHM45PAEBUfgkbUM2EZae
fwlHYnBY3Ub0Lq3LSxVcJ4rJ2eFm7S4S6HK7u1I9QdwAZa3Ym0fbi0528cz8M2GW
9TZagBYRP3XlGRQ4jw+aiKNrstsoDS7WefPuA71eWNJ+URd4h/MCz5UHRW3PPLkk
B9sSwHBwB3NGWdgZwPhDwLtvMREYIRw0UoM7N519BwWSl/Li8ZSlZrCwmbGMxxKD
NAIVuFrdPA1EX8RirPxdwFFmvVTsa47Xn9TzRZKWvrk9iQQXei+HZsLRqMI5PIRj
Ad0F9kfNPOEr7NAi0POJf/ffEkKmRdLM80ykkQ3YLxm+uYMhuHryjV6ihAEoOsWQ
6TrqUDxksbbUYJOgi5ODlEoj9s7FnILR34ntkDNUAplLofCGVknphrg4jNolzC9O
Hn7frUZ1pfnYM88K0ADIMxvNISOSyaQP1ErGtatL3icnw1TYZTe1rOEeoNWNax/i
hv9KTAnFNJ7UcMgHAoF+ltvqjrTijFo72mUeTLsVR4SuQQJmzPASkkmpZF84nNOc
Oev9w0zYRPHvuudBNiQclC122MghWxQbYtnGDg4JC1dpyCcQL0585i8v7O7exTtt
mrT2dBWKAMnqFtZpoMHyNWmf3yskf8QLAnn3OLJvCCn8ZWm9C5g05UV7LpGbZntd
sq+C2Y8M2z7AswUuOTyP5MRrFM9iGZ08RT8gcrH8Xh2Tg7gQRbgY02LkTlZuZFdS
S0P7Twizc50NJ4Uv3wk4M2ZOUPfgyUD1cgKki3VuAbS07i6ZEqcWnr+lpkcYK9V0
mrFh5CDAlQCQZUOfR4p4aVqSWtIHBov1LU6eK7wBGrzTb7SkzNro0D86zKzhzRUC
zi6k9GODzAKI/j/WgIaiVSYe9mfcQXZX9aw2kSHh852ixMuFVx1XpUg+DYLPtbqb
nAHPUpoG3p5R/X39mGiITJIDUzx9St/nbT/2pdP5oi9m4tH5GUg/YrEyl/6+DewM
dvkQVEo0kI1BM3Cn1FZSWXeeOCJ7GeeCNdEAmnc7vV4RSFcVMUCaDzkQiVjz+B7B
009UbhfXWd3pP1YT3AiccvNHclfXo/e2unptUEdh2YJA4d83i8UQfHoxbytT0uUq
l/aQiNeo9qNRSOReNaG8n1aiFWY0DYrY/G4Gg3yspDrLsDMWy1JAH7C1sKpbcKq7
ELONLN27Q3VWFxmDvI4pgrv2vXHyn7v76fGTjSOxNKvjYYHYRdHicDf5dVx7Amqc
UuOm6kwpp5JTbrRIgDzfFgL2urPchTTHbM3y2+P3eE/SCrsss5bRsROBb/JcZL5x
vs5B5VClUV35/jjsJsowUBO8lmTi6BzTbgvnDiM1GH5F6hF78Q6Fn64WbtpFmBrM
WRMEH8kDGVCbNiJkWt2cUog43/njmNfh4lOhC5T/dLCa6NMIl0tK5TmkOAmnRORS
ftGhq+AEGBf0nDfpoq16tBv9lcqqQWKa4MIFrbIiixZHIoxIm2LfDcZVflK7rLkv
C5wbW4F0H1x+lJ4pCIxA2Bzl31pI+vrf463kRMQZYSXzKi5c4vx2bj8L41+KVTPO
zNOzLvd3t8qdT0KY8xFjRfBMsBhPUwcjwJpXoSpt+MiyP525hpbvmZxc0ihrxZSV
xmkCnf264cH2XHJLRR7DLy74WBATWLfU27x7YLNKg17bKgK0J2NY/5VMEPS51XQZ
wb9QL2QPZeRtbHGnMrU/P/HCZ3NIgl2YZCShrEBfgKjGFqQvJkZMk4yJJhgzSkAB
MbTr0q+I1MH7zT6zUuXuT/v1gcPGxI+JJIADqOPTtZJQkdhB8mFXmTVPu5TbNqw0
zBuyr8ulbg0mEhF+n6ofh0I3Rfcwc4YF+2yosv860/BJ8Podkr4EpSNb34NFGUXh
qPan4QujfarX5iR53AgGyOas0QDBjptu43JUOxLIcFwmwuy5dlsfDrg3abTRV7pb
x+lKxGmMFhtvGaY4ID3awwTbjUG2DLjrfU9zjbKHc0vhOdPKqxjnI/VTGc6wn5jp
1XvHlX4RFK2qhWiSV/5LonRJWRAelFH/0GC1nNMLpgvs2DbnFJWDQPm0TJS4O6FZ
R+d/2BJIb1umqxlw37TamGYtu+vMVB1Si2VlXktEWCsPRb+SMXGFW+Xsxh1YzjXH
AzF8OGw+t+iCkviJ0s5m7gf4HEwqCrEHT07XHbXvOapxVmptxX+5BKd0a0OExy61
f/6c0INOxg5NgjjBbwWwFXFtf80hdSkdfVJPlZf3lWG0ZHEXJnwOyjH8zIbNoy8w
VHoVvmRFHIu3JX5ZrHQGbzrOMnNyv6KzOitVXHpOzLYCKZ9D1+giQMEGNU3zopIL
XOY89SEACymuBLVIc7X59xb0UMyKQ/vmstMXSWM0RTr+jFK9oIySXaMxi82j0KP3
UiXJWuyFCWIKoEBihCBB3FYNG463MTDLEcc+dyxrDHaP5RRopG79PYMJD6mzrDcI
69kkx+zdO1jkNsOJlNSNaM/b/YGU6w+S27t9Ft6UsoaPNelyvg2ujwDKve8Fcd+S
4uXbOyDZi1qav5QCG1N4+N6LeecwrKY+TtJD7XR6u1yFwbS+AJSP5o6Pql0kG286
Qpx0go+LEhoHHVjOQJH7++HrFhoAamLFXeNZzj3BA9fGxJNudcYpw6YNbhMu5fsr
yw0lcQ1DsQfflPoS1qXqquMe0rI5ngNcsgLECNFk6YcJMPUBRYZqKAh1bJzOSLDa
uqp4mAiC1Q8SeGajK5dVoK1AWHVYS7h2NJMJOzwhkAkUlzcD4jA6YAr4GEOn3nPW
j2jGHU/h/5EA7fF5L2diN9zfBtoJ6kOESESvcdH1rcFle7jm7YbJ5gSSK1T+7iG7
fe7jIcYzXeQBOwkNEmo3z8luxfYF3+0biqFtisJVSBOuWbu92kRlX6b4Kx2OXR3B
MXLp8bvBu6juNLAzDWYfvje6oNSbROThppJxEaMBE7LTzUUp+OxotU6JHFVG2gkw
8GiuDdWib98NF8+/hepRVAAszloW7XwnxJ6NOFjrBPs/4UXuI69xebchUNBEpuSY
vLERlUQcTKcEsjz+fJ6yHSTOCw8vgmK5zehN2K4Et0+O4+G2BFcwJKuVoIfGHWFm
d3T2ZsiI4U/KPqdcK2jHmXZrYsxhpV717dfc5JXv4eO6nQ2jGce9CkFRE6C36cfH
pU6lYUwz7hUFUp4G+H8OxlTd3ulrItrlgyZ/YLGt1G4ZH46YUDn5wZ/+INaPEEx2
UaylvCNiQX5yiCB8QcDX6Jv6iOh6fbfbO/ItlGoIQLt12E7FXMP7gKFy/ank5OT/
cHU4IsEE1AgUYb6JlEAwS1eIImbdENYdniXRo3epddIx1sDHc1GLCwgEkWbPh4zD
GAKG3Ps80HPitTrUduqVTnwlFNjJ2+NereAFuzVrapPVf8hsghBNRlkIz5ybnHi9
0eNAGVE5sSUiEWnKQoNcuWrgP8g56YHrHehDG7+4L2noV59dV9w+8r5zDsEFzJgl
3iSm0ciVEiEWrgNbgcijgbfAJgfCUwZgwnpcY0J3tgKUEixee2I+Xy8qA9iUxM7i
nQ4BfbFlqudozO9400y5SxGDWEYL7IS+gVsQDNcuQCa5/n4IrtcgbsFMndswmGxQ
QJxP7NEHSfp/MJtouMMYQ9EJxW8/ulyx4OwIFHjwDwSFQdybLuEokuTMuIJIn5BC
oO91ezgrpKIUZL8yBRYmky1pcdtttow6l4w6r3AQK//SFX3lSnRG1+SemoI8DqC/
orUScoL6mrMuy4Z7svKVVd/18DX8lNW1rAxhRJMIA8HpGOtntlE4a8nFOiYPe945
bhccRWFLjVVlnepbVuolAslz4iQNTAWS+J2Km2bYjxnRcnyRHEzD4itnizDdXSLE
cOA5NvkYLLab/nl7oC96RAX3ea+jt1YbS5AAot3obvpe9iKoXZ3mpDVe/Fd/b+wH
gsOctGOBquob3iia8pH+jStIFupuoFPoUzAnlfJQx+2righuXxJODzGSlTR06cef
Rmhw/7DlWSVVx0UySTmBWGYS3m6OAOP+siio3mAPjX0oiHcVtf/l2nR7MptYx6X6
95RGtEvEWdcMglS/66SCBYRLl995zBsEozq+rGJX+puM7aPtRJcOkOKIbMh6pTnp
Y4mPw7rzjrtCnJtSgO9KiqoJ6SZDW71kzBKhSl+oXOtvRql1FYrUJYkVKvDwfoaG
EsXvv3y/TpbvM2jpAnoXsP/82AKbdmcR3iish3JSREGWOHyrq2nCI32uoFSU4rFm
yMZnseuCZaf/0BIDM3m6Lk/Z18mlBbykZ1fCsiw2hJJRyKIi2/SixFQqtt1+xGSF
UkHkACcebrXEfnKSmIufjkJk0lfnKVYHMNUdVeAZ9hOktvNUPAHztsY6Tl51HfC0
lvn3bfp1vmq2Wc0WchUAHNAnmmq38kLSYsa0VNQcxUwhAISpoT10r9MQJ4tan2rk
uaGwa5NOqmzhorCN65qjOA52PiqdelIOZWuynfdNwx5qwLVbNSiq20eRIs0/7sL0
d7O4SoA5EotvBkMUbv9caj1XPNs3zt9hWNMfK2rL8mRuokKEob7b9JfDhpf4LcHN
b1nzrkcS6evUoSFHB2RNZFazKyiebMtOvbVJddoyPlxZKCGI+pJj+XXWaQxuvfxa
qliDjb9Rg+LuzjqxChirP0zHmT9zfDQMIoEeay+iFHqwzjTeoJNH5D9dBp4gFV34
qwlqO/FOg9QxO5ZiDgSA00pFMQdw9WUleaTsQUMkFo3nNpBQguyVPqvl+yLxp1ra
2svJaU/Ghuvv9+8xnKWX35bbVpdniS4c2y3ZbiKogKDkZttGVb7lgTqllp2PqQOZ
6nZkuT/cqFD9mU21Nii3J7WFj6gsArntijtw9iDCIsTVUDZobqlZ5aN3ydQDCA78
Lo2ZlcrJWsD7fo4qejVv41sEH+s+DXfEtcK/7lNolGyChfELo2aVFG9pvrA0/9k3
b0zwQI2m2CE1xdDJQvXg4ruijR4uEIn0AwjDXRZghgY7JQTNAP7Z0kJt69iExgBX
W66IOpS3OOTP4fgpLNliSshNAZV3hecwMHw5HeaDZSbLIFhJUdCIKbbDCdr0jsUu
idJwtfB/nh+lW5OR6eU4JOIfd/txY4IZ15GhDB9hKEFWtP1pxmj1ownoIt50tRMB
/AebZccAvS6uFkLU5R/qfyQh19PcJVA0ZIKiwCB0gTkix5bdaSPIlpXvtGvN2yrj
LZCiK01ULgCBv6wMXJgNmyEeDbn17Zlb9o15gJvF4MEfJDI41yvQNOPvoqUcYR4y
ba1YGze3NXZofA4VNu6YTjOeNzWomrlkR38IfQZiroU+ldJjus9oermHCM4aExfR
mR9F9oSgXJX9rcoa5YSswsj2qZf3ViKeNinMvjsWDFuAFnxAHv2GQI3MmxPssEyp
uTkXTgBqMa/EBPPB+865p/BUg1sosHRUu9xo0eTZdsNAM2ptiznBHQGL3fCL4eX+
Pk857eaEejRXQmgG07xcKEKvrl1qeRXAT01Bko+kGOavkfBda9/lHPkkZnfDYZLM
fHYGZRmQjsuN3wJUW5vLELU9DANeA1hVfasXZC5MswGoR+ikYiT5UcWOTUvzyMUi
1m5iNR6bL8Q0b12Z3IOLpd4zQWKDjFk6UlI857cDJ9tfoZG+M6OZMAXAZ5pxFOV6
4gxNbyec9YjvATLGv+sQLl3x0XzKoF2k0uMJ16450K7Kk5vHhwGrp0w09ei50F3H
nZXwueyTYEufLuHrPRrNFdQbF1yvoot5upqBMgr4K/Qn+SMbtVN8y+wXkrc5d1Jh
Ns1FW+pI8g1wme/V6pAKPrp0Hz9qI7+Sys5u3c3LN4qWHTSkbpS8KDr+Nldsee33
8ckGwxWOfk72KVWKt9e3XBBYZD9m+KS4DP76P7Bxb5Eh9ka2LLIJM7T2yxAIsF/Y
6oeYbkmKO4Y5sXEurbT5fjkb/DKfpcWw2WsL0j00oiOe4V4UYrrzhZl12/QUNtHM
t5JMh7M5YUoCitnoQ9Ew3vS0Yo0Of4tYPllAi5adIWRL51JIDOUwwj2Sxa3AGl9t
CW0hHBEUNrGiT/ZYFhwm3iiT2L09vUGkVyzgqVO8Ee4fP6dmzYFYky7LngCfB0ob
DOAyrV2ny6b2fjxktclD/BJcUQf4LWosTDWtGlwHXONKKUnzExICZzOaUc6FJqGa
aAq9t7eny0PGI6q9y9rd80k1tcKux8746+NvklPKPYHQbgEhYHpwDeVMBcYR4Lju
wo7goRRQ3WzG7YFvFVChOjcM5gyaoDh5qyaP8nxAjuAZt9yDmmpFNHvqjT5lM7jn
fc59Sh3zSpj9dl4FMjDwa3AaNXMwEiQTb8D8hU7InsTR2fM8mcCo7YJuqArLZxCX
IbcoErzex7jBoq4dlDgPPSOki2+2tCEJUlfoL+L3W2PkGtjCV1hcBwJ3HA1pkDuH
PT3O225wtxiDJuBuEQtZ6f409nol5RRJYR+ViRC5JTicFDPbKyW6g0/oQ7W6IiZt
M5jmdwDAJt5/iLA/lvFZ8nY2eDvGThZ8XZRYXkogSOjkvBJqO6X+aPLvhaKocIRQ
5/vzrnchfgHQQ3tQNYkLKhFCf2SFNeOQmTZRKnI643FbncTk/WClV3UYypl8l5QY
MNoej0DMy/nUVnL1+UB/7WnI3GJv63QXyhWBe1J+LBOb5+sLfoQZIDr1nWVKVaw9
8N/V7PZ32P/fqpK5DGFUBKRYtliWvzmfB+oc3HSEdpejeGCEYO0/dutPD56dniwc
C01AvEboXKRON7mMg2ljxWwtY0iupYUIfgr5+0TxnE8BsmNuI8SWX0heWigFbBhS
XU1RQrhtA+VhTkqdVIZ1Dnyu/rglPebNeGQVhwt89YYql2o+15mtsUShny728jOo
3ZNB3IBzGPRe/CAJpNDbf/Qy8p7Z9BodbPBcUAJXHm4d8Jr583Wp59bSSlcrSDbi
XQCg24oz1YxZ4IOJBEIQ3bimF3DzFpxKtfD6JCiv/18ufj7PreuNmREbzQhFnpxR
2BvZoyVSlVPAvB3PPM78jmfTq866PD49209XxljdiDGrgW5XQ49gQv82+UqJGDIC
MXeX5/hEPLxkNcNeymt8EP2Q5NrVpDY/129o47KC6tDy5askU0D+/hrRcOzXiE0O
tpi5Crb4njyVcGNBjC8tYJ28AkAuB7cyKbggsm1dCEO42J3epCRceYC52cfyjbtX
jFe6WyiXYR4/GHVgLfUYLeVtKe8scp3hRajcZPHVs+WbAG8jASFQy7I9ZFTuNPIP
uYvBC04b81e37ymcH/HsIdYqmnkW8LJg2+d6ZOvl9bo0U6UIAiruOrTRuqC5st0k
xszKS/mMKcWFSyIobDo/fIM8iZ0MEZVM5sEBXPebDsb7EQGoKdiGiw7HnWcJGW11
zmNrcWVEnTVNb6Ao0Y0nT5Sg+BNQG5aEmHQoZRMGUMey85kNRRUGfaXAFGxZsuFE
a+4Mmcxuxtj+ELVvoDlB8isFUo2fTaxYrGK5INuM3PAyecfm7r2jzVVba+CpQq5o
P3zv3EnSu6Nf3I6RXKo7awfFyrx+mFmWOfmOlvsYikMa9O1vttVkBhpRaQmwSiUF
S2SYV73dFBoValGKeSC7g7PcF+NvzOHsKFMx8eydbwGKmFssKKIvGqOeNGr7iL5L
m7qDfy7tcnQ53yFHPDlXEH8R63KdSIfY1BoCT2KMiXRnXqBTO76LkJbE2q87a9li
wSP3McmPJVYT2jea6SrQFwtUYgSksPdG10EDWJvgAr13sGOeZ+WWDV15jnpongo4
GkUMm8sEDgYBUxWccc7JM+wf0+YqX+uLNGIQvDZoNhmrtbh8HAyCNEkRURxTk0t/
6jnt/HvbJxgjxOas4hRWQnsaHmxI1YfaeLI71R8dSTxKl+fi7sgLXS8vTGPsjDRU
OXPnd/95y4cAh0l8ihPO0KXXtuFIPTCL3B36wgZhGnCwVmzQl82Lj/l2Of6Lvq6e
DcaF5FLFFSfTrc1KSM+CBKKiY0+J7tSo7XI/j6MN6AZwTv4tg4MYvmB0Nj074GNS
tSqcpHM4RWWeZ4Obt4EwZJB8JpOXLd8/A5ejGZttQ+zu2fv0ORoPuAxWygbuBaXb
XJmg5b1cWQ+PgRnYA7XXsswQL0KMHuONYyR66DPe6Iwbg4V84pq859a3JOCFc3d/
FhyxvRd9C8m1wLjxp2/ZfnUr8hp5xTBoEFUh978LiR9kCIj0q8upiLZzZhNtarHL
N3cYfK4Se48CASioLWEra9qnKcpzt3SJIAS16xVj4X5JkrhuPYe5XJWL4NbRUuSa
cOlgw2i1HKcYoWDhnUqgkppXpc9hdPr4GZAfwhAbJtMWU/rDtApOy5NfgmtJI0q6
MBshs8ivIz0O+a0csnOMkdh0K//MlPuKmxOqS6Rt9pq5yOVDw5MAVUADLM/Bc26K
Fiss2LSPOQvXwMu0teWT0QEgKPyzwlAxvT9qTWRIxucqdqXIRtWSeecrMcWVyjLa
YUUAEB4fb4dxfsgX9WcFzFD00Q1Z91EpRXpsUGLhJrxD7x5Qo+hPpEb/c1CD1p3q
vLm5ERkSCKd/M8cnF87HBAQhQdeC38c1d+c5fNYOKUZSKw4NUkbpXvyTKxHubU7Z
nLKWBZ5vuCK1ebiul/rIdPVVtVgXN0w4By7fE5GM4KQSH6pV9r2AKzoGwweeMfRj
mo9DmKpS4wkiYfVm1xmsewI+8+VtW1UJRz7AXQwJcgERdaUhF+tky09Z7TqGS8M8
ybAf1To63wdKPBzN0Aid5A+GIcViUlUAJIM8oazfjbLCASkP+7diK+n8nz7IWmLf
xXaW0v/5cdaM+YtYyzPFzqqZ3ShBz9v8B7kbolSg/GFHZ1TCavKHipR28uW+Oo2e
NoPlLC1u+kGLIuJDXZaaZVU4y8NR+K9sgiSCCC0T5sB66iaF9jQdiFXhUvkCTSMg
0p5o7Ie2Ov+SiR9r+hAOpv3v6yRitnaaJllxghnxshnBQxIwh8QozSPPiN+t7/r4
Q+uk1rcJ5OAEx3QQH5sdlz75EgK0p3JRvwMMvlvo6QrwjhWsqS3NDmGsLi6PYFHI
QInKJf/VHW9jDJK+zLY+g3Psr1lmoZ064ADGDaxitcy2Tylx2mWsj0YvCHKYi3dy
zKe3+3hJMfPu4poDBegvEtHQnatRMVkpSSgjpKBNHXVt7lcmROTtVTF2Co89HZOJ
iDFJ1OHzOIJu5yqRRkdF/v8kmOZGjh9aEN3WDNxfkH4zXT8bE+p9BusAU+EjsWjS
o/MV7jyszBoksr/asLRaKjhfDog+PEveubgSsNpsyuu0lM+032VnoV3VjWwi4sml
FpYe7IrtLkoWCO3pkudwOb1Li2GtOeg/JYhFQeUei4nzU7xkdwdbjndUJVm6m1Ti
+sfgUQMdTqG9cMRYS4eKKgrY69z3xrMUe+t1Tylt9eUcWdk4WgqgEINLP26jFm/u
YSFThUQXHOGbAVKT5D2YUzrKfow8AjJsp7OMOrLEE3GnS5jmtj1qvaXjKoLPXZn8
4IfPdaGDBfVkMOwciJ11go/lbBQ3pPgEgNRgzd50Z0Uerj3c9tze0VjvUdJO55V4
oILebgXHaaXCtUmsQ8KtiOOABs9h85gqTAijFiYUtNKXNlTsuTbXsLXqVUu1mZgu
5cyFlMMXnu6NW8TUbfGT0jLb1K/gRXQNTy09zl8TvEyn7trg/jffUFCZsoGIgjhT
rEtRkq1GYW/unZoOLuuxo+ZMBvGPSB5HDLoGo/YXJ1XVtFWPLC9kLHY+YNxM/kSY
HX0XTx0UX7hdRSrM9qg1+QuNkdkZtDgvCKNUnxVxh9rhpSNwcdIgT+JKY0z3IC6H
iNp2GtsDU/tHvHWEBvZvTI04Qqi/MgSJ3L61Cep2qy5BGNpihQGaAzZ4rH1Mtbvw
gneNC46qGdoHo6zw1S2Cey6a7mv0fDNjDE9q5zzCG8IJ1TC6SX6AR4UwTcOgCdZe
A+3OWLyAeqr1N0PaN2Jtz2gsfM8o+ODhclWklfju83RU//4DgMDjMtpyrDGd+yNT
1/Cb1+lQo3iz72IfPl0JcD2UYnKBaCW8lP/bz7BqmEk69LmSnllP136mmtntVxuv
n9NAbh01c7L0nyj/EjHcVfsj0VCWqq7ISgM1MDeKjXV/WOTYYE+EVDb4j2Vj8JFZ
ZqKs+dRL+afeWRwj3tgqDQGUXCwEhbs23eHLZY3ChI7yIYg5zix/va1lKaRIfnJV
m1OOcFH5rhddUlJWOHU/8acd31WRwB2CaaBWK+Xrnwf82KTaJo4/oMg5EUT2MoPl
YDVLwunuLtsDc9yI3BT4im457rmnGnorSVg6pILHStRiva+IwCEKXYcE9uGmD2TP
Z0vU10wHAlSK5/uTwiwhT8IxTsiYafa9BEdhQOuwwJD4HiVDyahwhCgmSoTjN7k6
Itg3mBNF+hgN/LK53LoXc3Rmwuu+2cOxnxvgI8FKnkOvncACZHBsyrxISgEftVnF
hP+9IJIi3l6+devGwlLP6sBmDSUpkuqlVHt/yzOkGunSJcK89yfb5ogZj1839Q4Z
IxpSZ03SpuWAP8we6aUETyK7rWhCi2VO9W9TxcMzto9xkln8zr8pJoYWzx1sylI3
z6/HcWp4GD0406cSDxwkQ9kU3EYabkIbDk7AYpeX/6ep5aeuJBn43n0kl4Wjwr6X
iP3Y0BHsTQ9rhW+vVsgYhxB9nCM0su3EPTuy4tFzL0RImYyfyIYJkvL96c0IcYPC
iSvjT5s2ui35HZveOfhAtRaiXYd6U0F/XFQvW+1DekoDTq9PMlRSHDrwSmbdn6lS
zMVA0HLbSKqXeSBOwscuwpvAJQT2prXfVGJbcVHhLD9oJYucNgS+Bd6XQSjvqBnb
A2ZP0y2AZiife/qwMBKPE8ezLmmB9rHwEWRxrUAHFw2A1sVvL+ERs017pogrWr9q
HnSqU0YAo8mwiopZnUMcxhInDp+23nMJ/ODLl0pR7WCoqRRI4yFuAyImXBPcQidf
uIVfomhGbrdIMug70Fq56PEQFnyxYBqD2saayQTK62qO000EsARIMs9eoxczxAhF
64Iw/invm5ZMCpqT9caI/wJlO5L2YM0vCtD4FMVK/VdB9q4mMzafmih5WT9R32IO
LmfkZpNvqjnPPFTavaGbnGMNTcx/4dgaU/n4HDEEll3e0OW3RpiHDeehl3tPyiVx
ahyzLrYN7Hzg6F7HhuajH6vP86taAhtn9U9X8xuoVkNAm9E4E+/q/BPvU9Q1dAwK
t6k0KfkMEjDFEDVOZWWISwNlrzH/2SqSABQfG6AzqXBe4UaNbom15Q8YOdcmBsCp
8JbM699B5IBtyGR6Ywev3Sm7h+rGh5r0i/ZRv6UHnKhhT3AwGz3Lb0MXltzB9T0B
etHMRGIrUZYUS2u8QET/zjUd3jvu/cuiT/V8lbaPEQkZUWE9+WlBhXd1jJIfty0s
SVgP6VjkpFIeeXT5Zrr2fi/2x76zlPmBgwnK9sN1p0t3BpxR7sU1q3Qq2PR3rwbk
CQmHjcWjkFOOOfB70dtPhS9HBAuB59H9isdu+bnoDrrTAeySfY7F6bgEgET6uxSn
N/3ldhxIr/SoszlLBkI/Q+8wANrnBT3ta8C7KA8dafttkdI3P+wc7SR/WX+w44tb
ORHOlEBfwU/YLeXFo4mUP1S9H0OO67o6wLWYRxYUMwO1dt36um/kej98ftYMb1nY
Fvb3JFCzbTvSpz21ezPmZUnB+/tk18VKtjTsIQF8PurM004Bi50D0NW1jk88n3fF
NjAAXY3iX8gxwEqej+P/jE0FAdmyaQ6WB5M0eo3P5aFxmjEFPIIfi0f7XW2Y8vgh
Yl+Cj7zXmMkEfDTW6PPkAHlcuBO+KoPsSbiVuDRuXpQmunwkzG9M1jn4W9y/4koI
mRcLN/cn/UxVEuvELIxsTRSgsOZIUx2+0+95DqvGjITVhXYygAkiJrWJCtadFIr7
FmkbsDR1/EZ9cPaOyg5mT9QNJP6i9UTgBdbuH/WKl8PMXJWe7ekkg6u8yaITE0uR
cbRxNZR3cojjdaLZ9r9fL+uKWZRB64CBFJShnTLkvcbKjR+q3tQRKa9XPs+21+R1
uxe8yAFQCXlTPr+9AJ97ScXbHdqCjR6ydGqN2TQcHmrm9PUKtgth8quXZfRkIxDS
F3UNju117B0Ae0BOYWfnlBOQ4aBoTWnmJdV4U//lskP/Or0gafq5oXdb86DGD9Th
XIEBSNDQaKFxLzAQ05CxLduDB11e9wxZfXYH4R31BPoj9MVaWaCMS6u/ojqotNq+
fzB+1sZsaAQv7pdHaw5ThNHiwGkNRn4PtCoB+xSTnkcWg/Ho0fiJFT+ZBGHN0TRn
0/7D04jDo6cjpt+K4yQV/RhlKqSoWoB3hvZWNoHL5JJ+xBd+qaqlw5Adlbzs4cyO
UzN1hmGfrEPXabpqewUzr50eYpZso9Ma0xvOzh/mzNNKZ4I+eBfh4M5dFVbxcdhc
12wcCFogO3D2dHiRVzjiTn+e0JwaJIIdHLcqu8lkkvAQdEpTklmhwNbErcbDKyYB
AEm2MguGkp2SSKBl2G94rIIsyEe128FFaxwZQScgQ2HzX/j9aWAdzo8VEcN0P4UW
UMdz06ZfxUQUIJmt6Vw76X5XKEzmj/o1A0oZkKLd6zhCojiUcMpNqYgYBtI7N5av
rkI2xWRSWr5gCSLvFNL7Ffg6iZXTyIF7D0D6jHtarIfDy9ZZCx9zK0IOAjTAuTXN
eL8DMb5ksEEhHLTH4Hrrg3JrgUJUdOCT9fVTCP220KgWNG33zn0ZamzgNEddNedW
3Z5cKEc1Gnib3rPj4XQNii4IW5vGBm6aCYGXn7gtP2DYGPazptivstsPtrFfUps1
xz3zsJG9013d1DAu5hgKd9hVhRDV5vGlfFNa8op9OWR7ojrkC9nC2W9bDflpSIG2
Vf/YCsDO8llpENpNsgfuhnAFvj6uTeFoIeg86sEeJRW+CQM/OR+AiQvxXZNTb+JW
10+nFCYQi9HV8uc0TMf31VwoH4l5WhERZYBVFv8DitpQnxRJ4EZm4hJJeKz7I+Jy
RQYo444OsFtzH617f7PiYhrWiFmg6WN5NBKYN3MNkESfrGM5v7S2Zy3Ne6LMd8T+
Eij1W4WTAd+Ahf+LnHUAqE2NRz82j90HtDYjsjvXZbSAV0Bi4WsbwUaKeUNk4EHn
6n+eQHIQl2ShAdBOMYOce1j3KHgr3uFX0x+990cz9gKSuGiG98Vf3nB3+WX3aZ7s
uyefIBmIlhwuFdm6FzBoNTIK4DbOFB34VQmLU/X9yKptMr6BbTobT1V7uaZZk4pg
MtAA/BzHy3Pp0kaIRVixD6CAR/4lFE8XbhFnfn9U2X/BU9ZiY4kW51ad6Uodkxgm
Fd3KvJPFCoyX5L1eC4tn6qzY/pkFcqANU50krPFNO4TKbe4kTTBTZW2Mc1LoHlDd
LgX03+tx7+jXzqTd72XIZz48Dq9ysg8KsjQuuVenoigN2K5JUiv+z1xbBwv1ZZir
LUfgS6R3rBxXyCtUD2b7vS1W+u52KBCa1vWl6OgKsU+2E3SISpDGFaAv0N3MU+WY
PFgjM2DTL83P/40Q6Yj+YaeYhA9tW1Ugw4CqC+Dk2kjSr4+4VP2AZrxUUyWCIFxc
iMttYBRkmGRwb0OPQ7qEMko+YjpVDSHRWKIaHouaStDmKpearwe/M/bUe+mUjnOW
ljDIbqlcL/3mgE8cIZESwjxl3bKuMunt1GiHo9Ol1oM9iRHhGApku50G/PhI9G1D
lTmy8L4FJhFrogGoxR0mj7zSzfP4aKLi/xrGAy8cAMTRrwRhg6+7pWhc18CBMESR
aXJAiinzzMsA6MPduJ6301Vus5Goy0SfyFl79cveOCTAzhHuevY0DYbx5m8exKrC
I5iOLQ+JTjHPQ/CtRZuA/4sQqsutjVB4M+80T+WjMysKEUPK9t2YAHNMlNfnCg4Z
UxhYr6GD9XF8Lb+RXF3jPx+LR+D6B5uGqeUWeeQ2IUrN4sDA7G08M1XPbWKaK6Vm
crJ3t6GLLdYKQz/rYrQOMkzOoxF2u4d1vGdDVes+tbUd5o0sh+8CsYfpJkwilkku
gcFY9QR4rq/CJcNMq5ggy0s3XBiLWsH175MPRI3NWZMqV4e5ZL7cNLQfZie0uv3D
kWvpMBodmaSmmdScwP/L/X0Cc2IXjXEmI6BypMvv8adqTaVSPHce+1Ayd0vsPGpt
Jvs6OiboFTp66/tlX/HWqE9rAB179gNkFgXCBkTrkfixXc3OCmvqOnvsg0OAiq5T
26Z1kMQkTPP9JVvZXP/IzooZOpN2cjQ/OLcvPQ4mErcxO05Tfm73NV0Iz2uZyRsP
2sMMlfkVJV+G7WYXTz16kyVGauWV1gZeW8QD8tgMWE3XYoruiOUCF41E43gJ1dhc
Hnw2Tz9fD7Nvvr4k3nLYJKfHrup//oGQy5Z6M9+Usa8eOPQ11O36uk7V9Z3fr9J5
avNCkf4U83V1Z2vylmGjj2ayN0QyaLwEeqERC48qitF0x/ufiDYG/Ps6BjZzKm12
i9kBIXbIiKFkBMJ/dqJoNOLlokWipmOJwnxLv5SQ2xtHYFmmx3Us/qmqYrHFTC0N
KzlzjKfvads6ZMKkStrI6R1zQYpEuZ8HEvERMD17id6EGko9etl6Nyi6aTVcrWtU
Z1e6ZNc34Oo16tDbSAC41QUda98xEjehDJQh1eUrqI0QHntgF4idFddwuBOLdSdX
5ZDMw7kiz+++gFentOg7tVMmw/SwXsGolUEv7tW/aQSQE1Y/7Xqquz771HNQOzHY
0xwbs7Svuu1fPtKiF/P8Vr7wuEu/LfCGrI8C3hWiC0yOVNyvRlHrrnS1Jtkd1FbQ
VfLjazrmIXi9nM1CTDgRmcKbnPeokQALXCYkKzs01ZugCZNG8ATJeDIWfB5tJR4H
c2ru3DXk8br2F/r4rZ7Wtz286RPll6xIHp5Iqlqk2gj/fUiZXe6IFtkkTLei2dsH
vlglfZB1qz7fKvPe6TsQxyBaYEBY8K026Oj98prBIA15GOFDCuvk5VL1QqIUTKMa
jeeKNQ8ApbDz6pmk/yyMeAlR6HOGFPozWrJhu/YBi5JNGLaOXNE62GL98769dmRB
2ktKhgX4o/AIj10U3ZoEaH2a6kQX730ewtIg4eq5ogFkEYImxzAB+6DqjibiRPRK
MhxpkGx6n1gXcxWZI792O/eC2nblKhIMwLWdekuwds00v6Qc7dsZjBZBzoNHN+uV
Y747p3lIdK2Mk8JQpeNyH1S1RPrfBcIocgpT9bQFSqGgqUIDAyde4pJ7R0jnCqU1
SHs0Lft/xSMzJSCjnVhhdJSly98dqsJTDEg+heJQCFKgPWjy3zwXiueK6qBoEXLA
zkE5Y31f4JjZTPzgz/iNNSJVuLWNL+qGEP3/iDbAwNiBqJ0wYjfIoPLgV2vdS/rA
Pup9KutGSVgeI8+i55fSEun1/xoqbUq7Fp/LDF78QsjX0ILbgaZH0nutNo4tgaqb
WOw2TsZMvW/aJgNHM8P9rDYt5G6oW+GiyPUsvCtVbb23Qo1Btd+V+y2veqPD55bm
B2p4WmCzVX5Q3BNNcO8Nm0IGYoyc4lGG2yplXJcVr481ijaQOXtbVxUNO43QbNAw
slKZag7IiPt+db7AUy7czaQCLpLROagPzGTsNoL6sQzEODgHGWzLSfk5Oa20SYYR
IOjJAvYqx4JOFl/qrgUtkxFGSx01LDrbwnsNhimA3GBGCw0XH04xawqEzI+KcxAg
2jVZ7srswqIDUasOiYrAlTxNKKg0c3otU/1lP88BlGxJDOuHnV4e7NhUBxEMhaAb
vS3AevBbj3TO9HPKlxtciwEKt+cYyRs2bHnxPx6h5kZY2MFfc29/hOpRweD19H/H
kjKP+J9rYhsPTUrqGqME6hUcrS5Pr5UTMpS9wk8N9h0LYzRrK+5K6q2aBMKKT2tE
+l/o2A53/8sQTeT3RoRHIEWx/qVyXUooYkAfnlaw6a6SsYnhCE/fp0oHIJym+/Qx
BfWX0ChkvgJj5/lg+SOVc9J8fk+cz3XstjxxuUXWCb1BUC4036nIcyW/Opg8Eedj
O6FpvVRFHZPWo7dgp4IElznRMc+YujoX9xofjnNZb8f5vdntqDdEH28ZHCUyKWr1
YkymNe3qtIsYYQRiWQ12u7PfxmuhE9OV9LsbvnZaVxDKnrppVAIFpjxe8YtNiaix
PY/kFkYWhP++D/FcW3AWiztjpIR6K4fX7doBM874Cblw4C607mov7i58jtcKT6zK
FFFctmHgVyCSKxkDR7Gc5oNNNV7wTA+j0ZMQu90DZivzagRsjTtJBMVGBVBQPR3L
Ztkeae24Qy/jOWhnvWBIz96Yc8kzL8ZfH4m499JiaUwMm8kT+crNSDCer/L2TgwR
bHEFMTMLy5GLY4yhFaqJk+ZLjwPVy1Bw13AeBb49yZhXASKiP0IuTg+T2hkGeK1R
+EJTsbe9eYMNp7vZv9SPOafZCCLQe3b01pVvzNyLbOT4I5y/7mB6LGFVK4bfrf5U
33y52xPMY5J4uQUvVuRUzcPEW7F7lt5oWpdX7EuHr6WSTzfSw9twCrm1j+eUSjtM
71C0ie5EMSFQ9uaPW1Ty+UNs//MbLTbT2Q5kfJwJg4yyL0b4XdvdUp94CvjFdNjE
RJCt9A1U+FJFdCvdNxWY8r4Et0pdhZ/gARprtLzHQGgIRNIShqcYgd1phHg8DxAf
XGWPR6gd9f2nNip9yIBIn42B6uHywpKylbGlOOuQ1k/+6KsaEYc+tyTjysEexiNY
V/34Bbury9OIhDGFN1fNB5srf6PiOlDTzcAaENIHCqj/FPs5nAaehHEPHw0hsVT6
bncD5YrJNQ9ZwVN5oYPEAZNeZ+KONFjs913JrEs5erRNr5B4hKuZZOJSagDuaNi4
zhf4b5FjkLR/ow8J6wfHykaNGPqxrpRcsijk+64VzjzVCuJspRK5+6tofWsCV4IK
fMil6nBywV6bbEPxJOlJG9PR54ZDt1NwivdOLexCt7SmbN46+NOEJkJCTudittnb
YO79NbPsAeAxk29Y/tpd5DRlCn5e6sfHw/1QKC37v7Znyune9JuKvYAFCa4WKoUf
Z3veb3jI3oFv5Gq7+qQ11XuX8elue5csW+iwnbEeyjTz5DqukxgMuVeO8oqGFd/1
Jm6JzEZo5wWmnN3gxKRqx+3v6NOxoX6T72AId+FFADE+rytDl6FVaxl6prURq9iF
sKz3W2DwB9/uBsuzp4EqkEjjTJiZ/KX5SHuYGJdwmrAhhBZOQhSkqVTn3s1DWfRO
N+DqodMD3XqPGFMa7oeAKk6dxzoIOep5pwfXmRbxH1ItJmW9WUUFWZvI9tykEtuD
TzoTYVxBbjLXQlx5qdOe/0P1GiwES11p1Sl1qHctO8lXXFO5uHN05mKkNTjUJ205
8d8bXZXixhnDPf1swaDxBxhOPncUmvihcDx9U+7Wj12fLSdZ2ZQfmv54wOhKjpPF
4DCobOGZUXbzLrPfwmbFWR0BM9tfOyKIlzbnSpp1QjaYB+DDjBLIqoxGnYR+Tt4i
cq5wH0CQUPP3k0UBC/KpKIzvGpl4uY7sBpWNo9kQMGAOWcyGucy8bdPz1RbuRJFq
jDIYowE6+qEz10ZyTsXgi0t43omgYLjv+m3AdnMt6hhPFFIXjAczmvjAEErdASps
it9aOBitO+1MX7t6IAYCPA4s2V6PapSV+sxv/8lqHoArG9xWdFPhXcHTBX4FCOpA
9IiboW8mf0L5eEcHx9GL2bbUyILI1dWJiZ1UMmSCbhoSLgAMsDCAKR7XJOyUhV4R
qPlPB2PU8CJ4rz0UIjEpToNxYxE5hTVRQg6kFX19tTa1q6kR0kB1qJtIyojiqhqt
X/D78uzOvfaamMEAY8k+TdMUQ2yfbZSmVkH+Uq1Y9Qiv9pBrryDrBmuBFkyY1f04
ezxF6ontjqMTuKfOIsHorCgFIdPa/vCCHrUmQnFO3GNZz6gAwLu9S7fhnc3JU0tc
c9NVfWKMaWz6WbbPpLb0Y1U3k7ZMT+u4J+piuygvnc03drPfBUCN6OWPjttHAof3
Y0+0dWBTrbPoVSyVN91mYACbfuS1Mn42Ny5WsPdmQy9rteceziqNaOA+Qyl1ssIC
zydluv3dIiN80/lIU8BJ6wOnoW1/QPt9BbeVOA5/VnYMoibqWWtVk/L1bBL82gZ6
WFozcihZUBEI2osXIOk0AXeQx9KXf5viSGgoJMyKcQ/2LaHTzGr73WfgkZHWRmLL
Zp2HqJ9S42cmrML9Oja+2N04V3AaHXVvuc8UN/wUZ8y5qbZSM/i/x/aN34q1ALQV
qu55rVzaGCL0nsHpEmk2l+KnERIZgAVmzfekuF7/KfV+dWbuj/z2oAkErFg+VLd5
X6lYckhNwx/aO9r5q2g/VSZtSOyyLh1q3z98U0Gc38GuqUmauyuCfHRaK4cE9O0R
zRowiihnJ/fonk3lwKheXsZUVIW0lZc/nFq5l5h6uzzZuH9ze1YBlVwgjG5PXc3C
BRI5bMXaPjC1KVcyf0FqpyJnR9nf+2QQWo96R2o/FKmhvWFrLahwSAuhaqYgIGrE
Qn89tER1rPXv8S564zPQqwD1xjnEYMdIgGrTHy5Btp8aQ8i8DBspv3AoqSkib5kL
TGm1YH5mZNMW/pfAjn0GKITSUeHgmNU04u6XSFMMPx7yghSJibUH79qD7rv7UIQX
g0ESnp5oWpcOz2xQBGkvLRWfu7mcw9zTxREHgBxPuZCrS369XEYESoAUOG/lqv5d
T9RTWy/mnVDBsykfawniIsMNndr0/QIz2Pcm+x69hgzXcf5IRRE7siYrSgJjf8a9
v5dN/Bgszz4+/X9zKgkHyh0tZwyMSHc3wsjyHHWeiPPEN8Nyaex42nrcDlX9IJ1q
sYQQqf2engjSJl4d5V85iti+lbXE5lvCYVAY9NYHRhmbwt+rzF+FE238gTDLJAAY
TD63bfl5UhPDjFggF3RzMlXlJ6rxzeEnzvFY72kQZ9d/AiQgGrWaIBhRL/pFAvF8
tyDy4xQpwpBfl74kDJabjL2xiXkEIqAne3whOJ4sVpsOFHLI9zcUoDzCsIk0A0bb
Ayv5d6VYacQjxGu32HFot2TFQnKzOHTkRxdl14Bs1kYyC7AV3kx6OvtRUTKaAtJD
SJi0oQT7cMCjlNRZjtfgpes1xWSuI8WYePl/9CFH0/FqNqL42oQDUOnnvX07vFFL
7gyjbNeTI5XbzY7V/YdBrQmZQCa8Ki5hoB5x6LwDWcPQuLiuPv4y4jm6A54sfOEY
ehMoMXiB5ZDyN4Fq5eNH7eg3LjfAbo72NuWmmo5q/SCKj5X8cnPBXMgXJ3s/VHcr
GOHsktzCfRCRAumbTAF9vOimKWowVujBR3G/dB2gtpjkhQvfavo5XJNmk+WSIHwo
X0tZiWNktBuGTsykAsaXb77maiXcfX59boWRLfWqS9iKZv+Wez0paF6lHZghAeyq
Xzh6XqeythfZ9i9rRusjIVk/m07QiMSyl+cceGG4BpRVMfMpvBXd2untZ5gIJX2m
XaP3JK2aNzwvqidpfX0Wb6xdb2EMgSsTUD4sRWxO1/d3fJ1aVItqnNjhO5J8mL4M
blTFHUBKRUoGOXcn4b2kuz8uU12vZ//CCQKKk7UNLvJOmZG1+eCgUplXHLByHvAj
E8QJihxFlPgdQ7EhunptvprZsSMD4lP086gqTfa5v0/2kRPxyRGvEmHJm9tuubrc
Gmq1jswZX9Avz3kePTlYJP8ShhAowGpdIIpE/4QtvBByf/bW8W2UfqZuUOBcL3DR
d2KwWuXToTrHX0l/t9J6hYjpf2FN88fn9TURYmtuEkaVD75cx9ogOBM+1DFt1dfG
oMJKvpr3QgOSu7hXVpeFlnwV6GVB38tkWAd5kq1+Povk4/vP9zusmZu4DlnADjvO
LI8Up2bOhbYHJsSWkCthxKpZAbm344gnrntta0LYD+gimIuWhZsRvJDXPzd2Zhyr
yTfSdhwxvAiII1/4XleUGSEY0daZasGQdgq2zE2zqEAj3XL9bTRH6LaHijq0pLXJ
LognEhkhnDaVYyxntPT6WQGAqN6hgrfF4Lw1loiaeFn3LdUK+9irxGALmJdHu4O1
PJnFLntqquqb/rP3uTOoYrPY/+qxxbzK0LV9n1CY/NFOHxvrhhPYnSlXpGQI1emE
FeijLCmIYtLGIMNiief1Pn6vP5VTAEAXT0dVE88md+756/smqN/bD096Iq7icVkB
aqnN7j28HXBkeARgbqixnvjF2BPt+ql5M5TKafFC6ON7MW4m5J9jio/jwUUnLOR3
Q/rCRDe7W3AHn5OW/xutFI2UhKF+cagZAYNg9RQ7EZ/dWyuUiLS+jFiiHloIeBiZ
6Vd3QvdeWpTWOq1Ge20DRcdIFNxJpRBm5qQUD4G80vCDwIo+jpzb8MX4JDxFTlyc
m9oTOyp/EamEcjVOYtEbzyQCus1YkMjBi4B9jRAlumOKVFl9sOa2m12pQV+J1I+D
sHi6sowB7u7Tyq5HtBTKKC0wPHcameKi8X+phOMwvBUPN1VZqnvqe606fqZ/JdPS
7L4vNpoTnZVe/ecE4ioPYpOqxydk+aAdRX8gRnUWmUzYKNMpUot/PCmoXnTyFeZk
/u41OQD6b3ww9jcrYqEo5TmaN4t93ZxxGQ2YYdiJ9Zc7BkvG0FtgxRDAJ1GnBQfY
W7l4TkWqsotJXFtmQvtdgYsKHk/SUvh6LK2ZWXnBQdCQQ0TEQ7CcXAX203RHOiPn
MnTzDsKF83UHlI3a4BbMEVEyeq96k/ggcx4FUq5oqVoTmRPJZ07iYuE8e2GKlJpY
v1TgwXELmIJRkSXqd4bsy4BxsDL2KkshwpxBtm4TMqLrlxwyPebYqztXy+bhLBwv
twVL10rxiYfMgnKSyY9bn93Uyg+CTYPv0QBJ7b9dO0B+/E17dc9+g/JakKRfEwax
+XQiameSheB4+W+oSWTbL+SAlQ0a30fJ4lu8Y9T8bwiFmke2TInctfq2SbLFLC8D
qQtdhA6DCvT/lhLCHDmt8KgOhD/Jla0ae6CF8QuCuO9luks4BQp38e55YUSUPVgG
CZIV/oAskTXIp2QMjpAXc2dBc4SwMzooyU995UQv3WV4WdAjGDjHLnUaeiDhTndQ
d/AKGMzrrdQcyuqiU7/DmHDCP8DYJlsmhMd4eKdLCB/IUbNgPkiE/DEzKjBQkyAH
T5C8FdZSx4r60hK3cCX3rSrhLo6TJQmEtoaCB+z14Z45ToOkkMuQL78ECGk/gaBA
PtPgkWanZ1q1yZq19kK4ACGslbQ7UyitXWO6FdbOxpNqtgTvpeVQvm9DgW/2DVcP
jVajQ1d5BEBmFHmBS03tpsqLXHvVUqi9Xmhh3MLd+fk6yL7jDFglQ+TXSVK5K171
Hw/PIfze2YUbN0jSoHHLI2gSHaqNPwTZr4bzgnb2XDu85l9OXeWiqELbHbugRsqM
PYatVz2onc198vWuCTEadXfLnsauh1tBw5HAG0E9E1UqXMh9+yz2U4HglZxHx42h
tZeJyQUy4tpikjegjhnIqCw74k32LKiTXIZ9/ynvMG8HbbIpNeC/UBn5t6lYnzk+
7hQaVmtXDSC2+a2EdNbOwr8zDi4kbjf+BUbh3zMe2R4QBL4NCDHlG8GklvdQHjuE
O8Cd42xn0tkN/GM9H7lNYiF4I4CpU+P+FHOwmnUpR9rnGlikjmFg74/mCuYdBObD
9L3HQtI9qVYzUcWVE24CmOp/uJVATiI2VMXFncVWTeFoNZ0QGdULCz6SFuaLlF/T
QBgCKbjAQ5t6GQ2+lLk7GijCSj9gD8cy2xtHZs0dIm8TGgE2nUJAMsm/mcHkWWKw
6b9fmJiOhHoNcB+yyZJJpHZlpU7bZGgjw082Ic/GhI/EKQheztKuvyklLR35Gm98
xjwbMYEWQq8Tcu03hJg884mdx14+2MHjo5x/bdAnoLAoHFl8WDcIuVX11qNbyLe/
ESwZyc7DHUS4RirI7EIwv1qIvVPi5eBLW7hCkwvG4d8APzHBj/DWeNtytDI3JB6y
otU3CdUxpmpUprkOpYPeP3bEsjllon/0Pjo0+twTtcGLYg4e8mSv1L8QzXETnRLP
2mvxGinwJlqexOr14IWt4AbH3iQy09kcx1SmCpxw2u8Yu7nVvnfuqgBVUdjYEpOE
f70AHw5TFjUzXwCUuwpqJoRERJ/OnJ8Su47rbiqHf4o4sEpG9iGmriY0/yCFLk9J
GRQOhN9Z4NL55nlQ2a2TbMgjCkVKmvrDBUvtLtFH7Oem9mizatTt6XjeNbN/qUuR
M/4VqCP6/G9kODz9/+Xd2PuWcgpH4mHkiU3DzjEQ4uhyqbbPbutJQ74R3HBmTDZH
+JTHuZB0eALuO5R5t78qcY5Ax2tPOtLgtvmEqAWinHptuedoSj6RSmdmSpaIEaCy
qvVKC3miMwzqMJ3JsogL7zC2Nq3LdSuj+GEu6ApDhukcxASqDiON2XNjVJo2DnJJ
ASyQYVC7vq0d/womVzpOiPM1Xi2eJzjPPyVBTpk955ofPSp/giD+F9c1G1vXIftF
sucGijUis61NCPB0GRaJIcOAegb8W/U2FmUMx2V6Shl/PLSgPLQ0ypD08C7Uc0sJ
zNABFvv2p6wr+A8nBxSedSoDKAbpZ7oPy4fYqo1vuRDDZHkyQCoJ1BE2ZjkCaItE
Q1vmnPVm8pbDPCzqDuaNJLp3bh63zp5mTU0TqNqMlR0/5Ga1JVb4evaD+SlqfNxi
GAH+qrqFuUIWmRUpT/EOMWpr0hN64Zd8Zx0w0Vrhvz3OfEcarG6uoEc2KvusKHvi
+3I8dfYlHBRO1IunR6j499M89Rl4xMDEkqWZnytiLVMSXR2htytK+K5ZeitG1FA1
cx5T2BFu9HDQe65RZsba4+DlBNFN8BzuddFJehTBztdN51eAcUSQ5kQP+K2Dohi/
co0sDtNKk8P89Z8Xpa2BpEU2gP6H6mPhc8DBsPnCI77TOLQt1aeCuqpwlx+RMMTL
wXtCyUUaxhJa2I6fKW4BTjti8MJAJ30QZM7FVbxD6sEXKjDPjWzoPJdbiTdi/pVE
HY8AWyeY610INlZoXHhAVwhoiFvUjZDa85r1tZ68lZ6hVPBHLb3D3pZdSXrjoB7O
x+PAkvW7QucKMSaNBfX7WXONL0MWJT1kO4jsF4pqULCzwo2TpXh+jc3tGVJ5mSC4
Frkb1mvItzFHNQX3ECQtu8J95NayV/YtOLA+nuHykj/UOJDXQVjwpQn5OO+DH7XC
7BqNZAaORspFiJTzhpLTeL7FGPKIXk2DP+6ewEFYnxvg5H5FKxNFNKKYxrqZ1Ass
lYn4xmdmzTHk2ZTv3/INyj9IAHv3r8KXxZcDYExBAROwO3GhiDt7hygIig7DxcDV
BikedswyihsLTy+BN0P/R5tMWog6U6BUBTF9pJt0H26zYPgLUrlhtZjkCRMhMv6e
x+KkfL2jGTKwMy8u2KlNTHRgAtwGiAf9B118gfrPLHEqFVhtZ3HW7RodlGeCTGwE
Mer4NDaRhlH9ZZ/rIa/3RVxMn3bVVpivv5SkTU/Uw/LKnOP8RE3L5Cg2Poeu7VHf
+0leW1KlP1TBgxiraw+CLmdSv8UyHgQv9HD4A4ti1ESI0ZuhH0XdzLELGZdX5lVN
OBFMOodcKDcQ8WHSZm0uQVmbF16nM4cbFoEFxhk/R/il8bvZSTDf09FNAzzHqIq0
MuJSwB0YmLOVWjIu1nnYnKgIgCbBL6+PVKFA6S6wUOuIcDVX5fk5a+XjsTAcarLt
Ev4rUWPRsWUiUumagm+WnOl9alLGEFFf96AIx8+QjHlTOwZ6Wdxi4XW6Se4c62GG
imRwnVyg1l5ZRecpgqohhQdfnHRJkBmhJcO+YX0bgddFFIa5ACjJSrYNY9+uuTZi
lsAHqtQmooyopLtcYpwJqvGhHo0+dudUV7n+eU3X2vvCK+MsWCfNAyynQJNfsgQ2
mdwpBt4we9QXNuXE2B8kuLFeUKfh7b6wfxgisQDoMQcl6zOfyeWdDV1sw6o2fmAY
/Ejra0eDhoYTUemBfImJfapkaYlVpKbseMTiq3aBK5DWmfgZ+oVHsN+nuKvj8vLD
IrM4kxnDA/EB1SAbyBfUYt8qis/WSVqrTloPemEIVBKu/ej7/z7UjmXmZk5dv0g+
JxEA73QHi+j9O9+mTk+dVuMc5X83sjSvXFuhYPYQf+X57Ch1FH4Wk57UYm1bqGUv
kaHZ96Zafd/bLKyRUc840rD0syW5N85Mw3k8Ptq1pC8ejIcJBpTHs75PU8CBLwK+
C3WdyRr1AVz2Dk2xZ551Le5aRYItYczSlFLP4yNXuDeBsmYPhaG7FRcobHAioJd6
90dmZ6OJuDyC5btaMo+4R4SDMHVAlUvc/B5Zpgl16sHHG4wAyYm6Jafxwt11sDkk
dimMGLjXXBLUcjWpBqEsIOSRK5817/Htj3svNsvifjdGaskehPk8+CRk0kdgifQC
lbiEYfRDfYtXbKIvlMco+JLBMVIIhCZXRbIVYlem4hXy80A5RruRJG18AHplycEo
f4ajr8jDXcXTPEahA/lB6zLoBJP6Jgch5L7rqOHuBfXV/6pOyAnV2BnItcqsAG97
0yD0h9UQt+t/MMpmEyLtQQyBG/wmLb1oLcZx8JnF9ZspouzqTo5HPJk8TcunAiQL
PGS7RD+ezrrLeDDXPBnwQ3VtpYmFqRgDDQVzAmDfuKVrp3BhaMrGU/v4bu/pwszm
HO6mUcFtHUOzLX+ie5zZIstwx0op7d4xQzJF0MYPkwQsUIaMvhNKJ4DEDrnbpKKx
rR4DE0umO6y8n+AFsoARk7fV0MmvNrK7GA7f31/za302l86SXAgJ/O5jPU2fQXrC
cdn4+l+jaYRqWE539jElS1t/SAIWkdjPtaQ63TViu5RxwFrlZLyk4+WYT55aSuRW
rRIMUwoT1G+UusxKrb4NwEfe3mz1jVPkldThFkk2fieg1QUnZ1CGz7D++x2tsKFK
g4sRhq+teX2vd0usu6u0GcPiONjYnDKdDZkleOmxfSrUDWeSOQLYue49S866da9B
b+z4I/J+9x5mbESH6wNVlkZSFvGILIpuMvNIMJrc851H1iMe0wE08xaN9zOAVIXm
5htfGssXkqk59FLAkkjvKsFob4ockomMtEiufxYQwmMYj6Fr/Vie/Orb4/2u4Y/z
1iqsYr+7zrb5bhWoGHlPPhU6KEn3IGXOmZOYSRjA2T+fApbIQG4W3gDHdFGrSMzc
2abUdAK8P81MpAYmIqqvTCPsWWSn1ft6ZC0f3juqFbbz6WsP8bLhPfTbp1KZ9I1N
wn9LTuGu6ypBuhcxdihXhXpmN7nWb3CquqCktQt2OxtPCo1hI6iPzz9u1DkowgKK
BmX0c8Gmx/3JeFvRHtr3GLPgd6up0CJuaar66EmebAuXRQ+b4a3N4vXAuoDAFDXt
xQmjAyhy0VP2jBI8l4lh+FabViiw+Rgxw4mSoKOWLJS5rmq3VXfawjaNozHpDssR
KzY3WlshRtywIBpYC/Bf3/Z6XmUAIiRuBF4UD8tW1Z0ifFG9cC0jJw5Z7faQg6FS
6kLcgIudo5kCU+zAnhsrh1Ym8UvEmE6bkfEc6OcgeO507w6+ujpJzvIae0u1aYPD
oXhvESOrSmpHYQCurk80pVy/cMYT3zIG/s9aCYP0H+sCCBfI4TKIIPD46NhtZnaT
vKqJgmDiyzyssZ0yn9wvJB6bBm/7N/GptTgytuwyqHMZ9VL97qsPT4bQK5FDwSRp
jG8gtUpJHPmALc4FT9mEPtwonn1mV07NjYBNXxSBAeM3tSRrXLXYC2Cy7eQoBqdi
Iv8rJglEHtCh6CeneFJOqFM3l85qQH4gncdFG6S5bxWPlAq0D870jnwOdDt1NCNL
nvgOdFRwhvf8edhTsaAjMwspjZ9Tb7/QK3SRlPO8OOSwYu/jZJbF93Im8V17P1bS
R2d8lRVogy8nwA++RUHEM2hBb3g06C6LV5K1PIZcZvGW1hFw3zkzVV18kFWxysO/
vWxm9AsToW7YTIVqG38+MMJf9tZ1efnUVeuNYhtEOQtjRV7OErNbaqoxdLILpZDX
yXaCPT8MoYoBVLIynR46ld5/mK16tXZ19viDCAmC3I0R9lGbOjAIYDwJxNgApeDM
WtI334tpdPZgu8zt1wlb8ts/XCOIp+Z9n5hEQrT8MDrJ1cwyR4b91oyBegoO0dGu
IfU/KK4lSG9acKLiU01Vr2Fs6R+Efxi/8bKNd5/nYKAyPe5jxlWczTZZihZbaR0O
ShVeEFF0ZqlBjuq6ZAd6/E06acajH8uiIFT/g1gHJ/cEJvQX4wC/8yYMf1vCM7qs
4T8k6GvbYHGSFXk5s1ztkLLEs6iNr9njoD3GfNHH6ocSOYp3d7aGreAi5v2efg5b
DqttuUsNqdkwUFzBn9f0Qg==
`pragma protect end_protected
