// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HH EA7C,U62EF9_HC&V74\R:AP*7:K1!<GC\RGQ22B #472C:&Y&=]   
H-J4/;**S0>X>=MQ8 ]$V8@):]KYB*:;,+$27E9&M:E*2%&#G8N9!1   
H#JVTEBO)/[ 4RA!-(1@3C*$_.KNM1R<-5/3Q9TM^+QK0.\'"_@JFD@  
H?A#*RZ^("L[!:8H%2KI>\03C(8KGA9D[C,()/WZ52&#AJ^:&_!L=7P  
H=6L>W2-P/[A6O3E(S6Z.DH%(I(:#([KVRTML0L2V^QB[PD2J,!>^A@  
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@8JLCX?DV.?"(P8?%@^\<23MXAJ&N!JB97\I:#^\Q<BD 
@VGLO1M.]?=!?_CB#;%7ZMOS=WK[3(UF< 5X<#7W*:=@ 
@>HC^:QT<SS=FQM'KX.P&JR3$L1-HZ?L35)B-A?42"8$ 
@JC,4!9']%2R(F/?RGRZC[J</C;#'<E[9+9@I^S7SBT( 
@A=N^C,5D;1%<'^FD$? 4]S03NRC[DR'$M#2PG:XGE/X 
@V.*Y7>1R8!6*;/CK6ET;R7*#-)*+KS.4Z$-HVJKT D$ 
@SF2_MDH@X/C_O%+65<\4E&%@T6"%$^>*)PS_[& WDP( 
@5.G1_>I\T[MH$GK9/L )9[X(Y](H7@CZ4K(3^(@LK=P 
@%_N 19'HR+GZ2=.DS].%>F+$SV]#O$@WR8(260 G!R< 
@E5H[DDH^0P7TN:AH8?_WBK[;&7 .E>.+H@:[).9<@YT 
@WM/3!#5>;,J0M8S=,X:XLH]MQRUMG>=M"]-)J\E&!R0 
@*K_=&&?0U3HQ;'\H.YF>428S<[#9]+4+8: RXR@8CG  
@<JR,O!QZBC!NV5ISL^$2;+B-80ZKP;K-O804G/1<W2< 
@0BE>RT110&6T29F_L76V DN>Z@78LA2&T6IVI&_T,*$ 
@85F-%\!,J?DSHB VSN9^2;C+?M2T.P)\,/ A!W^25RT 
@Z]K(I<C!F>=.8#_P@BD)5+TCE\>$H3DQ;'=_U-XPBY@ 
@7TE]K:<QCQ+B;R1GX'.JL6W;3V5<(CPNWYS+#J88*SH 
@-*T3Q>7/Z@HZ4*);;=KK."VBR!C EQ(\WDID*68.5)X 
@C@.W./Z]W19-,V%R.1900N_%=G&$8-F#1M/^N,@P-X@ 
@E*.(2,<).C=&;3R,:#G'F"J:.I?9GD9(WXC=M:7+Y:8 
@(_"<[TXT=N\_4*PR2-FG'NE+U0?3FO/*ZYIS[$/5W+D 
@L^&7G,MF$?;N5JN"Z(%N[2M,;$1\[&RJ)D=8"P."9SP 
@!^I#-TY#AMOZ'&6;XQA)?7D4>$$Z!/L-)3E"P@RNAG  
@GIV2@N)H3N?PHU'H;]48OB%9^4P<CIOVZ(>Y#TV(GV4 
@\DT;&2X ^2ZZJ<2]5XU9_>ZS]'K\>Y!'I+<S"T[6;AH 
@T2L):.2T?@,JGRGS*2D-?T#9\^! YU'%)?>?^GR"IJ$ 
@=V/CY;TS6ZY;2\=V48".$?GF%0*WF PE.W$>EKFR$<$ 
@6ZVJ-LVNAET]"'F^QFLX8C9PP*,\.\T=7F">'Z*>VC, 
@=##6<XX5+*S+(5-FAAEKIKJ.UY<:BBBYCYC$2- =+8, 
@X$#*R6,T]P#O"]40YZ+J(\_U#1!:&!<"*8(/W"SU) L 
@"/YL\K):) C^&L=+S]\$ LUH$#532!-LH>Q(_B0T"\  
@.5J'X>HIJR-QM^PWO*7_=:R6+L+Q9U_US_E:+F9I:S$ 
@"Y=0'?;OU.%%OA25<XYKUEB6]M^".@:8^Z-3Q,9LS.$ 
@T]/.E7,)@DRQQ_36XZ6;6)%2"0'5J<K2RKP::>;CG!L 
@2:$-4]/Q<O*L#QA22W)8&+/#&I/M@%9(T,#2;&D4A_< 
@+_RCENN0KPI/*0[WD+Q%4#86-$;DI[IX-^ /9*R_?8\ 
@+2SC!UD>UQ0MVJFO[_]N51;$M]YE5XG6J6U\7!DK=-X 
@=U%L'TP]K3IK*_&9X"&+ZW[>9BCAIXSHZOMK?H]Y*[H 
@=A>I6G"Y>+]G<?(2OZR$/YP2L)M! P\TE/-5!M V*@H 
@<4%4"(-Z/>BYES]4OQ&*?O8ZMTWG-=;[)F>!V:^VQ8, 
@3L9!=1<;QY8+;8[2M;QL5N/^#1-P]S+<'-]3U;8R]^T 
@.%!7U:6+NVR8*^,#T07H<"(Y:$ID9H##P14*I\)/@SL 
@'3?,:QHS5^&NGR:.,E&8(Z)$:,B!9&HD$,"I,W%B7N< 
@I-* ;*\QFWH3+4T5!4N^I_S4P\=I6C3O!TEZU35E7_H 
@V$4KO!>'M!HB.YBZ*81\@S\PPE4=T07)-B[PFOFY@M8 
@;)=[2@>?2.U_ ZX;"]L6@;5'H-MN .AO#5^+H/[!'K\ 
@=LRUD6)^'5 Q%CP3$[=<7T &)171J8FBV@4A@H=4H1L 
@>;LQX;7Z(Y"IT=H[-?K9JU?GXI6B#:TS/.?D0'4C0V  
@'WAEQ2L7]H!8J6QG*DE+'0@_O]80(KE#4_!>$++(RT\ 
@."(]\5-3A<M&Y5==-0RQ-*I&>IDL?3</CJ"KH=4=;40 
@=]^K#(7/(I+@%)3]\V%M?1HMUW0-_M]YEZ<$J_TV6R  
@@K$05?XH!V+U#_ATB84WBCQ6E[*40BZO^(18KNLI7I0 
@YGI (5NP&ED#^K- M.)A#TS[<CO]902_^K;\YHS7T/@ 
@/A9 !^BVBJ*(0[GA7;QF)%>^?)%.2'U\O6G$)PIC*2P 
@(:(/%*LB=)E!6HK6P8SRSZHF&@^AF/_79)U6C4#M_5$ 
@>B,4WH4F0&*Q+GD#,Z"&U!4##,]<304XH.RAEOE<420 
@>[:*+1>%.)10[1BMG?0DE&X(-XN\3 T<&QT$/B$VA+D 
@K5E-@S;XZ?0T&D*6U=X^ZH/NG46$.3+='9WQ&2G#<UH 
@H]+AKNZ-*3><NG'2J7;L<01A!ZB_SV@S^< *5WTTHFP 
@.,IZX<8R(/EVA]OBEHG5OQ>D'AV"ZP*\"EV0R\RN@4D 
@ @\,8#*%=;*K=RPNS=>A5!;3P*F#'6WLCCW;?/AGIUP 
@IY"0NKE*EHGL!S4D4]L.T-1B(FN?TGV-R#5/[38$!C  
@D05#G\<9J]TH#Z<%8P"R0G+F@]*LY$?T*Z0H9?J31%L 
@H8T,UYLBI?V=,6QO%;3PQ!%\".;0N=2.30AI.WH%X'X 
@%3[Z.MGB\F09E WPEKH5OCF(9T+CNA$2NNC @>L>X"$ 
@2OMKV3%1@BQ%J*MO[97KZ1R4X+7CX@OLAEF99VKT&50 
@BH%1;!!"@P$'3;$6&;4'6;*3NUL?33-M-5LDDHM[AJ< 
@9BDH"6QC,/^S S;:1C#0E^G3 8;'07_ZRY&HCH;2WQD 
@&DV/BJ?7B=HY0\J;(F80N$0EN>;)OU6;5">.=87E6[0 
@G])I>8L-'+B;3,;1VR^?]B5-&"J;7+"R?W'L.[%J@\P 
@A9M ,A1N0ZZU!)I;30%8WPJBW-))/^%."7T1[TDV\QH 
@2D_*^?6^)#"-_(/6V3MK46+I<DKG$\'(_9#XN>0+GH@ 
@Z%;KO6>LI2JBY(+-[U">2<)^:9P(@L62YRY^K#E/^^P 
@N FH:KWM]OHM7M]%/QG>?>AGG#:KZ'8Z"="*&$#B7]P 
@$OM*E,K>])6FR=N+:+T3Z(HM9)@-E,=6DZ=-^MZ[?,D 
@%MI[4)TQ1O@)L>@#+,NPB9/1EMN(1#VU5#MXU/G "KD 
@&5%A2HD.S?J=G]P+79);AQ?/5 #J=V,:U'3CHUU<Z)8 
@_8.(@G)V#)6N" ':FM\!;R#&NHBK"O8%3.\,;.973O$ 
@)IZP9)LQ,N@"1,>%/3 ?.7$PX2N"_;%J03_E/6(@3I, 
@Y]UC"F? 'X!/'[I81O3F;G^OT4CLM35AQ$\_2+7L= P 
@,>%7KAU)]*G?C1MV>Z,OW%-Z$(P0^U/7OCT;YK:C<)T 
@9:I$6:128+#&"*/5\F%N(W$E^]F!38 .&S(:<!$,2S< 
@Y*_J\U&0N 3R^0:JX60 ^:][H66J8*'^]5'&X+<);9P 
@-P];K6]W$/8:(FE8\L5IK)Z!&R1.F]^1=03M#^Q:+@P 
@3\ +NZ#A=H?<RQ/M2N5Y'>%^3U"U 77-]B),/=7DY;4 
@54FR[P-*@=X95*ZX4-92K/)R%JKB!>8XE#&NI?+.%\  
@HWYO/G!5Q#@)MJWI52\.6>CL)O?&3W(DKN6,VU?%K8X 
@SE-)Q7-P5DU-0S-T10T<@%"3W%"X[-.C_9_1P-V .YT 
@CZ+@9U(-<%3UODI'MI?5&Z'<9CMJQ4&'.U!39U8!*^$ 
@S&U355JOF-)^8!$:VIQB.A46RE1=+%+VYK_@_(P$->( 
@'I1ZGJ!]N-TBLI.L_(82]Y5E3C+ \(+&T?9 ;F:V]7T 
@/R9ZK+HHS)\JO9 EDW ?('?',U!6_\P)-UR/RX+,.[T 
@E*,Q?'P%A/0W^%YEZ\*F=,7I$NF5[^Q)O*/\P;[D-*( 
@97@K+/9F%P?_JZY)$J42BG^T1M8"8T[J3:]9F2\!,XX 
@SVNDU8FW31Z65PZUGL5Z]K@8?1T/9($LO0WD3:;3*&P 
@AZR+Y@,D34<:N(8/JY=C"\7],LEDEG:F JD^\=7W86( 
@.K/GYWD)#B]TIO;'#+ 2_*<^N,U7\9!*B3N59?+./&0 
@Q%AJJ[15:^L6[M_UR8J?X.@31M&1[M\H8^RF]UH8^#P 
@5$5=GNN@A<:(7H<BAOZN?1:@BDT^965(?&*]&&S$$O, 
@2 WO'J\/DINA3S$,P9HW<:G*,&)P]LA$?J1)[3>=_*$ 
@T=G$KCI=JQRX)$K*9S6]]NRC@$[IM<+\&;0D##]3JP  
@Z&;CE8&-X.U"<RHNA-P%@62DM@C^A2W!/'DG+1Y?%]\ 
@%8>C(9WWE5\9 8&PK+^7!?+%A"%>7?8HTB+)0 D]L?D 
@#1LI=<7-^^=;!TVF$+&;(O8$SS2[^/2T^AWW[/)?G(L 
@J<%14'ORKHD(A]DL=6VEN?VIYPSI[7!8 IB3I<'L,*4 
@GEYYLRP7WW4H#<2T=4<B?NK7Q(V[XFXP8 R*-XQ.I+T 
@GPN5V)2K];6MTCNE%.-BAU8M%]IP%(KND_5U%:-<W$D 
@T<LE$MHYX/32QHT9XW8AK2"#Q9:)(IAJ$ISU%F5''S\ 
@ZJ%XL>N)Y3*_K8#3&&,GN4M9U00^>VJ,: NL;S_:W80 
@I0*S%T.M5<>L M)9"N?067(L,71!MI=XTE"M%(%9<"@ 
@YU,:I%%=4MDS#9,5A\7+D0DTE/7__)7UM&,CXQCIGP< 
@^$HZ=5-I;_^80:3CQ_*M?$_I,_$\)MI%Q&C<-<!R)P@ 
@2%R2J:UD*U[$,F&..:;(0[^GKA'GT9BHQG/Z;5DTZ+X 
@4&IIJGQC8=7&3'S7U>+4_2^\._474Y#CMX#$!^>:\S$ 
@[)9'8@<&(<V"70+/VP)U.*!=L:MH3NNF-F<U:+'-'-  
@NN1S"0[")7@B0FJPU'WRA8M-MI:+[/]-1'!ZUL1; !8 
@CR7L17.^$#W.70DVZHB(#?3LZU6!)A _.-IWZ2 0C+4 
@!?Z\Z>A>1 NM**\MG9A9;<//^C;$*(J&&Q"G=>TBPL( 
@ FMP&R6G;3U0,[ZH)LT!&X5=D59+C*!"$F5P@R?;I=< 
@L=V1#]T_#?HJ^4T#9ZW.Z:9?]B[? XT7747R7+NL!]@ 
@5N&9R=9MHL+2!B)HA8H_<*BO<;!Y^X.&3)%GG--'.R4 
@/$#Z#1_8[H]K/+[.1GPFTRTCGRS8T8[A9J2\G#WN26  
@;_QEJ(+\6W1.D^FXWAA9VF\"[^W^7\H Z <@X]($G28 
@N(S-NJ=72]5? -67O<XP$2LO/E>6 ?5Y-1TL48+:Z!L 
@-^G!_B<25=ZA2:XO?8 DYA3S/"8+5)/Y^$Q@F(CL1%@ 
@[2IY0#>AT\8LK<Q-P@ANHH8;,[HJ;.G;4;VB['<_0_T 
@.=:5W@=?%:K^_QD;X!0[O&T[4"=L)(6?>E,FNNB/-AP 
@^2_L3I$1X\WGUEQZ[ZP#8Y)&M5W^8 O:N=QD9,R)PGX 
@,2IQKYI@KZI@GB81OL]7XSX=\Z43:7R*&F%:H8:4E2D 
@*;#KC"+R#MV!EM1@P])VE:ID:L,9O-),>F9K$Q.;K7< 
@NI]ET[%)>D=VM9>P0J/5#-B6_4@[#ZW(::L2WACXX6T 
@-"*Q:FFRS2+S-\$[O@!F777E-OM&L+Z@YN,5%S[/V'$ 
@^7^FS(1I.L+1TBO.(?.4ZX';M7]).TWAN\3D%87,EB( 
@(YDRS =T5Q8_\.WA(-X&8=U!R/",A.-^DAY;;\@#E@T 
@/YK%U\W=ZRN:7*2NMBE*!).D"TR7CN62?HJ* ,A&G*( 
@/Y1*# 5@(AD385Q8G0>BB3K\K$A< C7(6X@R3_"S=WH 
@7A.?9&)\F#^^^VU0GBA]RB\RNAC3Y4FVBWQHO:]+:XT 
@BJ9L5G\?M0CD^T=(T8(O['#4RP>Y70'9!I<5BLI%*(T 
@H7D @SJ>9K3NVLZY^.\&0LZ#$4I7S@-P]FM2*D!!4-4 
@5>X /37Q).7V0M,4_.H65##.E&W4]*[(R]0)[#BI00\ 
@4P8NO66:Z\W+7)QAZ2[B+!LV ;>5QS=T1S,/]JY(-X  
@;,E-(J9(7;'APBXI@OY %F.]L8)>Q5*T,\]&(H.\?$< 
@5FC9DJNFQZ1HBV?59)HN[692VES34?;Y<71'2<M4%9D 
@\CQ*]39Z[>6?Z]R%0P"JER3\O\6;^CRP-4@\112V"A@ 
@3)69YAIK6._+)U5]O$ZK?J:C-V[7+$8*2V$WH%KNV*4 
@XT$B: 536+/(13,.;$7ZTO]2[ZXJX$Z22JSQ<']0*K  
@-N<)O:]Y&Y@.\390RA;/MC;10U1BC\P(*9-RA]F'ZI< 
@^O=[.X(95V%\3Q%Z<QDIZ3E.7 & V40L\6C^9J8/]>0 
@F=6U_!0Z4KV2I83DKSZTK )KTNZV>'772@^R4#-!Z]( 
@C2]:+\T[!.?BXV?JQ:?C:>5[UPP3[:P7 *+;:LDZ)(X 
@787TH]%E[SJ#$TDY>P+U38,/+:5_Y4V?B5*8WG9_&M  
@9[V T#F#]!TI/ZSG)AQ9OM^HY&%CLI$ [74;H/)=49  
@-@G0Y%>KHE?[Z)W8 ?A>5CW\H(U$_A 'C+=!; T[M H 
@BSTC4@8@.Y+;'+9,.87CK\_25($EU)Y_H L,1X,[?)\ 
@0&L&DF"F]OX;B3VF@P]L$&#%&PP4RE_13XE+Q]B(,RD 
@7WQ[Q882I9UCPU6J>[9-X]L)I*%6O&Z\1--2_ "X)VT 
@Y((P *G+K'K^'(:.(S6-#R2\K0PS=U%_)C@8Y6ZRS>@ 
@(@!$4@AH7R9^$_'"KM?2C+*0F/E.D .H.2C,WVPJ2BD 
@M==I@%"%++_W-+;6UQ=;8!)YI+&/[@H@:G>\VT]ZYW0 
@94UOL3Q_4/77/"7[;NR W[SWR6.F.0,@J@#3 P76!2@ 
@$I1!<5HT]BNBEF?N_YIL!O6/N;657B$3&(4/'Z%]!,D 
@2MZ.J;#*3R'&&4*2^!@3>,D\#!6E23"=-<Z5;P+QM$  
@6:A3<3TR>MG!";-J:]H!VMBAPK6L'%A)1@@SD&MJ7-( 
@6NH6O!.JZ@\MZO=EL9E31/G=RW@];B'/4$>2:FD %C( 
@SE!#!#7"3"9%L":6\W/4;M%K%M 6%76JB\2!EBL;@C< 
@^KIVQKTU PP+5,OD/N=XGE))Y&/Y2NV/E#N1P<X"(_L 
@=I^:3;*\IU! &26)!@C=+4Y6/;?^VLCA;"V? 842FWP 
@H8WVE9(52R5K =^&JYG_C9+MD_8T_%?R_WR4'0\YS<< 
@Q!GT_5H5J4-TJU!?[+:-0U\.K]J/>^R&(.$MR\%IAWL 
@0F.I&PD+IQ;KVM 7A8=JER'HGMTT127W9?F\/MEOTPX 
@M:2U'49Q["GUA.J1F7(76T)N+X)50!,IM<!OQF#W3T  
@PUWC4($L=.P&1RUIG8;?+TBR25N3))6C.N/^/@]BSU  
@N*L_J/33&(N\BL&;)-9^?1\V<'WI:8()>6)0OQU@97< 
@U1[,L,.[:BK'1@KG7%*>GDE?3GZ1?MVS@/&V[U6);;  
@:6@DL L"(R^:4*7-;\&38;E;CRV&M'UTBF#&<6L(X^$ 
@:&ZF\ICP-S&4C3RA3EBA7/L*NB&N!C2A=*@Z/NAQ4;P 
@>WB+N_6H:\;!O+0-U")928_\S6MU"06R&NP5RX7H(44 
@6T,HBRK"6!R6IN9_!S:+/XXA@)=OK^6"0__ JX7(4B\ 
@]U2-];L,T9U>V&H2F>"9$ TZ'@PN5#CRP&YP+2OQO.\ 
@BZ:;,_=;G6[XG_B6P8;WWR:4!>]>W3D#JUL0&F,+WA@ 
@P,4[J8;P!ZP?K[" _.8]^JLVMN!9CT%5W&-:E:R15C@ 
@(@CNL&IW]1F.%7PUY!22LNN(P"=K>D4C>'.-2T\:$M4 
@'I_YHIM&##;Y09HCJ ^JF_QL!+AM\;0<C1UL)W_Z@*L 
@.MYFKUWYG5*+M99!K)F 5Y-":">"P!/.NKD('G*(WVL 
@T88&Z^HMXTH^0.); >V]$R*$96!/7+%/\E@P3P@I$AX 
@KNT&=/S?N0W8K>>:(FW\$4F[*('I-([CV:[9OCA2T_8 
@;?=#.C1%:CL<J2X(GE[KUM56^GD\7\3'=/A5?F+\;G< 
@(LW(O6EI.L3BL>!\R3:@JVP^$MY>SL>MG-#GZ+S-@P, 
@\LM26%-NY]DC9Y%;%XF46)G;=/>&DWR#NLL*8MW=E88 
@+9L=C?V,NLYFM263,-X$(E:;,5-(&%N(-GL([ZM;=P4 
@EXT!9^Q+>9G_E(0UKIR+]%@2>,(*^X#>$6!(9C#L$*H 
@J5+J1X<@Q3-?8GMJ3:?"]]TF5004-[5_\K N4FYBA6D 
@9);_?_>=V:<^M5,7#UU]"DN;FW.[0"AIEI$B11P4A3$ 
@71'VNM3CHM=8*K*D<4G+=I+53[\C(G,E2BA_!AZ>Y., 
@OSHO"$@FM9][$BA2*!QC;F--!BSY'RBIZ7C/ZMHY'L0 
@*?$OM1_3\<\+]^\**R,I?]X.OJBY><-4R"IW88\>)0$ 
@AKOKT:F,]BH*L-_U9;P8@"U<);9LW>W$'R"$WPIT @P 
@XHWC?24O] HW],4#S4&"@4<GK \MDLN#G6>A>%2#_JL 
@=C8G:#^Z3TQIK<<<K/ ]9-P/#'&R9B6?LJ<._GVF]FX 
@%>1+QGVQM?EF(F-(1=>TNA),J2XU9,5$$B BC>EVP;8 
@.NZ^KD"NK:X"-=VXCRT[FNO21C3LK\UZ9%A0U26AI,D 
@,)PVSV,D8TWH+;..O)A8<K=S7[TO#'2=Y&TA@"!HOF8 
@<,&LP9>)Z'F 8-9\HSSA8LT=V+F?1)_;?*6&()SYT!0 
@IU6/J?M/@@'X!L30-J]Z8*3UU\<*S;'I=]1(P<_">*, 
@F G<_:C>,<-[;TB6Z)U*S=C\$&(*&!K<O(\C%[T)?!H 
@#^-GN $&X.]QD7 (&O]V]4978WI0[J:\.\[D::TIQ;( 
@,F[9^,0G:;>E=X RITMU#'6+H@N?3,.KS1<IM(N-IEX 
@_QLN#3=]/[J\GG54>#[R1H@XE3T8!*\!BH_B&X ";0D 
@E.3.@8KXOKK""93S/JQ0>C2F(T;5C.0LGT;3BR)2L4T 
@;JP=&T%>JL1P9<I^K#=H>]BXT\K&K";,/F1 ^WL!S&  
@BAD8&B=0$4Y,<.WYS\:$RI(?R"08_B+QQ"K(0I_5 !$ 
@3L^!)T4G/#I@MZD_.3<8^J9'[RH#FN@!APPVL%DF!6X 
@.,94Y/2O%T_,B)6 BNB#VA@';K\+3+X,1SI6 9O9\%X 
@W%&[IN<MD,PTT'/J"N: -9;T&G94TN:&K/VO!^!NQ%8 
@NS'?V* T<UZ!641;)"(R/ 7JQ^I>B%TWHE1> F.)_Z$ 
@4>+[#!)..]6U9=:P&^H-*?;)7S$@G5IKC8MZ!(\:)(D 
@#RPCU'0?>0T65\FT^UVR2%S88,XT?(]V93-",5"=#G4 
@VZ5D]B!YE6Q@%F#2=W &G.?)D#;H*I,O %&^>0ABRM( 
@#1$78L(!S> "R)+*O\CZK-KP(]7F]UE0<!#IG@E1POD 
@>Z*!P$5Z^8@5TG\VCNDCH?N]QMKSGG/Y;%!<UCJD^>P 
@0YM/@L"/ 1T(](,3#T_20<V$J DD"IEWA+1_F >' JH 
@_K:S(U%2R]XDX(Q?85Y7".B%//GZ/G7,ZKE#+U^27H0 
@)<A-9G>;8,?OA\GXLGZD1U%;5"PW3' H;Q;>$'V94WX 
@"#+Y-ME%()]B-5US$?C^HQKR0/#"Y01W:[#F9$G=1Q8 
@C9=%+C*R8XH3NXWWD)>4%&9V@220XG8\G$\%HGU!X6( 
@W6=NWXS"30WLB*,")FR*&-SZL#M!>@'Y4BI'V>6:]P0 
@EK!D,?<=IUQMSP* :@,/^1'I,!:)Y2[BDX?LYMC;MM\ 
@O5&D$DF 15@%@SXMO2$)@R1_=HX-BH&[E73&/Y!APS0 
@3> )ND1HC:FCA%F-/=Z$:@_O>7 ?>N(X3 8M *D0KH, 
@)'P]"'QQ/3@YL[32:*T(Z">T*<%ZTD:5F/1W3%.AB!  
@[V<>&@[6T3(?=?K!.T# -P1)9O&Z75/H^X,8K:MG/B@ 
@\1=QZ.N+T8#K8(TT)G'$4*DH/4;*'M=X0.AB>/)/#U4 
@5"0S.J^:*H@(2CG%:#"(3,,G60/)=P<9<$CM6ZTQ/90 
@_ZILC#556I6-[Q]^"TM0HB9J)\S('HQ#\WP6+FZBHHH 
@Q:_)#JS(>;?PTU>UL&:(T/JO#)*T%O,;G4R'U]!P-4, 
@+Y5 <*AH&DF,*"]F0B$_/6?%*?X2RT][*IU=/M"#RKL 
@ K?R?/1LTP?0P>4I[X\B']H$B9%1PTP.F&/-G@TCB]P 
@CLH;&49V'0[1>C%QQ;KSI[R<8BNBGA:9.<2/<HE$Y2H 
@*>=I5%.%_20S&U]XNW(A\*1V!C5H'C8$P_K%(2KP0"( 
@4%3QHR4XWV_4R*J)=;@?LY,Z?KE'\]=>^:7K]L;91UH 
@!/$^WGHE^I*-=\L\SNS0H99PV<+O>:7_@Z<%S!=.UAT 
@$&S'G9@A*"Z&]9KZ\F.H/69R95KM#N>VP_$!1+> C\\ 
@!4=*&:P4R1;=']N-6_UU*[_(K-;A$1MPQ"5-PYN7AQ\ 
@VE3[3I9]^GH>_MC//Q<=[-KR-)#N=?<6<92OM H47[D 
@S3I+^Q&82.%GV!=_,HR3P<YT<""T?HA>*IO.["_-X?P 
@MPJKVT8^]9<QP+!HG@NE@1E''>I-NFBZ.1#1K[9-,V8 
@3; E/*R"[YPCCT";,=5)?@8F\^!@5(;62'/!$#'R$0  
@!Y6"AV2#U0S]"P1/E2\$2YX![M+XG,+YG3[W.4ETMG\ 
@7$=Q2*@D/<9;/!78LBI%>0+H!1<1_#")([2T]]U!IWL 
@NJL,IW B0YNB1*^',68.HF%0"L87\3IOV#%PE2]99.D 
@X@W8#C2>,3G?E4#Z)Z39/"UW5C*PAE<LW$;%KQ>$I!P 
@HS,>S?A#,_>Q6._@7_6ZWV TB2MFX.$,O%P6\#$^<&( 
@*([Z#7\(*71TUP*A?'L-FZC$(@0.- AE?%YT9(*ULFD 
@+3W2EY:I*7XU2SA0<D3CB_J65%!KZ^Z=X)GD"_B@+OT 
@ABA>L1C5(RP@TDCCQ>Q[;-6E@$",XK9UI;T.^;F]_@T 
@NI:AF4,Z*\$B@=E?%#UFFU"9LD^]13=,&T(1N]N2 9\ 
@#N?<EX+41)QB@SSJS6IC'_([$&]CK.7#&?ME5<"<]2P 
@C6[>JH*_T(/A&M5>1TSW.E-N=!PCC/<1Q$R)PQE;KKL 
@\*5?+(>TB&#.J@;;KJ8GR,I VL"HB<-5W "CGPN^^F( 
@QF2)?N?I8KD[Z:83TRM.$).3O;3LE8J4ZT??:O*E5UX 
@Z]G OG/SHF:/8)%I:H<0+A^>))5&TES/,(6K723XY/8 
@J54R,@=5==U/]!%LTQ!'^QNFFZDYYY*!0)(NX++UZ/$ 
@4-A$H+>/)-(*FY8D.($28N*K9E^<=Q%T(X.EO-85/H< 
@>MT&OP*L=64WE!CRPEK!FB-G^57ZQT/C= ] PF:3>%0 
@ 2$%QGJ!2N 8')&]LKP6:;"8J+X;EB!XSR,"3!Z^L,4 
@"TG+UU#5;"R]\"D'2-&]QW)>*H:'.62Y-#*MR80C63$ 
@:,86C:GIO2&JH'0ESS>HWN ZJ%YLR0]!SG34$M6!:04 
@6=^+8-6!.[V1('QCPSB/K#97RNZTP.<;2'#U#K#Y[/X 
@?6M ,&!X5)=IVU\P?$2:FM[&&K4VV$H6$4?>'82>5A4 
@P,WQS_B95DU9N=!76:";3==(^ >&Y0VH?!X!R6Q8B$  
@36!"1O^I).J$%FYN4<P<.59];4T'B9>L[XOL-J3K(+L 
@&0Z]="(KY^OLJ(4/](0*1^Z=F8<: M(@C)QWH.# GR0 
@#O1H=2,2O74?-R.-?F;3^91@ N+3:32,7V-L1P=HTEH 
@#Y""N@X)?=^!@2%&0G<$<"L+ QN+WN4IZ#GD^UQ^C+4 
@=U6@Z$!Y)G'2+T1@QMOP)3\'YS']&$.(1PZJFYA5]W( 
@VVYL];D)0.!RH[ZYYN;B%PP4#N<P&>OOB)ZG'</(D:D 
@(#(.E+JTWK!GY)\!-":T)MO&PWH_@9EDX..D<GH# 9H 
@ .5\\URD+Y;AEEC/2H!TNL&RL<N\6VVZ%@^+(N!G;5\ 
@$=4#"$0<^KPJ;GH\WT1J_:LI-M10S _) :5UN0@Y@KD 
@N@@]SI1;DR6-GWG/P@CU7IP"=,V0YE27E(RIV.=5K-T 
@\59_N("'M:YTI\O+,T3X]^!$?D2G>'.,B&<5;=J^LC@ 
@"^%#YPC-K@JJYD,=!M1IODM#&+PG%H#Y?;C9PN&(?0@ 
@)00?U9C9T(B;TWO4'16)M6=353\\Q.%$#EMMM.7=6BH 
@X>! [:LGYEZ<@$L=#;19*>YW7^!O7ZFM25Z)V2'Q@?8 
@N:":41\G/IC<E4VEZ,$;G=[\%5\RY%W9.LAB3%"T(>0 
@9G31MG5<I]/QQ3YS.I>9(Q0/;9_Z?+M"L%'">_3O>&D 
@.=9ZV6C!!_NG(L$YX48"ES>Y HJ Q$'BDDO]G^VH46( 
@<',4XVQMA$^WQ>1*4TODAI=M,C+@-H5>?/55'P7]_&0 
@QG4[CB4+1G3U2#U_$NHNS,KN =V6]=9/&?4 -G2%L[( 
@B&C@Y'[D$;BZ_Z;X'X2%IUORWG[<\#;]KB+]$$:R>?T 
@KB;=-(^/K8"3SMR]T$K"/,'FAM45?)C]P3F6])1@1\0 
@Y/Q,<0'T=-ZO#?(!OIW53KGT!"W"^_MCJCYF5T39T"P 
@:4!&L%S.Q$KY'RT]:08:@<U@-(<LI5-J7CV6=:FNTHT 
@%,,S<#9KZ+9Q [-[G^B*<X#]8]8Z/*BL4JGXA^X'?.@ 
@FC,BZ<%"$;<Z7=+HY7M,QV$II[R1S95NO\_"_\QSJ;X 
@3JV#'T1SZ$&RXS\<_>1 \LP!22IM>25X%#V$&O?;8-\ 
@( 9+H69^X&W@M;]KY6T*.,]@N2F266 P^85#9F)N\'8 
@E=I7;RD<)XI&%$07([B]Q$FGY*0(+P]!_9MBX$R3J^T 
@# 5[5/QG4J6X&W"0&;=*@M,UQ?DTJ/BM[M$O1#48!$D 
@,K?QD4ZRWH[$ FFMVU\Z>4<[],XWUIM13YVNZ:[9)"D 
@E:,;+20?/:=4>R4B2/-S<!ES.<6LT_J78)MZ,^CJC'T 
@8Y2EP@3FT+F02$5[MKE%I=LO/EV[!EW\ 8V5L'9V-2\ 
@I$@OUH!' @MSS.Q99PGHNX=Q[H1Z6%.:VG3XL%VE;Z0 
@\UY(((JKX[!GA.$\I43R<_NJ+_!<B40>E:XL2,PMX:H 
@#'&DM]-8BA4?2L1(Y!"6Y*"L%JMNN^>O_UR8*$=3Z., 
@1YK@L3D'6[UNQ-R4EH(/;9UR'!C72SR:G+/@LVY9#4P 
@&" %?(0>;.QF3!#D.ZR/@^@PV4?7[=R4F)RG61/$\R4 
@:XF<N:]QZ$P=3&FEY=81*MBH=@0KK=]]TX/DTL(5MI4 
@V$H,)>%02#@LJ-/?JZY_BQD<AR^1WL#\:"XFQ-^VJ2( 
@2O]4,:G<;DIVCR?![P'<#P:E.M!]=R*Y*8)GFZM3)KP 
@V)1F!O+INK;N_7B%TS)XJV>/O<'^]0=>--1R/BWNCAL 
@1D7RLF,]'.,[YMH=I]^TIO$ZAJI=R*%I'H)Z.<&B5.P 
@#A=Q_)I?M\$6V-1V>?L[%?"#J&O)1UU@F J3>Q<Y6BD 
@A0DT?D2.!<7'8I"5(=PFRF]Q'+*!'%5W?OJK"34*V(, 
@TA*UV9CMQ^]EZ* *,*W"W1,DEMG/<FR\LF=1RK39Q@X 
@D/?O^>F_$V4*%?@!NN@@_IP%IT!@;RBRWHJ(AI?@Z,T 
@H<PO4W65&,8+BR)%[W$_[A=5/#&\JY:7<$EYNIB+BW  
@O"HW*Y.UC(HL(N,'D1+Z+=TV%"VMG #L@72DPR\T^U< 
@L9!"(#+NT#&,? (8%R5]@41%SW* _>86[)M^Z%WV[YL 
@04@VGF7O*+C/ #QD'R[UZK\;*>8FQO;&IYCD6F.P*PT 
@Q-3"8BNB5993R4;L8CN5P5#=A()EOA06<X%0=A*QXD( 
@]ZJPO<D.)F\EWK\:,-D&%AF)HGMT3B4#8,#8*FCD[J  
@:8Y1M=V(PD>F"+EF)R*,D(]A0NN  UJ=2-#"YCDTVQT 
@)GVRC4'LB?#8H:(A]5O]X9KTXIYN\9.HYP\-4N#B.54 
@N96>(LJ% I_?Q%WU>U/%A"?C>K."O]50G+4>?H\_?FL 
@+"%ULA*H#D[&/DPCV7STGM@@%+IVWF8@5A<?<#RW#AH 
@\*KX3V]@7IR=$AX,+PD7Y$7:N&68! 81B#[PZK3X6[( 
@("4-%K>4D#>[NV6L[XOG":.*Y(*8W:-!V>[O:3?B7.L 
@W3*?941]8Q (5JG^9 +G)^8.W0,$[27OV59R9UN:;)@ 
@PS<$<Q;T&^%9'9L2ET!>760AM4S((N&=J4=HR5 G7!, 
@(B4!T'%8:D8EI\IARAKHNS=N@+.@%Z],7[T53Z]C++, 
@SAR+;DXO=]JI8@-0\II24!SD3^( "7OD@[:HD;@ 0J4 
@7Z*]0_,N^>A2Y<MU-4Z=<WQ#04-B5,&OT?;1Z;C?EV$ 
@B7,=G@#D:UVPL<QRO6P8$B!"VC*H$Q*:K'Z([,5;]6< 
@IEAPB8\[762'@]1#O46VTLG\+@453\1*'V$*F 6P)^$ 
@3' PGJ\'!?"\'$K'KVK91+@+?'[,UL)]QZX943LJ[0L 
@;I(YHP!N# 3K-NK2>TPN/]_U#I!=DG$+WR*]$%.=+ 8 
@*UQV7\E\U'L[U34)"B/$U2=>^2I+C^KOH"<&!_OO*,H 
@"QF7M#=VC56@Z70QD$,8N0-@&\('ZJCE.]*'1V<6P]L 
@4W=DLR!4L 0\Y#5V;=@)6C56P,8D^'.0JX0@_TK$/Y8 
@%EE=#I&8FD4?QZ6F30]:!7>T'?KX]!JW2OWU.H@O#>8 
@8QN*_E=IP>4!@M(I[8DTK7#"(.>K#*SOP/KA';/0>SH 
@OD^S'BR.X;W@V$:GSII'=LJ8HM),<&1'58C*/E.MK14 
@[Q;1LU'U8_9S@H";J.)_X)F'(8TT7X'U_!:>'6FMU4< 
@?/A8W=@/>4T(F-&R3A4[><EWU$^V(6!L LL\A$=_$AT 
@AQ]AMO&#+*+7@E+PS0893J?@&&B_HNWXOFW,L%XNPHH 
@ =O9>HDW4Y-Q@^CC#",39UHI,'B&'PX8AO*/E*J3SI0 
@I;I=*"IUMN[>+>WX #^AL"*".-:OX1#C:G-?:;:^'C( 
@0M$QP4I_96RF%+\S(K24/ T2;'N\_VO<QD4"_.!87 X 
@84I08^M.,ZH5P_7D(:LL(9,-27:EAY+H7@-_5AJ4PS< 
@7]S?!@B+%N9<%WK=?\AJXV#Y7@\U:"DUAO?.KNQ#]EL 
@4"AZFB8N'ZW85MY)C;VW!H@^(3[:%\3\VK%(-XOKK@0 
@*.W>5X(>?O2N0D-U'[M'DH9P4W>+Z)&ROS+RR<FXX[0 
@"GS$9H0SI4GRQDNU!>U-#BC>W84>? N_'R/"^LH-_KX 
@.N(\9>LU%"@\']JS]*07W)B8(QK2%BG1#X^OK+.FF%( 
@*)H5^F7V"?'D1E ML@3F8%7:#%H+2Q6XIOOR)U)#A$4 
@*(O/>LRI6IO?R#X'"6805LXKL$F&YP"JK29YX_S%R[\ 
@2K_8DJO#D&)./!<BU"MC>C_F M1M"QV?D!V0+?P>(L8 
@BK&A5/_R<+ 8_*[R[[FY;]E1+>DDZKO';H4R)YHQ1?4 
@Q;D-<SS.6U*':_9\ AV\W^<40A0("<3>LC& "9+%R^( 
@HT&R@.#&40 N)=OT^ULDX5)V$?:'FRT275I3W(GB5T\ 
@ZZ*M31\7:.\J[B "'U=:B,ZB#U!0UT*)'X5AH$:NW#L 
@:O.4R(HLTZ4L7CRS=/=6F_)^@A&7<.".J*A;J;VTB9, 
@7,I\DU^^\PKH#_-1FI[>@I<2B@2NBQB^\(.*45J#SI0 
@'OU[9%7K4 SFY/SV(YRF20CPPA5\A7+(.QG0M<>]D(0 
@:?<M96GY55QT=$V[P;,XQ&(.G;Y'46",0QM\DI$YUXX 
@R5O&Y$?GWEC-=6P"/)VH!QFR<MJ/O4YJF>^J1$^!9$< 
@[XD<Q0_66Y*':_+=0U4$G1R/L18;J03_.KE=(8"L\T\ 
@:<)255>SG"_J[\SX0H]Y$IT;;Z;@=5&JQCV+I(!+!F( 
@'WU'A_?SUM@2C)>0SYF&(HJ6O8RING+K<K_I3*:\W5  
@0_M\TC'QVU!)RAD)@;=W4/K+_]'2=S"X8VHD/-_+2ZD 
@A+L@MP8<AVYU_!WZ<+G%6MM!&$>@Y%3NYLL+6@?>PXX 
@+#U9^HK>]8$]5T *#->X#?1"P1XA##&ED11B@N@2$^8 
@\O-5D4L,(<H8F[O.8]]])G;<[@Z"Y3F3O8W&)9)!:WH 
@44S(2Q;OGN0@>9(QH.^]D/^6RX<\LW,^1)6\;(#80]8 
@#;)N"#96<,G,,_"=V;K[6;W'A%9SU706F96F,;8A.., 
@DM@5[>N-(X2KA/"(P'S\6:!8 9$7/*3*O,F59Z$U:'4 
@8"("($N_G=TC9)DWC1KBYA-1 (G4HI_8'4CQQU2Z\FT 
@NKRJ3G-UP^-79B B)^>J]JM6TX(;0SA-N%H#T5S!Q^  
@O^Q_=OYK,H&/,XCY8*V<_OYM<F(["!7&4UUA<8]OD3T 
@1?8MK9E,C$7"/_0)HV5*P5U$')M'C_0A]&8$&?@&J'4 
@DQ*2/FGR^5B-V6<G6-.1$_TL$\YOX*&/E;$&<E&FY5$ 
@)?*1*D):R2.E@^-@##+WPVW/KT5D [9B-2=6!F)6A/, 
@FI*IH21;AN]$\G&#2Z,)MS9O(/^QO7HLSY$,Z5 +;#0 
@N1=@:=L!06$PTAQ/>33N9P-HGY3Y WDIF]&B0-2);H\ 
@T".[6)"E3]PZ]+Z^%_QKC+YE"F,E[,I_;3NTW7\ZT?( 
@:C=WY>A4J UG-+T(4"S#EB'%Z-!(XJSS-8S2HWW ^ID 
@%OA!H7@]>\?- MJQ <?!9ZTL\D\EVQ*Q5<Z?#Y.$ODP 
@54NJMD!-9-YIH@T= E=H_HYVTK)-1(APG^$W.5P>&@0 
@#8$L8/!M6))*:KAT.=>3^5\E4K!Q]/T<G%X_H$0*"T\ 
@B^</_:Y:#$=."_OJ0J(2&I,<)+IKHAV^?ZO=%9Y6DB4 
@ IN::Y#@11<5@FD("=\]N9N5QI$*A^=Q^1J]@&1N#.$ 
@G:'X_":QJQKO+C;4I H?"1RRG WEWOJ#/A8VL5?DY$8 
@*42$A5,%:;XG$\RVD2&7VK91SR\9;YF&DT.E]&M*]XT 
@'M-88D6_\5N*S7BW)@'.5?T)J=DJ$@M;B>'!4O-;K&8 
@4><DFW/W UEL;%-M!.WIZU4)/5C$,>T4%W4)7)R^,4T 
@?.+^VHBA6FU%52;Z3$*B2_@^Y7YT<Y%VR8#058/B:/8 
@66N2C\'$+N(>*U0UX9!W<%@",!/>$I'W),8^JL@GZ_$ 
@P2092'TA!A"W^P5K58]I9 4Z[;?E/:(<R3]K<YN+N\  
@0<P/9+"F2?A:HMJ1TF6/&OP_LP@@<:D=NS!+\>UQR#D 
@$:&X=+R":*LQV>LV ,I0=\1!7M"D?(D.';1>0''%@&P 
@;_G^6(T/("^5Q&'TFN)G>POR02$W#J1'*,HZKH< ,S( 
@M8 Z/(G CN[;XA[?YG3L[B:TJ_AIYB:D&5 3=";96J  
@U0G#Z%C1ANS?[(+V=O';AYM!]I?38GU!I\KW&MBV(O8 
@YY*H+4K/PC=!LKU<X0N,Y3:%^["Z!: '=,DYXQ)MO+  
@<Y#&-JD EM\RJ/J1>:UU!\IYHY32I!&@UEQOP2YW,T0 
@Z'QT_'B;]44]9*Q8MI[IFD?#W3MWB7$^GCZF"+"%%3D 
@OJJ]EW5BZ:?\;\_@C<Q/VG^7=V.F@CJ=H\*!KKS<UN0 
@U5'?-R@/:"%6-U[E-*H\18BW&_;NIQ%*4I*26.W!NXT 
@PL5U02'=0]39UY^M+BNO>UKFL*:!?9 X:]OL\@@]T4H 
@/EQ.G@#N1(TL:9+MY8L+\G)?9A4NMA3FLNO(&;( X7@ 
@%+*:/TJ9>$8D+@77SBB3V1AT(DUR%V8Q6CX!@@M8S#, 
@36V<W"(3/$8Z@'6#%;=5 C\0_2+SHG &&0RHB\?9E;$ 
@B]5O'GC<[U-0 N$A<?&%I</<O%PL< L[UP-O7U[X"HP 
@$>JMZ#V(&EGUKZ*G^+KKIMIK#2)KOSQ[XTBIJ<L(3"H 
@6RO!*G>F.V&G7V]'>'W.OJL:<X\"^ -XO1"'-=529CP 
@ Z<Q:;/UT$;BY]%'%0*=SUU&KBDO#>^50>Z*%=P[KP4 
@"1EL34>P3^)>U0A,WAK8OC:]]DFW3C>(WWFYGHIH+LH 
@4<X+@QLN],-C/.J+2L&0QX;"IK2Y&!K@:V4=U%:8W*4 
@_>59I4=L+*34ZQ<V,W:33GJ+S2YIC9O'D\2O20_:G)P 
@ET$*A'_K8E"5I+2%)K%72#SLR3-71,/+.>5)8,RN4&4 
@\VVRQ/RL,MYN$&RA,31E(S [59PZ??&GN=JJ75&\3-, 
@IKC\9&Z#&+84BRBL#CH-*% [GA[>'URSE& :+3+2O"( 
@-?*90=U^Q5\E.8S'TFQW#:M\X=ZP)W.+,&"3TP'@6I< 
@B4\#)ZDJ;^0^9)*6ER<H!4IF+U.7UDK3+%2;8?X9?EX 
@8:]&B09@ST-8UV!!;O0"";<C^UQDDM&!&(]K,!3T^/T 
@"3ST 2\>W5!7V?VPF+-R)F6I:!RSZ*"&8/_E+2 3.F  
@^I>(9R(%G&LL;<9G490LC)RF>+.UTUB] #0X\(GFZH@ 
@,)"!-0I3;!O#L$</)O/74HB&L?X=A.F1&_-]:!9TR;4 
0@]*;K_$! DQ@^4RSEZS4-@  
`pragma protect end_protected
