// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
FIoC7PrK6sLzCVb79+PBWSMASJHMAGV14fZv4DVAEr5zG/Aio172pha1U6zvW566FdrZSEvm3Xhh
xv2tHRAColzOUOg/gNmlN+LJ9NTI9+8ZGVU0+PKlp8c5/LuURR4FbYfaIU4w7WglWotFqvvmq/f9
Q+gTFL7ZZfewKnwootS2r7QNy+Z7zkRh1TILUZif50sEfGRCchEd7BByT9EzH9NTyAsoNZlGpq3c
VM7gu8Nb/BARWyasDIHXA8vcEaUHBbjiC/NYqLCNyLdR+h8YgvmvFGikYocu/NM8G0mMhwbghvk+
GSl7zCYTec9m2F4IhJlIPsUxml1gtTqq/dX2rg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29408)
JBKtTfHLs4h4LC1FUYqzg6XC2y+L7zkH5fuWWBsTN7pvS7B4/j7vijYJPBzVEPTJhGEwEeFwX7RF
iO5sWn3hx/QC43R9ek8BPXp5bIRZmc9scGBke9dlQMxip6F6yyxnbOYX2BljpEmBnlxyz2DajeIP
k3SbTN/0NWU2OVwiZNz7werIwt31kE+/QydqYCqSYbK8wM28WrKCZdovs/AKCEnq2GLXmS5vKlCr
VHCQvanZxEN0jMShEDd12mmg9JYFrJx8O9JBdkahnlcL8Uhj9oZ83m+/qy4TTG+2ynTKQU0xbRA/
O4+yH1xp43eHOaMMDzlG44B4HlHDMwlQH6qmwapwVJIah9B3Yl/ypBzEPXunmJQFC20B4lvCXhMO
JAv831KtyTR7s47skjRRe6OnT9rhbHAqmdV/l5KNQCXqE/YFvDspExHcBTkv8mXzUWQg2HnLk/71
qwZnEa28Nq7JvMSVna3TB/piXlo6G8hhCjogdytOAtXRjG7EQz88AWSBiPtaD1sNd2fllIwT/Vrm
yETslMuWacFsEYD7/txjSjRgY+MJ5Jnk2R6U0Wle5kM+djd9CUNbOgABxXDIHZXmhW0Gy/8jL7vI
eIYUgzfOJQD0808VZIvViGmnDzvRV3jvC0yVwjWzfmGqRkpQVLoWwmq/8Cqv2+e7ysfH+eTP4vI1
Z8PXUi/VZRCdYz7GgUvrN8G99Pe6U6OA19uF+na8EY90c2YSMNsw7Ze0ddCdbj0adK9S3lyH5VWn
uNq3E152K2Qe8jC2tkwwnN+t+q20ljkFkNoA8hZPb6vrKkGqvcKbHxHe02LqS3kfAdiAce1RBZRK
1ytNQbgJv0OyPDQCz6IkP46kSlHjCdAOz++KFL7KJfrikGj4TEiFY6sbjhHZRWBshAu1WrqHtZ2p
t/FWWGqLI3txYN0saMV9MylzFY7P5YHrOHYVGh4gWRIA58jS3y5WOp+2qiY7lHCzUmUXMel5f4tl
lfendhdMv/PtazKuKqqiPAILT2CVR9JJqTBAASt4tYExPTZNWI37oyXO/WSkz7CmsM6JzhKpeXwx
KKgNkTKsMBMlUPryPHvyeM7Hyc75u/QPWuaiqfWjVXFJAc4VRbfYcrrISP9w+xahCTj44roZhwKn
v3AjPwEC7Rl7jA/HuBsAKz+UMsExEa9kD8ZJ/01XXCrXvumPsiXMdLambmi/xYcekQD2b1zYMdXC
sIK9SNQeyU3miaW6K3wCqhuDGESYn7Q1op/XPrpqnS+u5j/lKSD7lwCR6stxnDaOef6JYjdH2kCB
sG1Ew4sl9mrBay6mhXx3XSwfpnQibtJF3s3dzqienAdI7doZcqrwyXBEqSLDOOEhBfuM3Lt3DbZ2
46BKh3TQJXv4sOU+VgdmC4N9qvR5o7MTIryJWC2xyhc8woFP7r4k0fkLAtqHjRvcPVajo6ttVHFf
Uos4DBUE9UIdxNsic0r628hLYElRpTA1poafFhq+An4lZn8B6Ar3ZIuSh7vnqcgYpMzDpXrqm0AB
rvQJa1qcnblg8gkHxAGbx1CL3pyf1fvTdIve746HEqVmbkWLbazajWeilnAo+qhFeaYu0EhMhAeU
NBLApXmaPbqBdMx4wEf2hS2TVgyyeMP5zRrYrpP2zfIvlLfeNYU9oYctpg/ztfNlh/4+dSitUJdf
BXLTRRVv1nVea8yPVt6B6s4Q6byLH3O5wC/wwayxDfM2PwezrFEJgCVm/638yAN76unc2tsiwdXp
xYGR2eVuhQTq+csBE+p2esGeCX+FgZt2qsFzvdRVNVnc70+p8yndqzBsry8s87QMchGtFenZJHtR
bVNIJrPAaCXgmYaGlffnVgxy/hTaeV68BQRAGwIzORh9TSNAQPf5HjdeAUme0KL4/Ixa0lNV4Gli
N99wveRuwvcd/NZFoCmuDaBuTKO6/xHELs8Ih58YFu/C3U93lN7sQ6tu0erae4BVfRpxQxtgS73D
aSrU4WIpoBQQW6e0O3xLf7PqtyAryBAunxIdJrdklJCS3fdLVJ6zWcAOzA6yfCLLPWNjVJk/U0ZZ
zo1qIBn0J34zz2tBoe6ugPNIzyHWp2EJ6EcMR/pgnqlcAzCbuMIRS6QRHgSwvQX8OxjGnWH7TFfN
KAZNGlucEbFWFUhKCXJ6j7t5zco64yO05xHojuncz8nsvU8vzPbHqaBnT1cYlh6pES5A6qcynK0f
conCsNiatgvwwD2tPqMB7VJDLVbBRSanOXgP1v4R7+LAjdny5KGfcboEdSBiMCzFV41h8Vwfj7wT
wLpc7Zq3U3t0wA9Nw2n2tQqUwXiEu5sFNXKOqEFRZ0BPyoxu9TrQ5ge2ksp2bKg4LUACCnw9XRtH
o6NhWW8LSPcws/6ybwb8qytoCAbIwA11XlxdRdxpu5MxQZg73XDMr1hGJPIa+phhWlBMT8L5/Odw
DTcRgZXxFK8yBYJlh6kh1EX5uZ5AW43ro8gKaWaBDwAWAOdQmCMUH4OG8f1p+bY39nwk3T6TB1IB
4Uu6k4r9c7Ty5+KtKUcIvIcrIDBrPCgR6G7xfJTxZaVNyJd6iwVp0MSlnTGpGS9ZjK0S9YVNOStp
TgMB5PiM2/+6JVod9lEc45eU1e/Wav9oE5vFdFzNkUnMNvw6GG1ljwFQc0ribSLLvB397GaPfK4M
lrJQOKGrqhX3e40C98zeovEav/4iyTpnVWGszLK1O1hlTrza63XBZx6jwVHuoT2HbOxxaySCyERB
uu+hyaSkbr5Roj7A2o5YLu96k2Vp9pdCZvRs3VKJY328HUyC8qfCeYFRea43nrxbIqU0FrB3VOmp
/gMSYlDANYPvYbLewOw+1GTivL6dPnBL775r1rC8PSpMJnOBWoYlk2xmX3KtFlPP1VmU0oc4j+gh
mE4a6MO5sG5zn4RUCLF/lPkgYNRHoLhAo/edQMzSMniXzImC3Tai1Spvn4xJ6ZfnEOSq80Yn2dAj
OhWmQDNwTXEYZST9SHgokNVipSVD5m3SaZzSQaYw7wYSoNsd7Q8vgQeNMb+RFET5GsjMD0L8DnH5
aIuTcrQplOdoebfa3RycwgMdayjrgP/rTDHW/vGnw33uVpln6yyIvac+IC2pAEqAXKq0tVXktdkr
SgXsjmIaI/Bsv7IXxssiX8HJndwSyjf+5mFPdbKb+82EJ8ROuqpN6ZHo7c1hCM0OvIAmcNngbCDu
0Gdms2xDsgKZMvavuN6ZuIgED+1u4fvkMjZUDPT8GV1CYfm0Ayh1SqfIHKn278sMfkRqep6WtkW/
lp3gf8ua5dbRisjIf0wPDS2yXq2duU+fRj4ATprOwEMJf94SomKluxaZG6/UxMkO25hCJ+iTz3V/
hW3sQaBlQOmmyL/xUwrNoiVhZie8+bEhye+Yqqyrf+CiZljCtCM8lVX/AeQjibA5naP6jQz/wV1y
9AltMWZ/7bq3tFALLZyatGi9dTZv12NrRrxPsuo1lI00RIQvxdle35tBeN8hZ4Zv3G0ksw50ucDT
OaqYuSwt60FHDeDbFJKFdDSNQlxvMart2pXmETBc1fKadS1osIxbCqDZ4opgDPBIncMt53FjZmfB
M84UhQkK0ghKp1QzQtZcYeXcv6lFrAuJdXx+79wDpmIFQFyy4WeQ9o+1+P6Zi6vlPj7e5tOKa/1D
kUHTt4uhyd+Dlrje11K7eq27EL4FHU52rGHdiJE6EtEIVRhtzmkWNLXuPxfoAIiINKt5nDkfG+VZ
r6/DM+ZNHr8I/MqeBE00sV/stJXseTFbdRQP8frlrubWVFGXN+wm/d2c1/B1E10Xhdi0iLyoyepF
7pXppTAxCj5ktQ6hqL8/PadU5exAiJZPOra7hTVXuUh5t/ycWPGtFRwstyfV147cvi6rwWHsQ3Af
wLGekWzvWdj4+Oz9USl3drAtHndGpL+paK1Khg6pk8nRM9Pj9/CyPKpqqc5vVNWq76Zsn/edrgI7
PvWt7D23aEVs/GYxKKt9nwpIMsV4V/mr77Jse6fKhILIW1CiZAm5k08bZBKztmTlO2qDFyD3pz3+
igZq7Ob504whLKHFTmL89cHwrMCYkmEA+nFk56bnyHY/pTCOzyZLo6RPzS7IgQ+Muw5+3gZeLtDW
2I4RKZPZTKvFpgPaJBiEyo613BYHrGF7Lk39uZvmeXQwDzRulpukIxKVpfdPEunIP4fEhhB+UOjC
0l4WqiALaknsktATJegQMt4vXCRXxoiHyaVYFSfuxcQLXJP0NsfioP7wZ6PMWS/9ihdE7jNY/tl/
ifONj0+3EYGhnTFILnOKcd4GHhuIucMX6c+45sWzzoiw7sdHZ78IWDSvG+kUdzCmWxVsMWD42Zoj
d5sYUIXzYOFvTcbFBo3OEETyt6ZkkMeLMqnfgi1gjZcDHB8uSKUyMFDhiwbZjpfs0ZRK6iofyoR1
lpwl2HDx8HJ63pVXrP05LB4iHEfYdEUDkU1XO8aIF/qW4wPCaYDFGku1Vjrdw0Rw4XZ/xhbiGX7P
+6GAVpcZzcnWanL3J1fmqUSTvFNOdlf/5j/KfAmWPJ5BJ8Xr1keNcNO1sXJe/dTMxu6t6IZs72uT
YX7P9rITC8CisleuSdOPtKFadUYPeLLM16favH64uZhe0qeogEI0KoUf5KrMpMYUXN9/Sx/69Kd0
6KtnXKgZ/cQslAuXkZs6QO+aLS4GA5AUSVeWwy3dm0DL3E1TGvS4TXql7w0Y8NNZKN2JDRPTIVsv
Fag1zS0zS07Q1572AFqWqx194R0ZDcCZS+fpZ139AipT9cfn6KeoyCn5vqTvuyyKIEvM9ShbZZ2G
bfsAh5AVkzQLCu8Mi95KoNRhlOm9/QB+qRHgRDDsm3YhcwJsG2L5e6EDiG7UM86ZNK+GN4dvx4cz
sWIhWuEwvT8g+9NWl0GxE01rzCWHq2l/aGm8TmCzBtjwHp9kCz4pJyl9XV+aUjUWH/dzoGt9gs07
WDGk7zW4Gqrzx7yZib9Av2gPQXq0vA7fMyv31yFzEr1N2Rr8OElEUEfC7bZ82S5kUH1MnWozeo+r
p54E6bzkcsNbIbjXd8ZE37b1QOZM+Kr6qYNfgI3D8p2fJiVBUdwjlQaCZgg32rogFxFMaLtOpHDy
r9/ZYZ8tGWNDTuokgRjxp33N7AetkZam0HxhsByFtaC+tlDJ4bEXyZDKKphDSOJDPIwYDj+5P3lr
IXyVOW831kNgMbBQLXEqEO3m20nxHtXtPug9ZlIeFf9TNZmaFOP3faQw7kPbsxS8UyeZUVF3BrAA
vSmoQlhGOV2ozSR8lbdiFs+k0AxRts6qAuj2vw9kdd8AcJSpA1Ul1QKcic6GBK4tAkPWohwZPerH
uglgYEV1uPypYD3MoXguVC4tMg8sGowXV8sGpxVSREkBNADk9RXF0mTYxNPc4fAFN0ScSf/JWdkW
WXik3RYmAJrE1hw0Oyu5qfkWheXpPqpaNGs92EvwRpHB81AHGxdsVyfQ4a/01obyQT27rG6XtwV8
0kgOQ0Ih3JnGcSD4v8+NhbEcGkwTWQyd04dhovIhdn/0+Shw78EPFQEdyBXWHHK3XFZ2Ca5W/GfU
EqEYxgSaPBZxXGhLoTh9mb0/r+8/xDB/Mrg44DR5M4L0pxYKLvk/L9QaV4ZE3AXvbofx6eyBm60C
dXtAY8iV/4lZzejBBH+aWo99JchnvRwjQx33hL9HAgjr3OdIF2KD/nuQ7SQyV93KBgYp/q2pYN+7
j8v8hPoKPC2TRNkK02CYbyKKV5PFLY3NWfdwebStyeJxaalhLe1Phf9pH3gI+Z5DKSCKlP19Rhc8
2K5uYQhtgh4Y+21iDilH6lq5BbRNxec13Dt60dg4osCl1u8385m9K0Z5h/aRUp37/mTfDIYBpcC4
/MZXVVOk0TzaqVHezuZtyUArRpFITovUyRD1SjOonWGHunYBqeBsA9yadWT2IPZZ5+re3+uQeSZM
Kn+TnA6rzrbNEplFNkSXM7rze2YaQYDybvzGYjH5Nd/mM66CVoefA6L9DIvgdUGGKRkXkZF+uEEz
0Nwr58XVI0oQWn/0OPcVYiahvtFmQqE3cfgv7Hpw0Z3GFWuanmFDR3qQyv0eCfWs5jYSBSnIniS0
IYvD8Ap8/aJ4x292WhOhURJ42XIndJsrT3cq+heiEWcmd208796NarqeEdfERlt1dupoNXfVQS27
+YE4d/aRMi6gcLNOD2HYIBShnOS6AQGDBvMDFt1UepO5eCBe+hig5hMcLhgGbClUL7qMgmaWXT6A
15yslfIxb82Ld9oHN+zoGMa161zchRCyWvw2muhs+BOmazUcCyhbJ4tdsCigLpHzHlfzcR2A0bp1
oM0JjGt27ddtfXzNFCH7HXwCCxa6hbUBTK0O+4VAW40Es1f0oaDO3m+6C0UvTEfLBI4o4NPAsozN
rLkkquKX5O6J+o148/p2UkeW0Vs7pcoEqYOySS1UqkPaoNIMdok44cG2LPhPb+9v8EGSQK7YOOlt
Gav/KxJSc1wtyNwxN1Y8wWhvU8iecPFTPCpnj5NCTU0C9UiLCPsSblJUEtP/8A4Mo8JvLNATKvue
WXLGLRenZLLoqQW+A3jIaa+q2AVScEBJQnJoyke9aB7hH/ns5Tux2IxoB/BgyceTbPI17TwVvFZN
R7NwyA6XHcy0i2AaVg+mBR15E6LPl0ycTnx0akYsDaqsm4FST+2bxUbPb6TOgjNKYKpmEzoyiFYs
kv0J5A8mnY6PoTStSMJEr11ZY3UJItEoVoMuEomO5rvq23n64/IQ2bV2Z8nFt5NI+JBt7srH/i7d
sgzRxbH80yLd2JT6OTSzjdNIzDR/mvEDNAYOJ00B9Gbz7lTHWrJSegPk5E7/QYh5mELkIt/6pBfr
TPCcAlOPkq7pbRHNtYoEOgklIPW/qLs5k/XLNcSuMVmetJaBr19nWHIqUx/KnW4fMJioTVREljRT
G/PIOVTvxUJY6fRBFdgxF9yg0ZNLeeCw+8XevHzswDhKYl/fcrPT/3kbFBxuMaESGDwDsttSn2ss
flCQAVb7OSryC1a5wEaV8FpEuaGGzZRVOLiyga0NUZjfDQzH6fqrxEsUVAKZFCatAOSm0+girFQ2
YmoQ58ZVPPYTxVQdEUCRWoIAeI1eh2gp6gGOOghGHeB8v+m5SXFbxrtWM2DJqtaulA7+eMCeghWZ
SR/PoQp0+0B08qGGR6atmZako+0TpnkK+nwXd4UC/zywavxms+0D8CGHHjUJCXdAUUBcrzcEd7lD
zpA0QiFQFSSg8co9JrYf+gfAPDtjvGL5quh1W9QvYkmdGj+3hC+wQv/54kjlsMt08eCFK2t/AOsZ
V9X4Jb0xaqSnIfPQMfbfapIOQtmAEtaj1NqeJtTAN73Fb7tvFvEGVsEYewOih+uu5ybb1IRjbOaZ
hwXIinCaCqOzxevnGhQk4yJF28YfP+anvD143B1DpS2gEVMP7HVlOSun7GocjLXv00YcFH/4fZdj
YdHoJa6Af3LgHx2aACfWWwuhB7k5mANl+jbjr2HZFeILecrm3E4nbZcBvmswOSaA7zWlKaB55RBt
PzJ5IxGjJUZDmFqWtFckx0b9SXpPxDwWyht176ZE0V1h5IUk3ZMxAerYk8Okw0O5lCLAviAcSQjU
ayXvtlDgUBhFvp5LyBLABYVyIYCbhaP5ymuIxIzicoQEFW7FQB6wCWL3MB8bf7IuUpigt9i0rxmK
x8mz5toyVsWlAKgWTmVRrIp0rDWQ1F8O6rTuzQCT/0CgIaFreyfD8qmV1YGj7cyA/laUMwFIVG5M
u5PD5DF5FKmHPTMS78m9zBWFupSoHHzPEMumVh+aPJctTCfZzcbkB9d9ClKvKwXMM2y2XLC3ik6L
zqXw8aUwp0QzSYe9RP39+wdbsnR7m5S5kDEpr591GYEJ6skBewbwMJI4Pb9wyEqPQ6Xywv4FejUR
c7qCTnfy2oHpyjSyYMmp1ai4L+QkOaAbp+of4/K2egLEeHDjU7A2aJD2I5smu1eF1LscwxqkRzrD
FPphXRJw/J6pgeaQCtpc1UrwoB1mE7VSL26xqb/rwO3n0blIKhnlrjMCh5ceJ1TywT3Ty6Gixb7O
Ig57b98xto1Zm+CWkO+srvZSxu0J5Sb1/0tqd98qe9Jx1/reCV+hzeJj80leV2kSUfwkEGQVHrbv
0cQmXqJR/8JoMj5unm8LlrzPmo6xn58R763BhZn8Q2z91sqBScy6yXytffURr+ZifmNPlQs/EvnE
Lb+qkbbPD1wnS00bUw4B6iMYg2U8UE2zG+Qu7CuB08s6qt6rivYLXSHenKGvWRmaHYkSBoI8IoZ1
MizbiDBsa0rrqXmO0iSE532sBmnfe6vU7ck1rv36KXqt7gMlGubAKNsMw38TMrK493oyVr3Tmm28
eEM3rMYgVFjLEv85oxNg9QEMGE3WL8vfpRj5C/Hi3VitEXkQqdGPZq5+oZXLhYWyNsnRbYBf2GTn
1McYm2u6/3ir5FVNu7AH02OZVxPhBYL58IO6Dq2euTBa3UXtSP2jHKmhwF2m/1zqWi4Pzxn5eXgK
61n37Udu8nSm6ks6qdQtvSoptWTNnC1HS+TriK7uwL0bzHusHklbmSKIx3IbOK5C4scLMKhSilpw
rBXpvpP9EhwAhUrpcEanAsrUUVxbL95Oh2gKihayAXd3puNBGlhrsHAocvRcTD6d0GBhtCpmZOLJ
BvHGNfhPi4Otkdv2QHbqeclPKvVD7bccpyRKXOkxJdKA2lgFtW4RAPQfuemZqK/ltLUzQiiOHv4o
1UrZjdZofoE7QrM+xcEa6yK+DAVvhm2DZCvubuAyaFnC191jx2LiHQUjDA85bWlsU+LM8SGbm8hk
EmNhFz8OSw/LJhOX3S8OAq2uNRO0ZZORszOOA36geVzywUL5gPUvyQJ3hwb7OKOslrl6Dd88tnF9
qEV7n91N9YPRL2xi2WzZBS5YMwdj7IQozr3znCJDh4/uWpNuF1hSBTkY0wuTSq7jjqrSugnwW1j/
o1NdwdjtNaV6S/CFuDBc6X2/PstMu35jFw5sCuJXS7E5r4W4pSCuozczJcLtimhW9eAIgi6AXgLX
wyX7n4SciQbD2uGTf65jB1LdhhdR1mCI4YZhM8AxHg/Xip1+NM8aKa0XdsfDelFWg8LHQWt22hhR
fSvMxQunZ+cVUqFiNdSsreD7xMHvYhib5F+by01HBm2ekcV5Ia2/w9XNJrGOaOcsBRb+9Eiq2udP
nX7MJA2HJlpwxtRqEXOTAjdMLzHXiI30lBfKFFF8nG4sdY9vL2ac1+bujHPEPPVCxZ/DhJ0uYT/o
np6QEkb/RAgisp3viSbXe5WTowQbwdJd67hLFiQI0/9fXkPvDz5CwKACpeuMQuCQSL0l+4WbseEg
upnxhlYVrEQi1e/umawrHvrVLA4IfnN9HKidBTouv0iqa0UhL6T6Ykh6jLVrzVBDZ7wHRchQXgaU
oIZ2lYLnQ1jPZij9AQ1Pyni3Bia9bQaerRFymeXXmDggkIdvnK3kkmIegQKwi1f3sr4fyNGBfH/6
4g0ffWB/ENPWoSg5ppRNzMOzFazdnCKg1+lO4E04eBiq1viioRUdNPGkEA8oZPf4RBcZlwxeenRO
BynXan3NN6L9vlQwdzCbMiGv6FEIfiU1EppuemhvAF86u+UQVVGUWthTJkYYPFevGxITyUl+zFrz
bDKaoeTAJwMPBtHYL5c5glp+Ye72LkQtpib34QdrfvXja6zG3lohwWYWbGmCX0n6C//LIjd1A9wl
Vio6jWZMkYbByMH9WoqUbGx2S1IWYHD7icEmYKqQBf7RdrZq+bzDEA4093rDUlBrnsP9zZZj66TL
jTancByhpu20DmJhc5xbeUAoT06aIAFQc4lRvo8OoArNIcjrSKQrSIzp/SOejWc7XFU1tnk9NmGR
2Mz7Hjj9E7+oGQLC6jiku2KV2uRpWnxrdvAmqPBdlTZAi+LVCvAM3AJRUuGOqKJW7RSqCqV/BCeS
W9M0qhp9c1ja4Uk561DfNq9qfQ8ILoarjGJNRxbuXiDXoeTWKovK745wViKdI6YagsUnz/3cXbzX
UAysp2qMHlK1S7R/10B/F1bgo9o37vWWJwts8Hr37PoTAcGI8/4cXIZkIC6o3dm8qN6yiHUPrmQ1
W/gj8aQMcT0WPdX2Ezhg8qOlX2nYYSoXPPj1iogODCMg2d4DhFwpP7TeTAMBQYWXLSxbYdZHwOR2
Suoy79TvufmNm28anWUAehJwXc4jY1mr1NSHNAsp6TcGYjfI30uD/83B4rAmBUSiC06TtV6UYbdS
PNmgYAHDsACRw0+2f9GGNLz5l2B1TULbPoQ91hQFL4HFgEXt2TFngAM/4S+35JAwqsDBDY2KBsDP
Ag1EkJS5Buh10M4+WmvyfLd/1ogjsJcHLAG39WP5NDntz6Gy1o5IJx8U7d1a3pCQuTrAohvsNsNr
fGywJpiAxQtMI9LtljIaAtkNeVxP0JYkf5v79GLnajqyxU+E+dFpsjzY7B0P0wfaxdTfhNw9yxVp
hjCn+gIPnK1RQeH4nlr8GfryB94q36gECnW1UGmB0kVUN3jh+BkwWupJeq4y7zaneJW6HP+l7x5F
BexkTynTLYGHTbJkPy/8+93QL35DbZT4FZZuqEbimxaZt3rrjTSm5GE1K2UGB3QgvlnQLNKdsgfp
4dUCQ6YDB4gdRz/ff2gnZvBhWONSpIxwjMiRMcaY4qiCbb4t7v7Q5zftTsoKpFJfAIGQ3AvIkt3A
N9vaELV0oydKzHPdwFuJ2wL6axmNUUU8wb9sPMqFDUXGywBHpv/gd8G/w1s5vUJ82ZWsiTQ/NBTW
EdoSOMSOtJmSv30XRbgLoz2gTvv/yk2ndKGhJPrsqVQAySZRqLi6QGKDEYIfySISC6LlVghGe/yW
dq0BZoaL+4ykpt3QJ3dQbtqaEIYxbyfk6kMsgPlc6Iu5Usvr9uxG7auwuZNBxUIwSTsC1QXKcgLj
FJUUcx5cvPjv6Qe03G1XWPUcda2ZJPZzYtc/UwccyT9PloHQqtkUrgRnkIldlMCnEReGCaU2cXvt
ZloibWt7zPto3sBLhmkN1uas4JjVRgZzdJAjH5NZtF1zVPzpSuoQPv6DxJyvQHUW0V9K8mDvG2ap
JWSYXnJg9UP+pECdJ7FwnsX+IDWJN7ZY3k3upuePRgB0nvc3JDBVRDSDK0zoPAFgvIv2yV3Vwt4b
+K5rrpdO2r7fbHp4bdl52zx+zQH/sHwHm5AMk+4UKL3VRUSZ1Qgh9cJ89708LPPMNNnvNogJXDzU
T/N5Hz876VMdmbP3xW6d5Hi6gsH20hEdj4MM08Ni/fX4wKxsAAACgCqDrrShotSlpGwbVSVmbH/H
s05pLwWo2lTBHoUTFOUrHGTlDpURfFJJ/zw1QE2MZuNfPFExDxUxxvW7197ndgtMOxpEq7neCGwo
I8qpclVFwCAIvBeTH7Uc3HUhrdAcs7X+MuELQDK4zGk9NVvKNTXWRAhbUVorB9gB8HQzo2I8FyLp
qmFliDNHH23hkLFSN2t4A68QTqhxjl9co6c8X4D9hLPMdtZNRRiDpVOAWQbNjlEnVqv74Ba+dDvp
zp9obn0aOSfdZE6o/qH8l7++/jNO/JT8tnfUtXpD0/Ytc/Ag1e5b6JxNleySh+cqDB2E5/g/EVWO
LcBkVNquI98QimFAHKC/2ZiL5i2mjJka1Jfx1m59UVtlOSPC4jFA0mt/D1Dh5vYEwU2PKdUjZw0o
q+yC4Vm38VAkIl6pkfq22qonI3J9wQLEI8o4M12ecT7qCtIzAtZmhHBStrDut3V2o03J5DejVijv
Ne+zr/kRyYvAmANzg85Li4vrl87S+l5hGMnYoL/0iThaj+O++rpILzKuGi8PvyBrExu1iBw6CWWz
DtcLC3MVbXuztoMncyqqvdSdhXdFZf9S/ZosY83FncrmkF38nhSwPATGsoyDn9x275S1CNDhu/K/
9cqUUSg6oH0+En6rDZCoWNvgZUehL2xMFAv4k3cmkfQHwc57z0MHKmwb9w6fhnI/VJQZJgERwXVa
XrobTMQOdeBuGSpMweYs30Q+Vil/3QXmmk8stK70UCFIFvy9j+4waKIlcHH+jJJJ6fWe/73n3oEH
ahYITKUqBNbILOxQE7LMY2vIlqCMEisqC/zWyDNer5s5OFAZndNaIAwBFGi3RuXsb0tnl+Vha33s
yFTtcXP+KhpdBPz+0wQ1KLht6m/jeEs73yH3kxBFIPvGVtViYYL6GxDOZ4phJ8eWSiVx18hvS3Po
442ww8OevcGZkvS+6WparhAyEWpHvMkiWasX3m3siHVGjOwOFhmdGfEH5DwAIq/NTYc1PoP8o0I1
6UVzsxHZluvOY+JTniXUwlmlOXAr3JFsGG9Qu6Hj/DGwU5sswIY3kQk/tIxiiVd5XSxyM9fz/Q63
ikJn+aFZnI8Nud+YhaKCaOTLvmdWvZm4mD29FkvLbpz/dieiZRElgYcuv5GHBeuCsy30xEumrvi5
VEyBBy2fVLUR6nexBYbH6EHWbXg6Zin6CILHiuPhw5kKD6MXxtVtw2cBhTSbX+cYDNiRnlkrO6x8
k1stTkLdndcIHXiRc3Rys680+NTRMkIwSh/LsgjTi/wOUlOSYs6QkBSVaT77rFkxPDBzOGYTuW+/
c6IQOw+9fMVPz0uy9szcrKR9BcQElTDnv9tEkp6LCcbBDl6Hbxo7ia0vGq/FXj9XIhh1CI8WSd3Q
O8oVAkTFm1TWn2fSjdXfsEBBX+ZyoV7+h1CxwSDwUZ+gzc8bgsmSmHAmk9nJCQSoYAoCo0VJUx/N
F3AEJpccPAhRBBjIT4d/KX0SQpqB1SBuTr+Zobzqz9raiTTRJWmpKc89j8IPwUIEXo0E5YNSXxQM
nesJdIL3rbNoL+oehggrcmETib4Zlbb9tldkuU8nfA1yZaJQu7NynaTboROWzeb/OELCSBZsXFs3
kB4EX3A61bTIca/C7CoNf6wCkZgzKBeuQQESrfxKj0MVH+4IrjKGKpBmBjen3a3r+yaOnIu51sd/
S8blNeuo9OfSGR0rYqHe8TRNl8uf4u/Gtad7mpoQ+h5oQKJKcZfxQaLf4lJnF+nUWQk379L2dx3D
rgRVTNPh76cea1kfTiKa8IDlIGoKluObk/EJSBFeJhVZmpgB5bXEYBhp78/GxZPO/GHvPX24EZ0l
RijSxKR5l2m7Xm4hFjCVCQPRdwlRiWLJMuRySuL9YKWfVs4HZ4UKIvoDIeb68sz1GdIJLrA4llE0
IQbdB4+dl4wRTKB1QsxFfwkJNiSgiY0lkWZf46kZG02XLqaxSMJyor6VJO7ePM47PpWME4MNd/uw
4W5PMYFNqrWvwl3u/0WDLeADhFDTIrbU9JJTBhVz4K4ybufrMzyx06KLAU+6Zin7jDu2I0ldc66t
PFZbv4fFbmNsyE3G7iLz3hSfrB09L1AQNZtV4nuJ5JGZurJQ2L6VDHUn7uLvNKtbJBEC3zkbFLrR
U/nooJ8ni3bS974caRtkenIQee1VaTcVH0uz0+goALVEv5M03qI1UAw8v0jY0RaiKMnqurNWnmn6
2dsluQkbX0AdHMnq7gR5+3NPDWII+J1/nu5EKZGTgpoFLpsJ70H9ekv4WJTiTsuTy7gPZ88Jbzo+
K1JAvs75LaU3yHOSgkQuqHzsJnNQYey7v6AfNkk9pnKgdL7p5aSXKELLzTfHYaTkjQDDzv6LCPZs
SixZkpN7CvNnflp9vUJ2LQXFlsTD9FbL3YjcHLA+9I8/eXvW2AcS4ZCxkmpz7V6Wt4/b52YZTDU3
YG0zmAA1TbrFz32nBfRIdJPQPJ4TTjRrUrH731dxXJjmMGfySLSiW0XX8ZKERcYNPxeVtyXc+/lY
LJFPXmDwsv1nVxCLfzpt0AF+X/VS5Fw04iZChpjIdHE/9fiIr6APzdYz6VHcXv/nOUMpI43G0UPo
hlReI6sMucjGTXc8JUDRHglyftXAhlCSEtykxCrpKQDVRr2/+01TJVmFxY3Qekx0oa1rGxPE2DjD
Uu3a95/laofDiz/BaCLDvxcGD2zArQ+yOG/DLRrbLGmQn0QHWeeBvOqVWdGigC9r6w5fuW5eYaBa
o56P+T6WymITavutDvonJB3g746lDbUSu8Ino4VLob5ybHrQ9ZrZ6LeSArEL/jI466anH+MogjQf
vq/tKqSd72taWwQxA+rwXPNiSaDVdaG9mTGyFGg39fPlC2W3uCzgy9VM8j0SSvqPddfz/OGGX/Kt
qx+YVJcqeWn6Jl58FWZBzbiQRc5DVqwlshlQFDGruVn0Ogx4ptzxj8r9bUqTLQCZAjinIyNxoQ6E
4QEe0AyMDRoxAHHFEn31P5sxMEMqYNZcqNVb+eb7pURztYpNzBXhyB39ko57XnKiQFSUBCc7y9zV
pjVgvApvg6ShrNDfe2vtZl9U4jrWq85xQv4mWL93BWYP255H9vS/byixR7W7iC7w5dhtd3rZFwM8
wJRMhW/z50SsF5XuvoUxf7Lba9I9tn8ry3az+GX0TAJrZD/3WSrCL4sXnIsyax+4XYaa9mdymxIA
hoXl2ItgLGf4e6g4RFlMi0tLG9h9VqacREx1C/18Rh1V+r7onUFzvI7UZWWcJpkLr6rHT+ZXYAzq
T+YmvsnV7SF+okZ1wP0JW369Qi8Dk5UQVuM4QovmeM5Xdld7VeoCIhGO/GCRYOUhOFhiHEZosy3/
svEmue2FsgZc6QrAH8FAGGD5DvKCdMEe/zJlNdoBjpqa3QfP8IwcVvC2WKnk6DIVG78aonXxRpp7
apHrkfebXt0g2/SBy9z8z/1MsLiRdfIGkFPZ6vXkQAZzp/7tRiqAT5MrPS+t3ElnKfr23CoVwH6d
VaxdNbOurCaSxWS03ZD2cCpa+uose26HzB+WEsGWglmeAq75A8eHIKSibOk5yBOjOXDw255gU5eV
WUiVKvD3fyYcuXC7zC5jf8EZveW6qOY+HYVa41A7Pi7uMZaxm/njenQokHSNEUIzE++agwo2Q7lH
1VosXa3rcs/RLcAVgfj8X/US6QYdIGfg9NZCjTsgACbMvMdHUtdqvAg36KNSKbwSL3aDNviMDeg0
l0Bk4QraleEHyAc73MqukHHN9+XzcTZHyPEglNmnS1cnVwBYMdlXfILjAe8hBjYhC+4GxK+toOZe
DcWhHTjfgFvAKe45owTRQ/97/4agxHeTLlMbz0c6Gxsm6LLp56lAZThQYo50LGRHIpmGdXUUYjVN
EKJlES1cdKhrTR+c6dXCyPwzvltnSs384pSjugzXWJCZ3pkTy3hOxXKCkQsrT1gmX3rZ5IftIvc8
DzMyE0aKnCQsGXVWPxNnvb8n5dWewkQW0z0g2ewRmrmpUiM3gGW/nFOBqHcfkQU85NaoCUNC3pNY
36T01SY49qSP0nKcXloXLFYBYo/ofmKOswKh3zgvd0YZ/4waDAPJJKJeOxOi0yDCLvJ/mpHmYlNa
iwkQ9icIYR0s8OiHiFZljnHVut3bhWXDG8PMBb6t8JytLEPbsSMmL+aVl5ysNxW46GKYY5qzW6Ef
rsJDLviEdZTnrqWlFi01XYe8mzvpDBD+7RE1bYg5kTdhAvEDLaNOPg/btq9K+LtTyxTInfHvvRd0
NTZqJ2/9FJy4AkwXm15cCm6pBggaKdXVu6eMRg4wrF/jDV3E+qg1K6i930CYK+LarsSjLXPqyIVn
PQS6rYy1dELATl9zePxXjQTk7D2dyXFyPyGbuUHOl7q9xIuZukUw9ukF35dwxWoOkZarwwkf5MtN
+9wfy3SOWUOPUiRau95NMXfQllhLbfj3f2ymtugaqiP86YWc/l7XfjGvg7KmqotRwa8Q8PfJqMKW
UB1D4Z4Q/1Iqb1n3N0eu8KNv4r64GQm3O2TBsNJf/NUhzS7JUqtrJoJXY9Px5zeyPJJztmzdTPPx
MJH8xVjYUbkfWnMWD510pAxX4XrJ3+5VvTkaCKxwq7dZ9s/JZJOTCtKwIJ15uLCcqVPTbx4JvKMm
9kMhy6uFfn1D+GnTEaD/rQ+BvLkkjRr0bcwQ24FiAp+f02ZJu4zKc/Vucg7kLcz4VHZX+Lf2jiA7
R8vo82+7qYrhHZDHtQpR1LLoaddroB6qhX/+HcqP3PsWdhtYoBFf3bawC8fIs2FlOKnXB12o1Tlk
j0b1sWvIxxyp3hXzyWJ5zvDcbt7YCchlTJkRr/VpDVpw9jFCdzgk3guJFvOG5PD/Z7rZKluFqmLP
JQwtX/mlCIPJ9nQiMWecFc8WrEkWLePGhR5fA6XsdDUlYJSSgAyx3gfZk2FNj27lAu/CTfxRYf/l
YaRe1+y/2GARmgC1+egLZhCsVT4YnC21SBMBOJzfYKZ8n1lf/gNgEnQghn7D00RpG4Nwgrq0587l
XJ7YzKgCDK/U8pLFK73uuI4dFiKJdup4YJQhJn07+JWEEpdmXn48h0Hkestjtrru4B6N7hCcGLtM
9jC74sGHT9/eM8feuWEhLxAKMS4upohwhhYNzMsg11lRCmvob1tSfmqz/gT6HQZTql+E0nKt96LE
e8SJ22eBaNwvJa5N4rDUoT9wlxivJ1YSwO1ZmTxpGtIKMgwO74TJA+1iMdpHAIyAUmc8g+BaAdS0
Ch/VZYaj80m7bW4jioO6uDAouXDwHpuiHTGHmHp5J+AYsIUb6xYH8/GRPkE/RIWQUXll2frXSAfg
pklNMvnAF73BOlV9HSOtbg0gs0cB8LLpUeuAY5I90i9mzZ/EScW1s+T+bopYTOIPiFeELDCPDaYE
FrE0U51znsQkRbocF7tGsDEipas0F0TQj/7QAhJSEedus1jmrwk0G+F8MVzRWcxbjPioh9eGelk9
D8neB1N4KzVQy+yY6Hb/Mkw4U1pUR5XjcsMb6YgCQRc5u+9bV+8IoyeV/PWnudGiY6H+jlheqrn/
GBxOAReTCY5eWboZXEkMNTKp7rR48Vh4qD4Bmggf92GpMe2QN5ayspNAUqHi1qmZGBKYn69qqQgz
bBvNl/6PF/ICB5lvN5ioPpYDErhJTU8n3x3Gf3mAYcwc/PSVXH8kZMoCRwxdCJ1sUKTU9wcCkZu/
BF6rvCohg9qhcGWMjyRsBpnS5u0jZH224LMgUvtavUHJTpDTgay1eGbtxgPc0E1nvJ5Z5gU06Bh6
nx/KHpMohgF8SZFDl/FWJ39zPF0DEPRWgKpqjEszXjKk0XQ2JCMpj7YTSQ/gEB+0agRpJmj7XSXc
4Qr5itmZ04mpyjx+qIqu6RZ/MY1nyvAMpFXrv3GV/9W6v3DsgJ2rANBY4njKN/muxk6tXWtB3Mtn
9dYtCzL2DQ8hXfguxJD6Er5BWrrWmIM3ch+lKtqmPlKTsJZeMorq1uVTRyEukncpV8JJOizw209S
AXEE6yJVarA8P89lUiOXK2RRGrwbGals5D6WDL0XNvPJQXx05IJhhO3cO0CXy5uvL+xxD4iD30xz
5D+vRdfelyKv/PoNzwRrpQV77xUiYhxRdoSMmowGGBlXOLBOsv63IAEF0BU1E326QQhLenzs/+GS
AG2aIu/uInVht0IQPN3zcExC8WfpfCj/EdmvPLP7+ivszpaJ6acs+JjMMxH7X8IMhS4oOVmFJKDV
WhPUip164svzvPVUqlHB0PsPvVr7VkeJ3vrjeuhVneBzUKG1e6R2vMyhUmFyN7dHug/WpKzzQJDH
mzYpuCDykj+BuboHJi6We0PogXvQdcXeeAlr5FBgKDi5TOaO0ZztBHLGGhEauNBxlfpBtl/mENSP
o5lO7nrTv3+4/o+4Do9V6pPHiG8wgx1/EdoA2bbMgMJvqlULTiTln9El6LWH0eLHZCQQ4oBt2Tji
PfOkDOXUO83gXUqW025phyAN3s4TaphfOd9O/SJAaVGVkBtSQzYwXCO5z9y9Dx3H7dSMpA/5ZTQX
LChkOpiIP7TkaCDH5cIISXpV8QxmIB2ZsnxtTZ9aYPw2SK0fbWjOE31VTG0GWdl4Cx6QqNoF9cT6
g/fr9Aes9coud5vbBXOVI6bJEKv6Lex1zkv2mZURwVWduFAb5f7cKvRwtphbj4rcI8H7zj/b84A5
7URw5f3+GngSlsVZaEAdavnJPwb/TrKz46yC0fnmXBU+oaFU6GJckTRW/SwfEzD00/BrgpPUVkWt
Px46gV7S01BJkFj+4cmEtzXZKkle/eNOMty83aT6du8RQ4NuKseURLMyG/qaXaMC9BVetJ1YXUJn
jztmqEc8k7Oi4yidFgwDwK18g3BLr+yxSuwLcfRkosKJL0DxG99bPT29UMjuSWMxtz4e0aiA+sME
Pzffcxie2egk+fwSFZnpRsxbrUTuIyTmp4XdHSJcE9SsgLI3NYcadMsAqK49KoaCRxDcZDGf158J
W+h2qNSB/6K+Ni8KEhofmEN9/CkUM2iu4tOR+ZsHb/DUAPR2DmPcj1Jq+GcHDnU267wW/GVxPz29
i292KLi+SPdBQwz2vIClPDeCEsIR/ArxQzkjmH/KbrPLcQo0eFDwYNQBk2bQgEVAJF/ybAmv0TgU
wT+hzBf6uHHF/Gg5us1dzGJu1jTMfnilr4bo5Hh4vi5iRbL8CwKkIUMvkPCQIeUCXe8FAcw3c5Cv
kFbgd0eC4IsS7IZCqoWoKZBDrlDsaGvooqqYHUfXmxBKkicFQ+9oceCQf5MoUaiOA0mKProcVsjX
CMrf5Ho43wP7lQqY2hJr2CvbOqJX2vIMd6SQLppq4Mw0Nu0whjICp8z0G7YSaiS3zqob4FlmAjFh
RMCyF89GqL+ILjbq96o33DHhX2MYUlmODGdB+c+L+CYfab1WuLa/oHXw3ecGYIT2nMHSDKj19wgx
CI9VsNoGegJcgKzbeUSBt/w/x1icxnx0FrbleBNwyNr7XCPSMTulM28BBDXV+LLB7adLi39N6NCe
of7E39KQiG298oBkvY+nK77DuBOBkUqOP6b69QoiojWz3E/DsfEzi8x234KM/muU9AoaaYx/IdHH
Qvf/nU3r7+uc+xc9LdxPDSACTaFy5Edlggh7y0Dx1g6mrX7Ic7XcOPxeiDTlZZEK/jzqY81Lhxyz
xYgK7ZDHeHqaHzOBR5tn7C/fHmzS8wxWxK6w3arGrBkBDWmA0aVLtWtoH6F6LvDlC7Hw1jkKHSNh
8wuceMSty6yiw2dZ6mdnfifKMckJmgIgCwmbGuNMF+UUAA+JSK1isyq8v1HZu01iSxOdZbli8EX2
+qWdrBMxkX3DDZHS9THnYDn3Oq0IwSQfQ2fO9mkHaNwxGgpokNvhY8tJ1qH7K/nBJXsyuMIi63SW
57itt5yw+tTdv/QrIBUIuX02EmCsf+8t0kpEUgkYdORd7HAB2uak2KaGVBbfNTE5D6zxerlkYb0p
hNa/qJ4DbjOpHtjawX/tAlRbAtm0l32bETsx8Ipwqvj5O62KRdj3FjIbLbcxEKqKbaV3xCCds+Dr
OfGZMDXFTczklkuycyX8yi50CrTamYasUpHUieMZo4gjZ05QDu23GRFcpjn84qklSpSxDn9eE6Cv
Ja5qlu4AAzaMJAM5EjcDkw56SEd2G9T2l+R5xOjNH7/7u1ZoyUaUJ1djwbIi2azPyClPXidhutc9
HyhE1XTi0BbF4feERD2zFNhkvw/cWbLT0b8PejgyWoleyFGI1FrTqGa53yZOCHggrvMSzeKTnmTT
lKyMUVyIrg3uLi5q8iKFHc1ZQkrohhG6MMN5YMhGFyTfp8z8YUGffZFk4jRomx8Ote6fDpLaZxPL
7yDCXUYk1bh74WkfAP365uxTEvtGYvEpk/td48uGZc2H1qh8dobIvuTVBqYVEX7+4o17TX8zbfGE
17o287tln0iKJ0F+E2oyAmacGS74gmlm8xiDuEMXMvcPGHpNiEmhu5jPRp/Ap+IoG2BhUoUV+VcI
fUT1MtxX/i+6wT1a/HFMFd/EkPKGYpWKieHH1S7lwex5E2gactgmKXBn2ypsPEo2+qPzAoalvdcP
E20Sd3tuGOSyUp5/Ksom/O98U7ZObe1Fh8/+KQ76/LIK/3PJ3kgqFJ9z75RNgWuUgiAGGyrmyaNp
kDBiE04hJf8p1ueO3z+4qjt8QW2UgwNtehn/+0NkRFvzc6evY6rXoJgjPvuW9jPiqDVSNXq/WgPc
9i1xP+ZhsjA0vgRa1hELhRXKUgb+3J3pf23z/hjMq286EYyBGnXE0Kx/6lU+jlr5wz/NISboy6oo
ptwTSXBsFkksC2IDHh4VJO+JLKJHgLPNIvQhHEYEqMNMcIWv9ZAkgMhVrytDvzaMH4cY7gdYDoaT
eTBXBiZ120ZcCY05PXqmlQ5UfYj4nN3+NPSsTcTH8i+HF9Fagrw8OKgD1ba+vVbdZgY80CBJfxg3
8IJ4w9VG9XeZyehsI+PskZpqSQWP52fLk8rL8S+S9GUa22na3RqbaUSZKE30rSmzSc+NuwRb43hn
uoLpAP8JOVX8z74n9frYluVfUpbQIexXpMJiREEVPkDWslBEzbycwwrvxOi1F8kCACmmH5vdmVnj
DP42K/3v1YxqaGq6gKPIwVgLzlYUAfkp/rr699HfdPDGFvfI2v9mKcuWn6ztkLvcTlQo9H6f9ZCg
zuNEJQFG8D4H6nCkNubQKJN43E7lK6ioSPOwL+DJq7X631jPu//UIMG0NIU88U2EAaTMuq2FIioj
GzIhQ0b7Or9JKaRyFkZBlxBXXJgEWL9g7U58wykFU85jc+UaeFQ6tVz2+t6fBRYwCSmjfJ3O8cGK
GT9k1wBvtFVeQ538fcmh5HDGSbnUuzcf3ctHOUQVE6bmpt3yD3TEvfDyUgvzO84zHPXNx5HGiRuv
GZ7qgsbGqrYQyqgS0cSv39hqBjQ9DNk+02v3zsrz1XayjCRd2pxlnHuuqJdQjjZjFSEl6wBzlufY
GNQdR6nGtkyd34OiRBEbUBbScRMSzlJxpqZGralrKeRTeJxMI6qJFnb7ocDoi+zs3qJH2dEOXZuy
fCudGLEeZ1SrEZdxsVxwoz3jl2ATCYtOUPM8H0D34l+8yxlvbWEi6WQX167vDAvoWz6sXPgxpMVr
nEHk0B1y7PH1T8OWYjdxCiTIGrdv3El8PlbcnjegKnLGdwbRwH6e5+PHSuPuSy/ew8auVwm9rCy7
Gbh4uS2FbXO8iDsRX7K+4nUMFuDEyugTFZrCvz2dhOznxLJ2IzB9nmlotB/NXUnI644MaNWsvl9m
yoQlmZuEZ3BByRvgCjIKbDZL1lyZlDhLIZVb2V1G3BpRomhDBs/0c01OumAHak45VW63NSrMGV12
g8sv1mqwpa25jGmeOaY66GY0e7po4elom4WyuE58RdofXKUMyAehFiunBEBOAYDVUMr9JkQVNelf
o4mi+kdqGqGeUgTNKvZvM/gwYGtpDrjY8J0tdNbJ16938pwfYq1NCY9TEDTk7HjUwq/kf9n5ZjD6
MNC3Rs2tGlrOb4RZ5HUhZhke5eU4Cp7zHQ1HZKI3tYvCmI/egHZOps438UMmt3GdUwLxImAMUQTE
+olEecRJxeqGhNQ7msyekyt/UJBWe1ySvWlS5ZS6tpNo4AIv2zN2XJgz7Ik4BUNy5brX1yRDERmw
NqZwj0CY53UsZ3DPawZDKusLkSdx3zq5QefQ5SqaH2IbtChFBAL/EZIzzXv1Pdw1bl8zIJPvdTcs
TR7htI0pFcrFkhmc1daf2re+L4X2Ho7dk0F7YNc5JZUnjGzwsyw+s+EaVFeDd40YEoUsq4zMgFA7
rcG/ZT+eMWni0+Zc6p30DrTvZvkzdgCFgLwfz11lFvqA4SXdF+eXhfMUjOi1mYHGgUHHE19eruFo
aVD73FRLhQo/wOFZM1zhpdoKf6dQYijZ2ig0VCYAM2apZI60qVEQUyOa5gt7e7bVYcdOtt/x5RC5
vFeH66o/WkxuHbiksE7YBPaSbs886uyTddoEMxg1j1rca3IXgYOXg3uf6nWoKSvpcdJKGI23QzN/
LWL4rzmyUuEnLedKCczfvFyLFFyQJw+VyviviCOAL2ybYSP+TRt5MQjzym+9GWWa3i4U/63cOrJN
tMa+Q8TdOyh6E3KIVAo5gjIsC/MTebzvQDA42u7syX7FKkICbGBzz2kjyTRcjAHrC1RSvh9REPU9
j9ZYB0Kg3y0Zc06yXAmV3r4ihfqWm2PU5qmeRO1KiJne5rm9Ay0USLthJyAuuaM6H54YmuU8H0os
b8PtwmvZ/3fG5ruyyBKy9e1RpVtdw4RyxgWXugxHn+iD83V25DUasS0uURtncUmAeD7aBMunqI1z
4OK/z8sl4Rzs+JjlqLaaYThtNba+4oYt4HDbTJAyi5Fl/lFL7BfnBlt+eQtK/ZHkHNLOXm9oa23I
IV8uYT0DCD5vZw94LuoV4k6/JbGOW9uJgnCglp757I0HQH8K8WbKwXKRXvOgWmRW65beXRm+tX2p
L+BgMG4ZaKig3q5UyTpW9Mq/PGlqr2VvSlLQjDZUjjfXxQM86atFXUL5VrN1knsONsQaek61s1fB
ARebgD9ZGZQN1ijV3Vchcixz97gP+EcIklaQgtBRnoJUEdBmyzZRFM9pL3J3VPYkJl5woldG0QR6
BzrW5ZPI9qf9ekfO7zRgqemlAgiXLfR35Hani2Ea05Z5wkPez2KKpQIYDN4GD0rBdzRlxOV7pDap
KZqProZANhTPax6F4dOZU8NJsjaOtEHhrfDs8AzNYppu8wjELjW9sZAuxsPR9blCakB01yuzR5kZ
AO803fAEfgwDUalF1ArJpPvkQco3VEmjecF2ZEo1qMUiG6ZDPu9zZMoz5Oz/zBGmk+BiM70aHr7r
pRH/wVI1I4B5LwTrqYku0TqH7UssP+MvMPd4ZoLZVqIKZEBiyQozNhVTSgHaI5n88LBpSwjjXNgh
Kt0Da3kAkRIiWhp/3pyHdq1FEThqvbG9uhf+rf/JFyGksozwOBc4ftqOfpoS2Pd5ur6+8kMYG40w
L808MzWLXFqqdaN5I4aTl02RkjyaFEg8sQu58v/GuZBn4V6APKdO34+RMt2CqLvvz6NKF0K11MyE
t6weQ99WENSmOy3Vmp+y+kO2Xiz+rAbypUl0YywSzQLjY6ui+eRK00d28PpnB+NV/r0APtnOhMiJ
vuvHyyX+EVXk9MFHJwDjURn3IWaTniu8Tyfknewv1GnxNKfbrY+dK41Awdz0PEYM+N+qPbOnO12j
1YnnHQCDS1OUC4wri6jhLVIECW6bWNhrMh2GsCE15V0BL8qGS8UL8XAJPCH3Yh86EksOKf9C3Ygx
eGKpOI0th9rZiljbJpkHPj53yo35D6489Gu63FZZPS6pKQYPuYwn9WeQftnZjKj+yZWos9EI0EgI
Kbt808MIknubtDLb7Df3OHr5jtOqYgGeZjMoH+di6lbza6ggLe+oHnhbD/RNBmcz3gYzUqpisEr0
fJA4hHQQGwqZYSdDhyrJuzqFAgdPDVMFet8sLYRQ32V//bQuPXx9I3yqrRU7nD2f0NZJqqYtoBDh
OR3Ydj2jgOyamS2IQWcdh8u1t3qt8Zs9q8xterys5TtSCItce7NRvMVTztV9U6wUi24EX3+2wzbQ
3sEYU0Y603y0AeyXL4wnkkM8HgDhv6l137bKWhuKU+EH3k2DRgBEC9uAzk3+Ez4JnbZ8lzn1q1za
4VPMvwFOVHaRX2laGziGzI/EZ2yxufzrqDwDLsur5SOzY+Qk8FRWvurobFoKDdf6ESrOYcU+ocXW
NyWDx55ptbbVcv9oRVfu/5gCqg7KsnHZk1odRLMex6UeGTwLIlq0PGpa3VaE/J+Qr8/0GEAwQq/6
6JDbTt2yu/h2te0dlBTKiMYbk7mKJ1zeaTiAfiEMQYzb2DObuHtBfp7FhDSeWHzCiOYrba9uuMfU
DhhANaSF08hnTj5YUDwUm7UKsaMFTZVfC6aG8NG+H20/NxziJzodDmrbAS1+q4d3ycd/ZevT726u
QAvFP1m0Pu/gLYDKvgBdRz81Ou/+PO7670W7jJizg7sng6SQyy1HdXNd3UmrX5p3Q8dPcmH8x5Pi
z8Qt7uigRh/+kLQ8uaLKawo7ZeEmSmNL0zOvN8/mXlM4rySJ49kdiTvvA0yf6B6lejY9NV2phpEv
SuTyPFXt6SybnL2isFZAZULze6cqtCJEFPfb+R23S67RvLA6wlSP3xZ3xsgslp4yqSCGVbc8BUcf
GQc19IRpt1qoWMoESKQzkdQyOSUnFFB+uTcEdaiadn4nEsglMz6aBknNbqSZNIAukE4uOuXIuB1C
sA5CGlNnXTnqaa+g1kKB7i54d3zeH0tcDiop6kVm1ckdYRzC+hqvaYZMwUpxP5rGKQfhk+Px4yTD
yIxjUoGfd2k/zHt21h8y4jLkiLPrSCwAW0XNNTJ+r0MixMJFOXIgsL3jrQkCdt6ch5m1Rq0pnx7i
klr4GXnd91VrAj6y5Bnkh3xWQj1GT0uz6XKZa2pLv7MS3aFLjZeJzp7sAJECKoyKuwiG79UrUPot
FMdgUOXNVgonOtaD9y9C4d5lr8urvbcqx5KFCC23Sau5cy2dc9IByucWI32zASyT/px/cguRrb8n
pSDFzwa+NqnCIstZ+yfq2uIMLrpTg9Ba9dczBevNYRQptwcAjDphGikVMq5UFS575R1Mv2cBdu+r
Jtutc0LyVB0kkfMrRaPIDurCGnBjHbuvCF/EudlqUAyQvdy7GWnFATI0qdpTTD/say63A8Zk5vbS
2ZiWvcScD5W4MI58NFw7nxLaq3WIoJkxN4qSyxIxvfJSPdb9tS/dPp+cEZo0TMZPlqVyJCjlvCcq
UUhMTlEjS+y57ihJtSHGtNKNH40ao9m7zsQM6Ro9eJU6a9I20nmlig2oB9VzkaOqppqjKGTA2HJP
OUHD41B5ZDqwqMyY5DQxz4NENhHxdXGh9uI8Wj77pFaf7iCj88EP/7DTrxU2gcQr4dlMXIKkKh3+
0tRNCdRzOMesdYhPHykSfj6g4K05X3rnuN1Q1Rdl/7C3aosvwSlh75CMVdqNBOI+wwhlxtSrbgqx
/20ptrK/ccT+PVG1T5keQSdJNZoG+7Hpz6jfDgmRdcmFhzdM8qmo/jgLAJqjlW9u/3CclL0Asjk2
6lD0Pf1VO014WHHwx3dLuQ68ZWY1AiKAJ1W72FpmChVnqJD4I5p7zzN2bBvJxDOk1nyAJKM/qftE
+wNuTFt0ew11FKat1WC9qm6oK40CLfGAYk2upSr6ROPiDRlPzgpwMY62pPS7R/J87r3KO2zPJftE
o2UjYOfbecsruVs9s7bFGZcBcrg+qpiEPWHBraEiJXIeSHVgtuDDtdQfLxOFMdCoK4v6pbZsr0Lu
HBFQRl/IHWnYft/XtT0VqMq7gXmoubuvJnq8ywM0a9UpN7lG2V5vQduEFf/SbfkyJVU40VEitIa3
/R61lORNDLoM7sL1oV1WePZgnObH+xWO3l7ArE60IosfJKivU26T4dJVuEiPIj+Ma+jmUa0AMFXW
Fr86d3PFOAHMOHY/TADKXSi0EGjP4iMDg0OF8F52wQkDu7SLmPA0Q31gKY2JmSm9322CQULGtbK3
9FLAj1kVIaDrOfSoOcu+Vr5+hUiEKtTkTwdLIvcZtz48DQr/IR9CJh+coAdydVoGmCWV/Kete6On
NSYxCF15pO75NRmW/TUeCXZAHDKyDoltlXnC11SmbkZlW7lG9WwoGAe+8Pt/Z/nUAOiAitvf+gqJ
u6SbqvEosWDlaRgfR05jA+IRTz5oB3I+qrFCG/Uo/vG4NAx+nAq/dN5yUGgzKkjVaAiH3VLlFXTy
CTl1g4wp25XDoaAVAtZUeBaLHzWrS0OgpdpJJBCLBv1TnQ050DBKUilCBK3xTM3RCYH+E3GVbVhh
A4UMlImP7tXBv0K/7S3LFmuDnjL9w8g2EQBXhF9wVpwNG2XR/pG1VIy1Uh804WRcxdqoEQyy/aRl
pK9dM6GySN+KlrmG/6pBtxR9PmMiyudJy6vVr4SwIvClHPlN1gViI/s2gsWuPAOFJJdTD6HMuUYc
Zh21iWKk0AoX+OkJSo609X/rkBrqzSqkZSvHr0Ro748ZrAYis70NbcaYYA8o45d6tTVaVvjUc3it
RQkmCAYtJqSCtmhx5CwEodOvqY+1zVZxcMwDzFsM6iZgJkCEFUekQi5r/CBpoOg6kKK+EO2NF9A1
0cOSYL2vESzI0P+XoEaigB5LQ5TP83UxCIwnFvzD47c/TS/0SlWC1R16sF0sJWwHqMMsCgw7QTo4
3s679EaAVgU/RmnxqvMmHK2jJxArRplzqVAAbfBzLS+EAXnf3GCCa0OQOCn1HOwkwloIM93ZA0Op
AjvNqbgB0nZj6ZzkkRO/DNJLfi48WBAgFHsdBSMoyptGAyGCGfCNzS0jOKI6X7C83Yqn+wm77TnS
TnLP044ZPBHQVZCUaRFJCzPV04DBxZgDQ2CfSgKrp+oMF2YYz/Raq/er2avEnvO9gIdL7MCfNnaO
kBYno1PZs5U4mjplk0B2G7uDMqZqnW3hH3yMWxtA5Ih3nh3PjCVvwi830tKx1IHehDBmmXOF9EZv
Ujt2Mk/5XoqLNGcv69pQZd7sp9fy3sGLQDXl6AV8Nu4yY4ElNfaDmCvTC02Od9DVxHXRLAlbnI+i
AqNuAgueTICml9MZheYyYLS0qBbEWmqHdJeHfLwXHmIVHBr7/gOc8YBTBjnlQpp4A8oHuQAYHliu
YXJhizJpGq9U3osnIHpfTd1xy+d0AsOspsYlq3isNVA8rjWNGWKYBwqubmD8/KuEoIBlG9nj+UJr
Ya1Rd5nSTWyBzgRTqLqKZAYviKw2ErA+CXEYFKs/NDRE3BIeBWXIB6twhBLsI68zqSUhVn0C4+G4
yzNi9nBStyQ5fDX6fGhqI3vnyD4zTASu+DT2EiOBfgga5pvp6TU6njkeKmnhMGGhfLSOzs7batFC
nAm3ybRPtm6+uncUpt7JghqyzGkKLD/M7UMJU976ZXNpwgq/37H74sNfYefyqZ7Gua+5STTu9p9/
KsJcHxojEI9Cpf4JJLnwgGlZd6Jgz8rqt/0qSDQayeJiWchr024NPKElWLJQhjnPUFWuY6ZTb8Kw
E/xYAJaSFvklkTc6npmEIgwpS8+uFT0QZLu0LaCmau+8t7qqZky9TIm8aA1cNJYOfkJ9kA/NvtQc
rJk962DjwYoCBJH5SRYoTpyGgXJseUQDY2IZWFOOeb1zPlb6wesi2mrpKB4r/LAik6izKuQNizBc
al+n4OMO2ZayHhqT5HLQlWPdWhPW/+2BqNCzwTt61smupYckXQ6viqWD3y4UpFn5p23pSUVah5kJ
Nppip1JQCD30C6aCKvs/T6xyK1Nof5ZwAdbeiogqU69bXZyO7+vwYfLtLTDKmOuDEovv0IHahDMC
zI8Jw6IIlAcpW8MB2yzovlCQRkozHB671VkQlSE49M30aSgXl8aLhxfeY5cqIpSRTknAMNhAlBGw
fQGWtI7bd+TczchGumLKQLPDTekdw9GMLuK5tXHWfRS9+y11yH1tvEwTmRPYfZyMcP/v08PP6ubr
xHCZfL1k7CnfvSwlwh6/YeHQaOlScNePq+zmdf2/EDyJN8WlKsKbn0R+FnFNi/nEHD5AHQxJhyjp
lTTE8I0ea0vbeNYo1z4VZLP9KFMfunMvTppb7XYfySmsSxLicVOFMrTVacKIpIDE3UMbq+jIZtM7
OTE30ezFy053ALFwquMZOuLYQRrJFRrfLylGFp+3jdZRdioXSOy9EtsuLE266QXZv7EGmFrMRsSa
+odbYoknlIfuBfe2JOlMdmSI5KshVoc2CzW9Z9tdm9HnsQ9Xjza2bC8i4CbtGaG1zATjnUOx6OOA
202/ACbBinQrnOZGagr0QB/ceo/h7nZwPtvLi51/rjPeZzcLpkXCezoKR+cKGg2g4oxPX7QgxQ05
6rovyLKI6p3QUCEcmy7jEcxSQX2psAgYFj//wOI+aYBj3PbbiNcS1vIL44LG4A/8xCS5q55GZR8J
HyOvsMiX4O4sIA2HA1KXrPg2JX3kKRikiLhrJ4N6Y9OM+oXdGk/YKDoJE8Hghxs9HuVJwwiMs/Ax
N2lQVLxKXS4mPi4KndKI+kVTd8gg/O2lAcNpAIl+eT6km3uD/Ns/VWtXclTWWjh1RBlPqHPUR604
UbkLSYbU92m0xKNgbsNZs5YJGXQHDJPH2UbKOVXn/7HSRqG/g6IAzgPbtfYnM061yLalTKI/J9b4
9YqCZGK8nKzMAINI23zsrskcbNrWXsSXu8WEaEoLMklRgLaIngwP0Wqh0SSzbGjz9VTKTaj6ZAl3
e6qD4IDF0HVwv+snW+zMszmLV6djvV/aWf3nDUClF5VPPAcT7zOAvO/DWCTft5pU+rIqPKKQc8Hz
Cs1PO5AkGgTsxFlhzX5oklzhiLdedA8kEvRHfuRQ0W5o518NrV8JVjfoYgDQtsPXxtOP7+hOwpCA
yGan2pZmeq7/RKnAldR7gJ5hqIt3P1KDCciDAxwP3kwE3XwDzdrloOina57cifgkVIL2yI8/bSM9
8TJ6wzLhasRIiwR+Q5sPCLTP2VgZGQ/xAhXBP4EKen+U2+7vQpFUEF+wttXOZmiVU8jbNeKxsONI
B7KxM5gWII7u8YNpMKlaq/ZTMsMkamDrzICTIaNJAVyDyAPMxwsboR0JEkfcBhCVx9BZ3F4Z1Mlo
gDVyoysrX8u8mc1LKf7msrNphpqrRszKrgBpvKroYwbQO8GBuSXoFAOn6CH3C0oMtTLk7gHTujCN
3E32/VC68x34A9R28XJwNrMDnViBSqKgmQ8j4L6Qjnt5STsuA3BrTMdRpZGrJlC8S9DtSeN9t7a1
FYIlrLUPNlNcgWQvnJpIjSqi+aHOYlFZtI8RGzT17AEYWwXDZ5XeTp9lOpGA+ExUd8AbX4TzaElg
yKv5c5XH902cLXm8LROCAlOuXOwZvEGWygnSJl7Ux4e9Ak6AangR8bJ8Bug3o/EilrAVF8vj+Q1w
KWANC3sx0ZKarIewOrUgfvgz1uOMWV7TH0gTDza9mPvHoDyTW5tfXIhTz3d1j98lbqPw3FnSXNx0
ZcPNgw1tKAClOuNgpxOrYgfTsLTowG2B+hsYVmfqwMmTxv+fQop1wbUiGhOdw3aF6uFvWecsHFfh
RyXATYSCHJ75OsjSKOs9mShqZmUUq5ueG6AJKglacFREHqN4h6z8s2H66Rk274eymvpLih5mzVtC
fbrKXnpkVxKoAh9Kyy+djsQTe5jljI2+pZaLxScPiPhFtGaVBG0G56HKt3RfxFdwahBptgKzPht+
KMK5sKmYsJh25a1NKXC31MnW+EaFQayqVXZmAwP1cG3Rh9wG5KltRdoUD+Dn6xoQRnpE9rk/iH32
F1J9rxiPu7zuhZYrsDrWZa9Esowz6Ucwp/VneDCQLX0yeucIrV2rToxdNyLejPJY2+PMhoR+F7qJ
wDDmq7bu2JTXtyPwoRNqfD/6Tz6z96lE7l8ZPiSNQkq6aWrw5uADE8CjFZtgWkJcU4InGn+t4yTs
u4NkGl/eeo0Bex3XMxvvq9jvREwjQMG94bXPc23z+6eC7acM75EpDelRvJLkIe5/aeQ913ysVXNJ
LDcIL/+n0eD9GaxCE2+K7+cBEw8G1mKfzQXnZrCmX+CJXMe13mWVOs1hSddLLftFNWHGDfN2Cp1s
c1smsJO6juUqmF11sG5kAdvOPIb0FtC1oNUg9Onl60IcgINZh4Xm5jSlBZmgPqaFklnk5icfJgwP
BIGgzg7SBnT38fWzKUNmyMIttK2ykDhc7vrcMg+P6022k2mtDPY6n/b8YUvUPB4rkawrsJjLpwuc
ddnmYA8LEGleI2GbMENo0RRr2W4I36p/v+FNI2objKXglLOiWZglckfOm9Vj7XMaegt+4+GH+jTW
r2KkMpKTc1ToDMGjLs9XlvGfYeWX4QpJUmppQp8DxfeiM7wJ8xxqrmQb8mzi2mDLxpxPRBaag/H6
ATneRRYMKAXfytl5wMO7C2R+njX5f3u49hV95BUn+Y8p4lXhZlb22UhDSn0CiZAvdW4Y2jC3k+pa
Ax1quMtejfbz/MoVTXNN+xu4yNKfWWWiw6Cftazi+fZpSDE68Wka0X9BvtwgpIrF/VFoMAi1lCw2
tkBEPnxhnfnPep4kRnX+lz2swEB0x42uNYpUBNBIBDoaUuHj5hzsNlVyM10CuUb24pzt9ggv8m+M
HgJXlvW1To/uSHkJ+ElW/tKNo4i43z2fvKPLenDwKcwzuqvqWeQuqGszsiJHb8enHuK4lvQA1oI4
96e7I7yqkQjCJN1Drz0QbYpilGKDP66O8Xl5wibp16iuH+WlKzLcT5mpgOa/SLHDTPp9vzlOPe19
i/XTzW6XNnz5FprJpruAA3q5A53a9Up19NGdJqQysi00FPj0lvTmZAKkACLS/8C6NF9OhqmB0jrA
juJ4J/RP6BKH+8rHIL2u0tzz4HheFexfwE4SE9VmWio3rdYusBmGE/GTeWxx4gIi6aob5AZ6qaT+
vIu5tKidbHYIfSi0/0Gowfq+64oDZK+lEIjQRLW+5wjG1TC1YXSww9iOE7/+h0/5ZYCdGM/Ogxnf
K6vphX3oUlvvhP389y3AK0KSss7koCxmzEKJw7yRED8sDfuQgO8mAqMWxY3uZRkmS4lo2yXcc1NU
16Qg10i5L3jX7lrCKu4GjEh5Bw0b4X1Ko1rsSsvMlIwr2vaAD2rM5ID72/K7fmf6D1SoyMfc/fzp
DPgUrkfcHfFfGgVaO6FHsOD6I1t3nZvMNzcSXFDWdxiFxWsrTjoxINuREc1f3wvN9AqiiMLnSNG1
VdYmTLdgiwjeJQ5qY/WjfPAA5ufHADfTod6r7Al+s7pUzEWFpyLBq3wqj6j9njXdM2SnqGXYb07+
U/Mq8fyX9HUYedYjQ3NI3Z+cvZR1oZp+thPkTy+sJLIATXu96eDjqmdOX+G/0inRBJf4vczTl9gC
dG7HIlq+k3P7KP5OqsapHmmXTQ7VaKYk3tzmPUxcAXooLpU+m3XgllMWeBp2Tiy4Up0aNXwDlIia
2DPzQknl6DEFeWJOq942zFPoOiOuHvCqGh9upWaXzwqbrb1fUd1nXrSwg20IJwEmIcE+O2RL9AxA
/W1Twsr+iordayz6sVlB7IUQdJyHdOi1XZtER2EcjX5DjSP+oz6eiAaeUxCLK9a+mk9ub0pcaOPE
q3f58uQPYwT7edj2LOi3b4avB+r8melJWpBKrvBIxrbUznCX68mRIYXjxJw6xI3VvgCwlmDHaP81
/b7Td8Si2sZw6GXuWN1Z3LgDGRgi0k+aglGGDvseCpoWerEA+OimH2ot3MbIQ15OGpDuA8ESh5cv
D3JzNFWBa/5d+e1Fz9juw5qn/tXYjRJCBVuGw7PvF+hc+OShTD4btTeXcXJ8DGcE99Z0BkYHA8KK
MlN1545L7V8altY8myeH7UwEDsAqKsKs6hZqCL5SsgDUIX/bXxRTSwqpHncXrn7KLjGDe9Bn35gy
W38AUKGVUeliFiILWHQNe5VBGwfP637yQVHZY84VTuaVn+5RuJAttJZOoHXT+d2CTCDm2Vmgxe73
of5Yv67gfdTO33COAiv8RV1BnzT663mVQNK/t5vDMfufuYgoQa1clh+fYOwukTn4zDJNiISYduvN
I6UKCxJ7w5SQIWLfohRsE0rCPvf6kVTrZm9S25ku7Y+M3fkXyya9fgTjUtDdqKR29GWdDDW9/ny0
1hQnOMDjpXq/rqtaoWD2gn1zNAC7OW0mXs6r3dIhKKcObzL5ODTJ02OAsZ96f1ivfdtsoq3sXW1Z
ThcKi8XyMWMy4E3LsAihUl5hJ7FCO1jkMJSqQYIGrKhyEaDrZOa1wp3z8LzzrXg0aR7fZ9SodxMq
cRTUD1wg1XLUhWOKcHIDdzvlI6XEc4z3ZVDoOWgT/hWnDiz15zlDKYeCOwv3R2lHP7lfjgJvBepk
zOwTXbQhQsVtsYzbpbRddFZtut6LFRfVgP0PtlbsELm03R3I13Cw7PUfwCyvK++4GWp1GPk7ZCqp
lZQj6WoEU0khpwmDx1/Jls3yDt0JaP7QfRPJJoyXiBysBG0Cw4FvSxU6WdrwA4Sh8WZ2P795bARE
tLUnmQliAKSpB9pPkOlMTRT54grEXIIRAfmCXips5D0SRVeBFr30WxXN0qFnTLi4d0Q2wIPs/N8F
kyZEdugN8vioUlGImg27mHRxVLPPx1nZa+6zGmCzOf14/s5pSjBc88Wb+78OkQ3mqKBMkh+q5UP/
B6v+yDmEPCJ7EA/kSNG10lfp/jqDVjUfzIYrcAWDxDbVN6S/WQKTVth4NbZLl0jrAAlhvqtPxQ+x
KsUp8XbBSXJOx1xbXmIpeeDrpRJR8Wdcqme0FUWy1G3bDVHfArJEgXqUrBZkDFZ605xRmv6S4XTw
dwqf3eGkVeoYwdzDs9fm/VQRhwJw/ZyhA53GHMgPl2y9ejg+FyFTn1VqBWkmjFPUvHHJLcnXrzMd
IUhElaHnh1ftccht8BdGTYHli5DX9/AyC/kUGlVZevDJr+tVNKO9eSnduSpyse7bFkVw8fL76D5M
TIdcxhaQSrMxpCYoVaG+SzLWmQgn+by6KmCIaz9RGtPpaKZQI69njzuGSykq4PXjvB09ajamB9/R
q7gLzwG24Zjcz1sXuXtqOzUQJezVL38SZ18zkssnqZnJbtJs4Z5UtKmDxWazkg4H4mDicG8jeCpJ
e/TI05qkBYtlEd/pDUmGJ12COHPFLV3Zm/06tvTRon4kZND1oWPO0RcsJ6SDXyqJLXACZVhfsz0B
kEP2e7+0GiXh7MAcSCxzAo/gAnsmzzPy6LqUGFdMOGaxMiUy+6ByTCY3GDOU0ESHqloRJVwFxtC2
QJ1mrHyAjx5mQGD1KOkTG1LooO+k8FYnddzh+LUrrwsWKp9oy2D1760G3l5kZ/pPbttyOsoaRXa3
+QxsizRCF86RhUCTCDnB8q8xnA/Fk0vdYlNMmpym9vu+ej/IyafZgdd+XskMqKWvYR17aI8fhEM6
Yg0LqMIcnkgJq2smOFPh+7R09BbArRht+0DZxVJbjPDHRCliYnR5wLobpSqxYlsvj0bjtyNuPw9R
xkfdmM+W4ZKFEbyXalAlofi7X1z4apeFmOOQ4AQRBpG0vBP4fXhiHm9M0D7Mt2IpxTxb4vA8xVTK
0ST+VTja50b1s5hcHkklf2CbkLgLslOpUv+9hUP+VE7G1zAeXF9N6+dy2gimtI0i2o9jlw3ouvEb
Xcc2iC/TmNnGbi8AGaSA+CT5BdnRDWd7EhMcn3vnRgcvUUkc+IzKXw6AETkWyJE6T2945Jzam58d
jATucihcsRY8eKsXR0LEE5krH+gU9G6QyDEX3bwFSTyKNRuOlQ6ri2H+KFNcOF2P6HWjAGxDZteL
4p6btyXu66vf1VaZaXi+jiYOyM3uOudcjIQEBmytdCVabIzxteZiBjp8DJOZPd0QqKglQF8vufSd
DIiUw2dYZwKXofPWBx57MZr3ws5iB7Rkn54S9Dl1VypzcSnAVV/SHdwF4Ay42VNE2uca1pyVm650
0MRartaUnLehJwnyrFS0VvAHMO3vwYTvWbDsxZ79/0sicRMQh0rZVq8gkkEIns/pqEugbsyc+s3I
bx/NVkMJf7ciMYVpuokoaQBcUb8X2xj7hABfEmdWuFZWx3pOhH1SFtsqM7wjvqjIZ5HvCwcCqxm5
SAd6C8g+Z4LRpQqiybyqQJvmWoCtn2emcVlzS7O8/mnzdUtNf1mWUlHB14MCGMb/ja87/3wde0UJ
v6NtI3UsashLo1xRWB2uVykiPqDbs0i2jIxzytRveBxqzDKoC2+43rJnE0KExelnpUWDYgV+AgRA
wIhBAWHUwE4t59xppZty8uDsWSBl/nbNBWK1y2wKJirIWFHaHOEiW3BTLuHXjOXdcz2IbuNjm12+
HrWLIHhLxSAgwO/BQVcN9sXTJt4oPvx2z9ZW7x0mhFb69+msvMSjCcMYViMEQ949GF2g/UM9DZ1C
ng91tmiAnySTAaC+qCtthIa6e6VdaPe2bCI+GHVw8iJRr4yuRvcG2hlNQTqe45ORZPd7Jl3o4KKL
VlndoheVhuZchGiGcYayXbLAOWKtNAuvHL4piZgW8umlgnotm5z0dt+JcmOlmjSm8NsrC6rro+Y4
vOcYVpFyhlNDbw81lhZPHmas3XdNTEtfltGyvCcayi/c35f1PClLKr3ef9Qo+TEIv+Tso+ETRFmv
yctOcNEC/SwPhOBWO2bUN6V9N1rGah3hwDGYirwYx+1oOIxUUXAUmf2aEuqxbZFatecKJvtE4VEk
tHOdqDDSd78dvJQjJCCb/PanO/1zcr+b8t1s8I8MsbfspZJFPE0VotJexaTx5taMSJo/1FLIJQQM
ys9j++c9UO+xF4UF6vj7p7cKAs9io298JLqB5cEjvrssweWcy/EaX+HOBozyXPfyEhWU7I8A8bSz
mthK6Ig2mm1SgM4hROyOCcKiexkOBrgQQRwG4kWM38ookRzKgn7M40CHG+y3u3hS2bQZwyvLbAzK
AKf1Q8+Uyj/5aucUhf9pbGMu5W8+xFOYFv6EN2LGHFYc+HoZlMDSDKt6sSVR4VRtftC+t+lO+M3S
Ej2YenWvWT4XOpJB6A6p3hkGi15WRlQ6DePAwB5z0jagX3h8zWL+H7w4wxmNc0uwNAGiEjR8pR1+
IpmuiTBPuXeyT4qi77Vno8CVO7HAcpvNRXZDVw1eEKTL703cNQ9NuH04OiRFUDUv9npd5Naa5Yhu
sT8lKiWlQuVf0WzgTOsjvp2YPAJk/fck0hNxSQjlIHduKSUNwF9TZDMAsSSMm5PiIWdT/tWLLXIZ
rpzWKebxaRjiyrKoTw957v7p1x1QMIuimzPa2kGCM4eJ2RUz6Rd1B84NLU5cwJTBDDDk40g9J4YQ
efJjBXbrk6QSaCGiywdgFYqsELTlIWqeSMXlh/9PWX3xBKBMNNftlJ5TG46fKX0UpQpGVkR2awKQ
Qou5s9v/hGg11Vbv64/mRiA9fWZce/gXT/xfUdaOb6Yqhld8fJ1EiuLaAed++Tibu66StfzJGzYF
8cqglx7X/D5RbcDRMAcSxUOu0T6jRueRX5FVFt/jKNzTK6PD/GE2BMUAZY4QFxcu0OWTdZKcRsEV
oxEnJGzGpei209BLigm9YMYMu+Qpj9Kzml0+TSBr7e+tTbjGIdKd2iLd8ZHjC4M0fgVjaIxTUD5J
dT6NJUkgTTbL2a7mAnqeroMlnqZDK93L4r0VPbOIGkCqq+JGDNFcD0VTk1zob+bZNaS1WVVsbWYU
pNsnCjUwggUMoyF+Gvz7yWj6V2dUUr82ztTvnZhkRa3PaNjHITBfPbQYGG/cbgtaa40k1ULvGNZ8
iidI178HfebJLOMM0j/iQfQ+pAd1pBW3111pvuJgojE3W8yo6QonSwc/wueqz0AjZxEqqfPSGpg+
rKfoUwKa6dtGUukB1zORPW82RLbwDbgCRM4m2nJahPB5gUkiKrXOAELs7M8NjizAUQGwPFoVM15U
z2cl9ScQSuUdKgUfxPjo4M2/aIjaDIGKPU2ZezDGmWZtNxxyztdZuhExBaZlVm7lhva/CEd27ETc
ODz/oM5+ZllMWqOzOTo/HOTIYOxrPU7Xdxn+Qda/tFFvWc/z1CjR2zwVjCttNCDr3Ktt7sdYrU9F
5mTplWEiJ6X9ZHqHDaUrCg6hTUsglyJP5DNZRKi7Cs7p3rNqu7dPSrkPeQUobfOzqWnvyPvMMXAl
0L5r+5QIBfxbGZQo53+mSBiFru0JiIn/qH43DCoYyARICX50mUSXxUdRrr+0PLW956ongXl9iqCg
4dTvgKqpQPTgos7Qa1gYZ1NBs9RGAhMRA/AQL/rZJC9FG/r/Hs7RRJeQExxE+EPN1tj9Q/PMPAJH
kwuROTimMgid9dbnd/XdB50Dgd42izmXdCCb6Tswe8X69yIa2K8B/3raauDsAxC5f2Ey8oh5MG+n
g4ZhtsJNLHZJfOMOpPJ6R1RxNkeb4vjxN0Wr2ozLrCrkZVjdeELMPuuyjtPqDXFLNdu613pEvDio
D5eijvVQ51MalHUdi1sBHVDbU/B69lBrU8JnuDgqms9UWCZDvfO0h1vKTZwKVby26m2zjDSDULn3
6WnPWg6T18w2ZtBcnn1AaHT23rLMzJjVLPueLGyrjVl+emVTcvCg76vT1LxE/6G6V3gA8xO935Le
f0JSzN9E0CiQJ3zS+XyzP0TR2ocLbHjuK7ZaDvuW8cyBLddKQdvceZePUMAmPwzcebDhJGcUMBoI
ckbDJD3WyuHjW/gURBofLFYQOp2k4hOj0Ya+73G0wvlRWGLrQnY1+62kDtYpgNQvLYqUDF+omVZl
HiNneFg6K++1c4qolVs30A1RoWjXK1NHgs6tpTPPHc8B8Ff2GgM6DRw93KfwjXw+rPVcwfynYXNI
iTGpZHRxDvLZVADypGHkNLUhF1mWjLzjCNJJlNmGOznfRwTl4SlnvQtQVOuHMx3lIjtoJMbLbUqZ
DmtDpO6xb+3t0BSnW6Vkh2nDs5sVrSeRI3pA/bPHojGej8xT0Q7ExJTU7iYzFDtgSOSskrphz5eu
sJk9nHKxjaoB5XB2SlyhURjEhmDGUvGCe4g2RP2/gS5M+LO7boyR34d7gJWGjZNN0dCsB4ANNuoU
zANbSXTCwlDNJM74VtegKZNV/zlQqwxy4z0+QZxy8X4kXpkf2nAG/FN+zFkt/i5Ue9HCwx0Q/1/t
ladjGHngPHbrjiHRzFzD7HKPahlPBDYhYPCGQo6lvCC3l3hUn3OGr9MOv81H8AAESdLK97+IejiV
+j6VRjj0bMugEdPjXMcWY7BH4z6RqOIFf6XfiUFBbhgSft06TGGL7ENBfwyB6RFAbkmh16ecI9VQ
zjzyJcYUabbZ972WrR8mlZ9cwOKR4sXCoc9e/QeVOG2RvrRX1yAr5QC55JK7AnvFgMShKPySuopb
3thHtr0ODNt0zDrFj9px0X3SZaXjdLG1ile0hrxnc60PMT9D3C+G/5cTpiYpzu7vbB2CjrGyXyB6
KU6MyGJBfKfwo91+m9eDy6SwH79Z58ETv9ta4XYh69VvbpoDPyOnQsQ5Aao+DlX8cL4mqoZOVM3/
SQi09URzcUOgDqt5+t80ThiRsvdDl3YMWbzN0Bg//DfQDmnM5wtnriLlGJHJjXFyDUaXTgbs8w5g
wpUsDWaQrGPOyS8mb2og0RHAuj1UchWxz1vf0qhmtoqAmOD/zND2C/Ywmtx2AveEH2gAsGtMN0SD
Qi4weIE6sSs60PYD5AMxf32NzXKzrsf78qyFM2cThlt9JrEI1eLRY6iwK0f9zdtXGkD7h4INtnx5
54BwahXdZAq31XAhtcEElqWVoPTp7sjFm9zPZI79iBT1z3xZDCde0+3kOtbALQ/uSVpqBr5rzFaX
IwxpVKVYth0o3ZUmW4FxMWv3wkR32M7odF+BLQq/T0veCzfw5Yqqki8asFJpL8/xT7e5dmBDhlLU
vaYlQVgozknt1K8RguYiBz6WqYB9uczgEclBHtauKoCL8f5/UFImM2aB7S2wLypwh1qC9eYWtZX6
CnpIi4QMogzhY/YhnIicjyxUdqgOHRjiTu6Ow8VE89lTnK3QvQ1r/Ujo86x7SdxfuCjFH7f4LjIE
QyvtQAQ4PsbHNLgZptAYclnnOtyGKe2wWX9yfAwMmQCaPYoEqyWzki+FxOBUHw/HpFTW0AqqtbRs
mTLHSDxODmQK2OoJMU4EaYZoxqEiLYSti1PbcX1XWr9gDZtoybkKSNBSqnS+Bgd8BdJ89w2wYXdq
fjnHjS9e/fEOuxHnh9mAD3vvBJS/4rpwCClBsPbJv24oHNDlpcaTuM0qQDR4vNUtSS4UJ9X06ZHR
XXT/Oih21smQFAe8CyNmELwMbPVSc1XWbvH/kSgQ2ifnksWVMqXlVbw7JA+xl57kqkvglD4DVVoK
kNzIHHKzBtkFr9MdFRarZyZOttGg+411bLSP0qd3rxL8H1N6cDo4dKpFHSgZ2acnB5OI2qJoIla6
LnTJM0iB51jbdpxQmgCan1a/MpQk0DD33Nff+oUIr3UD54fru9a3o7RIVIgMNi/IarIJ7jTyD9oZ
tlwH1gSf++2fp14lAjj86cwsUMG/LlM06HKQwizo/+N1UMB+KPh48B8tMqscdN2gV6HGBOcxxA3R
ncXJf3xlz0tDuiDfY3FTxLIHNZH2nQYis+TYQ+LwjC980ftIvAM3vutHHBJq6MuRev9HAyV+7tKE
LZOB5J303ASF9Injm3dqS0ze1UL/K9TQsAWn/K+uzLbi75RpzEIRP11tf6TJ91LfmdMJnXh4/BHH
QcoyNi9z5pcrgJNSRPxRvMIl2cNxaZPHS7yZoyNaRTRa6feIcg1U8Co7jHFyOT9fcaB/7lkCuxHf
qg71eb868bzEYA0RQx7feiRUYJ+Fu5f3G10GtAsqHbSUTz9jEz2mxj8YXB8symgNNFEBXURN4Yit
PNA6gFg4NbXI8J5PkdEya3jv88YXu5Rww9Z+mGLwUSVkaDY5HebCkwAkup0M8nrW91wds6q9m7KZ
uzaytSfMARL4A0YNSR9KFbSLLbAxcyLn803jsjM+UK9kYhjdjpjGjYjm6iFM9P8+VtPcSCvJRcNX
5/lP5lrMaebAzLtVHFqcUQlkPu+4nGkLhIK/xQJhQyug7YbMvagugLxiRZuaxfFERs24ZvqTRxbl
zlxxCD9+DUGZMCnGF5JmzXQ6tMh0xI8pbllMsSWkrLZG3SRgobP70VeasN0HxPaPNgU+e8lHbsjA
XPo/Hw5mLUBTIKq8fE+MNnYyijTANNFYhwM2FchQzddj+iuqzyZZpnsrTsAzig6y8zLqvIdcJgwJ
Gbow0KSqLvbl8pB+wVcZQm580kKtwwAUe+Itk/Dyg/4Hz6lQPzOrDmb8eZ9rf9LpKwNFR1W6jUHO
WEXo2ekYPXcaWsVFyPkj3xfFL0s8YQ9dGTyHdnW+MQjTuLisu6YFc47dvYtOWsuV3rVH3mBh6OXi
9t/CYKEhmxdoDLrzmVEv7lh7ZjrafMgf2p7jIgjaBwgfQ8zeNirD8gi5QuROrc5D14rZWvyDDCkH
V9uvsZtJm2fXT1IOAUfjTYhl73zqiE4Vt4I7TlpRm5t+aOhzV/Yp7BMPKADFePtG5vMgbc8i6lfd
u77kJC6sLtYzin/y/OJ+RmmML7tdjIJUYSM8bbh5nFfMWyUqUIygjv1/XUiV/IT8G+ez95Mip5cU
DORsanPP2lGnagMEOhl1YqhfIzoNycW8ajkoeOYrSVuu4q7e+iik03npdp2jri1WmsSjyeQ=
`pragma protect end_protected
