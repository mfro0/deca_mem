// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HNW47R=A01$ZO[MCVO##B2XL&GOW^!3 0?-9&/;[9B0H7#15XV"MW/0  
HL<,=M>^9,?*O_>_.HC/;5F5!4H:C? 67:$S-,WV+>FB2/&VO 6H=M0  
H5%2>_&4IY$S83*!9NMUS('RD?RWZ4\6]VH/%'J$ST!6D@4%L[':RQ0  
H4*717.#14LQ7?\OI*IU@%;%E^5M I$HR&9E,^V)ZR$T+AJI4&!8E7   
H9G/+/ROEBW /;B&8DH=EB8PM,"$0 >B-J=[U;K^F4U$Z=\:#;\&!?@  
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@3Z] Z[ +? 9VF?SLE0?%(0S>LCU]$9^4'Y?4]';G/ @ 
@KFM$<K'JN'GMN>Q+)&3DM+DA.!D[>Z>[-BI(N!>:?]4 
@3%:"QZ_N&W7>@F]+6#'8%UA?A?BL$ SEJ_;/H(/F9]4 
@0I8AZ2K#JM2.M.LZ.$P!ED!J08G1PY#4BT_@;5CA&N0 
@7H4G\2/)+E*G390]LC%Q\GF))-K_AJZNDVNJY[FT!O\ 
@G/OVTC^W#T1C5%WKF73(QT9G(Z$4PZCVZU6.,_H-1G4 
@Z6G]8-E*P^--<P3'$]IVZE]TDH)X"<D[3B=M[D$H4 8 
@F%\F_@?6L'";<-49IT]KIL[%4!\\HP:ZN7"V#.L8[08 
@X$&,R:3GUG@B05CO\3<D2[G[<0R=UA]LEIE6MLT.-SL 
@\*O?Z"J.BUHY[88-BSU36<U@\9S(W>CN+W4W&:C'MW, 
@S[^W%#US@Y62$\A-P8+0@G"6K=ZJW4%U18I$?AH?9"P 
@\WV<2[$>#Q&BM'D536,*(3)N >XD?6AX%$J(BK&GM>T 
@)CVM86*BFKGDU3?NNO,2^/0E0M#1Q/90"GI>-S'PMWT 
@T%^DHAR9]K-WV#S_HY7?!J"6XV0?4S7T&Q\4)97*TS( 
@9+/[@']-ULB:0V1=L\T-(DT$Y)LXSTITX@+T89N+M>X 
@;61 W-I]7IXYO/MVB^B \&\H%V0[6AS0,8A[&LEUSU4 
@HG]NE$A?#.Q#ZD^$]$X5]#.98YZL2X;*^\O=RKU$]!< 
@P8ZYV93"4<XPX>.GM_&>,,/__^"PT&+/*M3N]AW6Q $ 
@.:_I(5^/5 D'V9HHB/!5]$BMK[8XAZ'\/%!)W+RJK+( 
@OC4"Z>;U[G6GM.GG3'[]Y@6_FKAA<%1Z0OT%E@_JT^$ 
@8 LK*$WBD=(9H=\"\:_LYZ QT"S2 JH*]3T$O;2&KY\ 
@!!H0(@[*C:F,#2Y^U"KL.VI?XXHOEON5R7$W]2/0?K0 
@GOI'3M07R])K^DCT)WHK),<H*/?2(T^J*A19/=@%/Q  
@=W2+K,>G7D!ATO^V(V]S"M4J*%2*K3N3RN(O?HTX7&D 
@S ,NSCBPS5 )[>&>%#Z NY:+?])*S?I&J;:WR<Q- T0 
@8'YDM9YAU-ET(CJ/50]K+%-I8<&"KV_I;23DCFT.P$T 
@QA3G3L[67CZ_P<F<-+E_K?PL(1QQP2"LC?$R[:!^"Z< 
@([*<)1CS=\8IPYBA!4LMB47X8\0C46P?/Y9<$JHEBGP 
@EX(^5_?'M<EECA"=Y2Z21D*H#AC$U@M88\15WCQB"D< 
@-A'M9./XK%:K,O.R4;_25B(6IC4W3N3A_R=<7Y47.5$ 
@J@B+0S&%1(M>IQD/1+(C32,*2!<0ZL4TK!]1)9HT=G4 
@Q\Y</_4"#7 +OB!SM9Q/K_,I8 ^P0)++J%WQPZ;*7N@ 
@PP049]Y?MHH#WN1G'6X #KUU@MVM>I:95%5)WB'4D_T 
@-*D\9^B;(XXIE3=LQ(9VHP@X>&,!@@)NB'#24;6-H70 
@C'Q?"#<N;8&X@47^STI'0V51;?PZ$$\W @MZT#6D M$ 
@*36WMEQJR_BH&/(%LBVB=BLY+R&3>JHJRJLIFR6O7"8 
@&$<L&\U4L X]O^3NN1CC^FH-IM3-7KJI.6S7!BIB"RT 
@A\GK^O_[9A/$TK_4A!4;?X#:'K4#RBPU7HY]M,2&*AL 
@Z$LU;0>JTT5K#2TB;Z8O$PU9ZY5$9?&<',$J_Y#BAZ4 
@0Q:K[$M=D_,!?B/(V3FB57.K^MT\E:OESSB[EGQ-]6  
@'FX> Y&O=PXN*.?J!G(:F$NI6?>(EC\IG#/C;JL0>_4 
@+0UR-,D6HKE>_9C.,4\@2)%%67_65$.1>.[RK8Q*!/H 
@7NZ$]ERTA#@_P":0U)(BM5'/)D;_XXKAU*P$1)2I<.( 
@X(./&QHUV=S;=&D&U/D- .BO42300$;(81P7A%L"I7P 
@6 @XV@>WJR$#>"TLZ5BG1MG_^4#83W.E>H&02%?97B4 
@G+0QG/G@.6QMB(G4:F@M#^%P[_@OU+6S]QP<HW "#"H 
@?T0R_?(9&)H1G[ 'A12-?][N UT208'W1!\<8N]/ ,T 
@SJC7E[KH\#:; &FJ:6+\:-T4EW]G&%RO(X+U?1U5]S8 
@)(7G2,7O4FB39H^4N[]#&RLBD>9] K&91LT\\Z2G"?4 
@L46;>_M_W.H;I[>W]9PZ)W>RX.Z-<X7)[B<X2H*^E:$ 
@>_/,+[3,$N);R;B(-8?9')-04'55)EL3S?G?)I'Y8X, 
@(SOH_5/H2(O%TR:.:/59V=I#CW.\T@/0U&>.58C?FHH 
@GZ[/?H0$&;_&3*I2 G]W_$U<<])CHHN"UVVP?(;CO'L 
@%Q><.C&>/LJ9<XOMQAUU'LOGR,MM#O-_^8(7&-5/63L 
@JEF"08F<#H%C7+'[("_,Z3G;\++"9\-C-;CHLQ#;, 0 
@0&E.^&:1XBO'W6;==:X1_3<D<J#"9IYS5V,@3R:9D5D 
@7/JA0+ [NJ/T4%H)XRWW5#E*:<'=T"%']P@G""5>OG\ 
@?0!AY)(1XRO.YQ7+FFB!TL"R ZQA1)9% 'Q+\X5[=IX 
@XX=R+UW_9.'DR,/QO,2C,/]O,Q6]O[_.>R0XK[]NSS( 
@V%C1>BHJ^ 1<B_G9_&HF1MOI24+$48RT1JKU<EXH5R, 
@AIC%G"K]K4.=X+=;]U1%6Q*H0&<G54$ OE4$,)*$/<L 
@)!K\C[NN8PLJW&4Q9J;.7HYJ8(106/O:)&"DYD9.^7X 
@/)^Z9,BMX9" CICC%ITM["I:)MQ,83*HS!S6J3T,_D8 
@EZS",LB#7\A?&KOOEJ)'EF#_:*><G%%3E&5%WU5U?IP 
@=4-&P/JCI3Z>#QP<^!MRYF:ES ;H#R%6YD&TZ8<'1V$ 
@:&:>U3#M44'_IWQ--9I^1BT(%&LXW33OW2,BD+?.&LH 
@PBDVIPO:'&#\F)]? P0@V>GP08=5;TWA&)59_N.=.)\ 
@TO72%-+WF6+V*YN\M_2K[:JZ Z/Q+U6O+Z<7>8Y4#%X 
@, _I%9O)YQ7;H09]S_8<S+%]*+>L6W5=!5&]"2ZIWFH 
@@K>K>R%Z6KZ0 5 I2<0(=C5MB*:%.&SJ7=Y43C3://L 
@ 50M*-!]5@0M2Y@UJOTU, PU)B:FJ+3HI9C<+Z&V<(8 
@@!-A >R(UXHZ<)&I[%%4UO_HE#@P?KT:1\$ZR.9VP^@ 
@K<PO!KJ^JVL17\6]85I_?KWK?PLA=$E. YA]A;"\4F< 
@GL:^@$$/7FLM$JN='1QJD N3JYV^>$[\,;0&1UD!_ZP 
@.%.]JZB&B!.&A!9%\KCA7C6BY2@,$$V$N5I#Z4"]]VT 
@1#%3HO D CO,XDG9"*5F4Q'7E?]C5=:KG0HLDYYA<H( 
@V&.T!D_.1N^TTYE,ROY=K&@NBEI"/$7[RT[-G@W[KW@ 
@HF39VKG<?WI]_F=S.,FJ "W6L]/VZQC=ROA[$P?I?1@ 
@SS\,6$/F+3]?3XI]4][Y=*(G>@[:SY/?XCTA I5R?VX 
@'*76C#J[<,Z8]4\I0W]::_S68LA^'O4TJNCTB*PCJ)  
@'>WV62F=G9LJE8-$@ 5$MA6RLIY)$5^V/L+\0$&CCZD 
@%+*IS_,*B8=.=Y!WX0-C"\RPD3C?'^&]5V6<^TS*0+L 
@]/<'[YHO^F_:#YL?3(I/0C8,2@N9RBH\L\MOVCN)C5X 
@^A,5$CTG)6@R&(W5"WXTM<IG0636UC^J^CSC19.O'#  
@,_VU!G*/"MO8IP"?<># 9D]]=^3UJY;'0M&K63J=YK4 
@NH8^NASLW^>RDSQ?XG9O!DP] L&D*Z/W=EDIP76^"$X 
@ WC4Y$S5(7W''>,B\'*UM/1RM$MF2BK8=$[!CCP>REH 
@RZ1F,@UV9;.(Y[9(H%*%E(=8_WQ5[L%08%ZTK!-U4L, 
@(*3G:C_4O/FH-)]?M$\C-+1%>5AD^"R?O7""@>BT%?\ 
@*F'*/NT7^"C@5*?)]*)6 Y;H9T Y\_]KOW8RHG:>Q<  
@HUV40PCN.\'Q.'0M(@!\U*W#.+'<9JC\#DUP%_P=3G$ 
@HR)F0;@4B_+<?/_TU" _?J5SIX#PG;VPCZ!Y9V)11A\ 
@A<&(A"MV6)ORM+JSB,,UW 7#LN=Q<(*+F&--5T<(QD8 
@$]9)Z$;I! V0EYF;-N2;9-$2 >4/^&BR/-(D8TP /7X 
@/@"8"KJ F6^J&_B.4;ZI PDVY9%@[Z091CD)J(SF98@ 
@6R>M,[6*!E")C?T9/N1KH07^4/."BT!I60B!=2SX$CD 
@0FU\.T*R\"1L/YW#$MD,G&CZS[O =I'!CG,"G0-=$"8 
@(_1<UG04YPE@'_]@QG04 6J$N%TC&N4X:=P(5^94C\8 
@(W,'R#CV*:\E-H7-N<$4_E_2M -K4ARAF$1K1E ?],< 
@+>(E"O:7-37I45)9R)%VQ/F0G1+LO3)7$A!9<S*XO3X 
@P8!G0Z@())6TR+M?0+STTA7UAV._]($YL4!89(2X,W, 
@-Z#N2]GX:&?"6E\YR6WMVH^J8Q+$<1G4[6'$BVS@/EH 
@B233QE@X)PR]='*A3YHF\P^V53Z):HC:2</](AKD: P 
@**>]&@_Q^_?BYI"D?S70L)UJ!,,A!>CY%&:P.&3'*"X 
@.TR7\S: TF(OTD$N\R<1;28XJNLV2DNM@EP\N1>U61( 
@*GR__U,^!W%3WNA/*?BG;[FYRHQOB+'_*TU\VYJ4,^D 
@W,5UNZZ/PKFZBO7NM__8OT_LS?JW9 WW"?;;;.'NS/$ 
@TIU.WNHQ]LM?[O/?J^:J<42"+G.N'[?#].A>LH)?_[  
@ :MZ_S-N2D,[AVI-VXUI0V1%,QR7\N0=GFXS<MH )KT 
@M-QJEHISN=IAJ+Q&)&;DTQ-*JDR_;SQ-&S[[]KWJUY$ 
@38@*QOKZSN)ER4[1JE]3,>)BDU4<859!,O$EJYN=\SH 
@/VO+LBT+>8C5*#$(UT:KPNSOE::28'$=J!H.<UIIE)4 
@>=F^LT-]5F_7\<M<?=:7#,1R_U0+UKT\^?65C*G6=)T 
@TCV4B@I 169H2-5>ECFU56,H>IV9OZP2QLDFO?<;A64 
@(<(P5KT*_&GHX<L9"(-V,R 2V7SPU_8>4ED@?']-4Q8 
@:KK/;/7-4S80\TM[W+:%_@&C;)!X6"OE%W<%_T!NQHX 
@-$(OFI'F2.@@1-'O%^OSTU&.(27QU)2LSMKI>OEW/ L 
@# QP@[95A4YY:>G$29IM53;I>J8D.UV,6.:H['MBET4 
@$%MD:3)E/#^%Q8Y#H1B?#!YOU;V)K-K(M8C2@@=7O'@ 
@11D'P;)C277.J9>(UD'T1@Z4W9IO@Y(QVO8U*;(0L.@ 
@R#JP4U>F+7,TFK>M*%*+*%_4\X]'I.*4$;7"9(EZI@  
@6>UGX^IGMS284Z>57.S\ _*U!Y;H5__!'P#LM*Z^B @ 
@%5;,&?+@%;U7%L%-L<XV.!JWWHS%>T6DQ:E-'0#$ ), 
@- D^)]U#\3;4?3E0IKF1#'W-J8F5'LK&O!^$'B#J$ L 
@ECJ69=T'Y%V8="_MT%PN'8X'/W%;GXV8<5;)!=LW#4P 
@2<$+U6\>2CFT4[@QEY&B6/);B5B5^]) QZ*PZ=[KPN@ 
@"\1'('V2A0,^J"@$2%#>CZ;^9RD$E.M2'@ J56)2[/\ 
@+HXI=I_E2H%I,7O5MZ@Y,%Q$))X)4DVWF)4<ZO)["GL 
@GU4*$=8& @B6B"99&<5=,XK*OT+L]W-"4<[O*H6"(P@ 
@Z/1B)#QC-S/!S6NO:Z6Q,#,VZWIUJ;@3>)D0.\,HBUX 
@,W_4</(HTCKYJZ?H+<6&7INTI[X6EV"E'L6AC)Y]C!0 
@O7C\TI_"^*BYY3=)>R]IL*( ;D/$>HMYG;,);R8%>[T 
@05ZM3<*%V;M3B^D.TSEL$+[M>=A6(U<)\5DUF_[&0-D 
@LGLZ64C;8;%T"DAR.MG:77DBRQ)[>#$P:Y-&))G9CET 
@&"5\[3?D+=GQ;4@N_SEHKHPIKT5J:<-)0IUPQTKJ?Z4 
@$"&.XK)6V,8S6[)PR!6YF]89$#<+K]T%/O9CE\DB!O8 
@E6%!'M/S)*D/!>G5ET<J_D7+M&"R;J4'FM>L)&-NNOL 
@K_VQRX*'W58ABK>"AZ,=0M5A^)F'G29+E66[=P4NFX$ 
@L F+._@!5%1+>X,M3+M0B&)Q6.DU7FT@UEH8W-F%IWL 
@]E0S]"(BG!B%_8):QI:SO[.%SI:S($KF0A8<_Q_M"SH 
@3A30XX#+V\Y X4N1\RPKSQEE\C,WX73E<!=XT99#)A4 
@(X.1@L2_F#T2WN"<@,SR%'2<:H7X.GZ1K>B3O%?A\B4 
@#8@J? =I4 "!$07' .89AX909[.+H(7TY4KA2_NV%Y\ 
@F:?L2=9)+DU+CAN<1BG5\''!)\7^GGFI)L6BH4./!Y, 
@Q_!THGE6:O[XP#L><YA3&R[NSPKX0G"XSZ@#S66-5T0 
@92Q@G6L36SZ/PGW1/S?/G(.MCGGMEVCI7$9J49'@K_D 
@W>(E2#VS3YQ04BUJ$F?\^GDS/>8>71Z43=WNK3IU^58 
@.M2O$944<P 5>/?M-WKU;5T@([URW*R3*#^H*\E++9\ 
@KVFWPGV?1=26P0'\W@7E<$!PY#I=!*&L"1(]^@^G6D, 
@)ZU(P&N1'B.M],.BOK0 WSC!6+?V-^NJJ;96I7"UB:T 
@R)>K>%>/@3#M:GK3+Z/L_X A4T70)^\PF+(!?HL[ZYL 
@]E>8Z\=IF]/15'OR$C"8%D\AM('E@F4L.@T%0;O"I#L 
@3MC6>YV,)QNJ01,%E9!$03_YS<DTS5"^(]$_BR3:@=0 
@.&5**E&AK:RI=UL(R@LZV\&U('[!%/!V#-JMA\XFWE, 
@]CY6:!5GY4,>!2@#]U/NSVV ([,C"U$EA7?R/VJ5(8X 
@E^G17Y&4LG[S6I;VB6AA.83EE:M*G\/,]0Q)H6B2BF4 
@T-VV37.,(KN/H0@J4=NA):T$^7QUV>K+$8%X^4>,.CX 
@BO)F-8-<.!TIOM$;BHAQQ8*LM^(U.P,)TMDEH\(U,YT 
@:PUCD'*N\_)+1=I/B@;-<]3?J88\3]6\)SP*'LOK9*( 
@Y9HPHZ#A?FO"]H']YGETM:\XT7]PK!8A5#1^!7KRY<T 
@H8N#%4T#7O61?86&&=[#)X6D )+T^5X@Q@C2?\/3HRL 
@D_52<GOQSZ4']2J=T/#1?_^>A)//-Y[]^&"8U3D$V:0 
@>7;'R+F?3CA+#P-Z;#HN-EPTHFK^$N /I"9=TD <KU$ 
@'Z=[R3R0"+-_8LVE$<S7!0W:C3,&3$CUF=*#N,E8ED0 
@L8Y=LA+86Y[X4/PTKAXH5DM4HM#P1Q!G 6/'?T<2KDH 
@U5;+X9..[ZMP>=_^HX\5 BJ3TD%O\#?5(GM+JV^">#\ 
@W<PP!*U9GXW]%*56(@"\UNK.@+>=;T-$CH5T4RWKH)0 
@/VMRQ_W'NX0*=?8$;XC #HV02T\<OF__S>LVJ (!]'  
@$#P+O%[OIZKP=\BX[N4[,:J('*&F.:(#[$O6N;K4NYP 
@9 PT*DLOCW(&^Z/'H^WCP[2GIE8R)!V&\H19<MYBLXL 
@&%V<#O0ED1@DW4<S+I.2K\EM'']-A1QAJ[>HYA^I1X, 
@*Z.PI.1'WK3#/8W=B#2W()GJ3RF0,_N^]1K]6[ $^/< 
@.]2Z%.K\%M_A!VU%B$6++W]^Z]C.^-,?UNJJ0:.??DH 
@R?T^"(J<+D3;3?Q.!F8"4^T"-'FL[##-L^)Z8SP?6EH 
@,-V#T0?110+2X,8-Q)'7@7(SX:N^2QVYYJT<O+,WFX8 
@VA"$=D=+33@U(-X +OP I6J+$T5X41<CL\URP ]R;XT 
@/B!,Z,)2LVG^94EGK\1J9X>W<.L%*W!YN@TK:5_/="0 
@;TY[>C>-.+_EV%6AM2H)U);7ZJ_.X_T#KA4XI:8(4&8 
@\'+7UB@+<+S&*/82K!& RSPQG%-<K+(5?)FWE=-XVC@ 
@-):Q!/7G@%%Q*SSC(5RV:*+H;H2CI+#TD/N7S%;JGG$ 
@JB&@W&V14\N?/NG,.& AS41>G5/(I2,HQOI^_UJ>2\8 
@1-,)-D?T3C0V$X\-\;4M#*IP@!H$76=TF075 F!I?M, 
@5>2OF?[K2.QT:US<BE\:<D=<*<9/L)<#FI1-1@Q7U]P 
@#YU599X[T"DC=)G?2M62SW6_VK1*'^=27>NF[%> O+, 
@#*#G Q\0SIO]U'57A*HGTB^#)7?AC!9,'E@E:+?C.'@ 
@*R19H+FJPC0:9F;^.>%;;#_O[^@8+(V]C"')JH8Q/U  
@OYID@JK8"SP?77&(F5$QU[8.""?J;4G+_5ZPIHTONW\ 
@O=W*&NO;F<_PU9 A,-EV()],;KL(H.7'.+5I02L+B=X 
@,*;]*'?8,T:\ -7RZXAAS>!8(MKX!!<$$1J44V9DS[8 
@-W@$@A@=JUT/T7.AL@80V"QZ3+32Z7A;UAAD';&;R1X 
@>QJFX/.<!M7R=-9OI@1QDQ8>#\=<%4AU<#,>&%E536@ 
@0H+W9=T3O=Z%BZZJ66QJY@NUI()^IU4_BDB4I.'QBE4 
@_N&6#5K/^B#!NC!P%)>:+8,!PF&!&EWA;@15YS7[/]\ 
@KSAN,_V,(,I$ZPU>QV[??TG@1<F1BP;#H6?^B8[&RG< 
@A&)GV8 $M>HXVW%20_T[=D54[F\:+_IMW8\6%[VBO\8 
@ZN>HD'1%91)G>>G\/I1R61P91FKPCW'+>I3XC[0V8$T 
@F]5O)Y6\(4?&"NS/?6.YPG9L6D6K%0HLD^)BC'-QE20 
@5O^W?M066:967,EDC6C^#@07L-OZ/X%X(&=0:_-.#(\ 
@!3![M#>]WLI1R&NG$#D4#=CX77/JH%&A!OVGH&DR+5@ 
@,= R5_\G=@"\KIT;]*5.38:[%X.NBE!+U)F\>/9])5\ 
@/5@P("\6RR@56AK<U\)3SN*ZB\VTC7^WVG_,>5JPQ-< 
@'Q?UG]^-8'BVX*DIXZHE4UMP\=;N[U>MZ 4CH)X;.,H 
@;X&IGV"CE.$KO1E$;;+\Z@+T]ZRX(K,OP.=IMG;-DV4 
@],+H),%$%T5P'0)9<R6.J!@T1) =68L@>BN;#?PLHG@ 
@^GP#8.&"N 8)$T(EXOXH'<_+YF&N3:.B8>(1ZN 7&XH 
@99BFBQ1.^7FE&]/"KX%;)C48\G6V/6H @,,BW$ZP/\  
@SVJ1;K1+8G,E1<0LM*7TYQ293X<#FG5(OKNM_$"$BT0 
@CC]_LZ*^L#LOXJ(;H)ZVYCCJEG80+!Y^5L'V_D8,7R\ 
@D='E34);G(2PN5>AN!%19>5!P^HIE0@L9AKRB3TK*#< 
@29PU]OL5./F/- Q#4N&<\L?((1>XJ)D+CF:@VIB21.8 
@S?!3C,V>5#_UK%-8XO;9EE3-C6T=(5#<S+Z^J'IO2V< 
@V/H!SAKR3QT?*R2C"::K<Q$-@9!O 3U6$!:.BS;4DT0 
@0Q;H  )IRIBO(U#GNPW! $/IRP2G[D14)/#5<0;4@9P 
@W]KLS:@^ $8;3DH?JV3'FG*-C^426),E)EQ:2X#CGK\ 
@>N]55QW()#/V0(,^XA5W&U/>"J1UR'K ;38QMT\1U[T 
@=TJ<,2O[8>\V7G$=4M6AN27Z&7__RYD-'75T]8\C,O  
@GEE-&>.)K= (N(#2R) !.#$,P=,6L1E9;KWJ4;7A/X$ 
@/M(AT^K]P0$5[34>\C**O$I4AJ1,!![EID&LU0P*Y<D 
@R1D?ZF4MOO/YY&58("00GC'"3<,/,$.;\4))_PA'C?P 
@J$)QB*K?F,6)1:#QQ2\%-8Q .Q#Q4SQ0&8XD5E?HTT  
@\)#5$0DE*<MH,U O26; (A) TW6>$Q,IGKDXUF]TAW< 
@X?ZG_ODDR[W;OFR<EH*0%@":7!9*8$T9%D\DAH^WW@@ 
@5"@U<NYHP(Y[C9+'.T%">%24M31XY>X"?$]0*Z-$YV@ 
@:'QJNP^Y8F9XZ]$9J55Z@&IZ95#5:<E3%QXZAV9 X!, 
@;^6+)\ZH;^)!RBD2+3:]=HZR_E+A]<OUZ#S:D55_(DH 
@_L/D&^VIEC8N(TK]UJ:'3M']Z3)=5M[$)%HPV:L=L]\ 
@$B,@V!+5;#("NUB>R"2&/9;/7V*CCPRB4.OU="L\*QP 
@5RM@%P(9OOYCFT0<KM?<I)5N-@&OOGE6$T,AKB0 ('D 
@["$(UV9O(-B6WLP*W:%K)<+K&?@ P 3I1#"R?5Y#%>( 
@0!S2Y>,7/8#^NR::Z4-P=D8V';X%UD !0<_N$MU4$3( 
@\)DHZ+B"M2) 7VJW6RRECH-XKW#):!6BM;,O_X*]*40 
@L>&T#W]#7[A,%0&XF7@;]"NQC[R;K(N=H_L2X$FW"KL 
@^-'L\.<Y0'GE'=C%[(.48YA6P>_RUSP%FP>_1DLG@(, 
@%&;$5:O:ZU$G'Z/]9%T.K/W/*<[_^@TNK>RY[]D+4&@ 
@]'<H#Q43%FAM:4]&BXD?P7AOV=;+&P+=BB6/NUI!XU4 
@-9-G"3 [B>.Q[/J2]21F&RCA;G/:.6*'O3?V"8:<1*X 
@TJE::^<T+]2VG2AXV7L?_=V/?PR>Q?@O+YXD@$ZC)D8 
@Y_"0IP^N(W9![SLR# -)E^;A[TM[[6E#'B$;<J6V1;  
@\U=*+<;<Z+%$TL>>P-K!#3$F&L![["2R^-6,18MY1XL 
@=)N[CRHX QN;B'!SW82&,E?1P^BL69\YHZCNU+9EJ%  
@L=%3!(XD9>]0(>4TYAO'Q[9HX$6F>T76F)*)CWXJ?AL 
@+ 'CQX&,5'MB\GBB*>)?E4HJ,HZVJRSK)0=HQ4*!QR( 
@LC)QZ>A"$=5A6/L1,S^G0%WQ_@GU_2!PDJYDVU9=]PL 
@Z/IJ'W@+&Q0J1)?>X))-%$C#!=LTF%\.93'^_%6"M"4 
@\A0I=!)?C6ZS0D*Z2I'3NDK*)9]YX6'<.%.CR\HI@=L 
@I#XHT2U_6E0 /US>GG0*OO! &U;U:VRNPB$B@_Z6>K< 
@5W(UM\T%6_)/YDE@ \><X@?]?,<=7SA66'3"(E\KM)@ 
@,0XCP]#SD63^K,>=8%G,8SS^K^.)V$#)^VH OCCJHU\ 
@VA&&W+;$DD)4_3@M57CD?W]]]H UQ7OIN"8BVME^@-8 
@DBLW38T"=[$CQ.ZD@A)$16+E86^F:Y4Q[X"?@5/%-&\ 
@16M^[>L*/U&;QY[A2(_>=PN J7;9$F>[GYO^(/$.6"X 
@F1N^]7/>NOI]Y*D/*[0%.NC^L#N+H&G]#OGE!*J-O\0 
@H\$ZUTU:S(VM'UX>FZ<T!IR1IXNCB:V)MN_!;!3GS?X 
@V/?077C:*,7BF-S;!_S'=D_;C7VN847\F\^UY_QK-*\ 
@?3.K[V4T 0_[S,+.*T9WLMW^[QZR.)74?&8@^ O$/D( 
@@Y:6C+"'!"Y\-6NN"'VX$VR:!2P/> C>-M=_?3YQ*V4 
@F)M=@R.;A*;4M 2372S-X]A*S!G1O]I,NK,;%<IOVG$ 
@A;&":-ZP&P@\D&#_1A<=O+.T:KS@'6L[+!O0ZU#K0AL 
@B X#+HE!N[:CM (T\YAC17<9:@E%$V=&GMI^;1+#%$< 
@WVF]=L>]+HQ;+JO?O=X&G&-H 8(.C&J)"3/H79W2-;X 
@8_#19D\+MLK>^?.L#@:T#AW%J3,0#4B[\AT+#P #[M  
@[46*3-$CD160@7'?Y%#RM11[ Z@XZ$G/#(J/T_TP%UP 
@Z6T)O$4!@=%2'=//T\1)U+>GX0E<S5ZGLM)#K#@MFFP 
@?#8>T&)V/W6:-E3P,?9N.CPR;9%U_R>D>Q2CK?;"HMT 
@9"#_6[PP)E"(IZ;4CBV;R5PALX8KIJZNO4BR(1V^C2X 
@A/6FT?\2N]%@;NLB/,4H:6&/'A34?Q<6":ZUZ%=S?V0 
@52<;M*N'," I'[9R# <$<=V$X822!Y&IJ.8'=5B^*_< 
@0VC,D1O@'#\%S0/7EM]F+RW79_I!X"X$<@E5P29FD@8 
@GH.^Q5*L5 B8_IC*<_LD:W0 6_I,9 Q*: ) QP8X#?, 
@+<CK(<.,L@(=!CI"HW'=9Y^'YJ=EEZC\TA*7: MQEO\ 
@O8@/X"AW*0.2G_";@#6TX>:K$H"SA3K;&BG\:$"/R<$ 
@9E/P>4)))D%"5RQE)9CC\;;^HHBX9F?(@/,;\_P$%>  
@^.6_=YV2T?9;2)?-'\9FW1>2F6G%I7=!MG]#0"2-6J\ 
@4M1WP.E,@P"]YL5D]T$,29OSR\KU& ,CPM=JXK.AAB  
@P) '3<-_>YMZY*?\;8DNE,?9\ W7B'7XTOS5,?$]%O0 
@PE#-"6![E ^;J&>TD14B4N-?)U4WQ_,3N"$-79V4$04 
@5XR('&-B.FE$9&>MM@%-$)7Z-2?,:^,_Q+WJ&=_X!?\ 
@R5&SFTK<<6S,#A^8<8C\@0 ,7<^!"]<3)40A359U8D@ 
@&&.5E>]F[*(*49YB73#F94H.YIAM/&)7;,X3(C(*WP( 
@39$Z>':B290#)73B6>$AK1B)5%R?N%_X\*M:LR.O0H  
@H\/W#/Z6MI]9E-*%H5#\:HQK85?VO+1I%!ULM/>)]/@ 
@*)G2=3>@AV/?R6$F &+>\)7*'QW5\5Y)ICZWX25S>60 
@JP>@0YAI"V4RWS6QIEP?[QD4<PU(OWP ;$BL.9>#)L8 
@:" :_/V-$2P +?,R"NR":.W4"8Z"PH;DY>Q<N [-IE4 
@F@=R[94=6KQ;\ /9\0RU, ]>5GW'4S_]UZ=+O5$FSR\ 
@G EQ@@I7KH+%?!MY-90+ZME!;G(79 )J''O[")^N4_P 
@0-C;3]:V!: TFG2%;O3HW?26K/?_J:R)*BGXH6Y\JE  
@[ZI#*&?M1XE/$:'W"(:-;M5VJ-^=;G&Q[$:=NAGM8$H 
@>KPC/<%+^6\0+=YN1*<28 8HAT4(XGTM'S._CJ>4GJ  
@.H0Q(B!R2?PCO5O.R!">/U^755C*P= ':1;+:W>&::4 
@E=W!B?Q2/D366#L?F6O!'O'.HC7^IJ-I"(IC!,0T2%4 
@A(^:)HHOD7?Y*Q)@4+4_79F)':B'>?YKI@9QW1%RX,T 
@B6R6@98,NZ=5(PN(?52Y487\Z3,#+G^YY4EWWG"M]@$ 
@G'!D3G""XC[5A-;(1;J[#/&%]6$1?(ASX,F-U(A#070 
@9?EIC<18[9@7.CJ9N@CY\\]N4+(9"W)N2Q JVCG:E/@ 
@;5-^;?. @KSTVUH3?1[-!HD4;2Q(;GG"'GM6=^@]4KD 
@9.(AOT:LCX<$FBOR(#KG]M](#$QBZFQ"?;OAXB+UQD8 
@')(KF.^" .8MW6S#P.C=Z2BW&9LOZ,JHUG@KGQ2 !B@ 
@ !USZ2+!D_ O)2^0,=]5/#02<O9NKK-+_ ,T+)DA!U@ 
@4V_@%^H[UAPY>,!*9#HY'4)*RYS\.5U*T;WH\,,'($H 
@GQSF,*Q%!Y]G=;Y+ZN*9^*!JJU574NZX*"?X\(7.8.@ 
@^!XSM)J8*'HQ!62*Q>2G3$!R&YOO(-U=&Y8\Z9<@#QL 
@4]RY,^T =<.6I-H?YR%+/E%XI]RH7R84S>9A-VL3"-L 
@DDO9*=Y#4UN+/#BJ%8H2J+QL*CL(_-<2V=WS#5&>;C@ 
@GQ'?T?'"\QI!2;K'UBN$(T/L?EV6IDBR=3T--2\>JF@ 
@G/44+".A>;C0)\#BM4PGJ5\D1>^I>79BA,<4\*QB4W8 
@J5^7@.:Z,O36[IE9^P 96QSXKW$<$24-V[(2^*\'KA4 
@$EH9?==TU+5I<44.8-OB;LNC,0TB1JFX]T:>*\0]$=P 
@",N8"J04P(L1N^QM.==L&!.,LQC[V]'G(Y1YRNG9!=\ 
@M)14A= >O8!I1,S.+(CBC)\;U.-K1CFZ41430)4@9GH 
@P;9CQK=WN(=S>IDD I!-YYHX D?$W[1R%]5QH0)/@<X 
@<UL4&525?F97F\8,T@C=N1"QWYV=CDQO0<85IC]%@_H 
@G65-^M+.QZ?SQTMI>-$>''GT(P"Q@\>H!*JG>8V&] 4 
@/R1'<O$WE-H?I-*$5&8CTY+[,MK3](A_\I'YV@4;M%D 
@5L=@%IO>O00]Q!]YREB@]8>,ZP%=6^^U'HTK$+:?#HP 
@N:Z *5@Z;KR/(8H#.(6:+UWN_># L+#!8P_.3K$W6^\ 
@369!;A."P76'=I06M%?4H>6(EER1'ZK1TJ'FKHA[N-D 
@3G%HP'_LP2]2\#K16AY-D^N&T(%2SB\R'($HG4L$5-8 
@(^@4\29?(,21:S<@:ZB-'%,[,_@*T R=DH4] D>&8NL 
@#^]^^Q2=>LNDB&KYY''L6H3+COHH-QF$Z@N&J-C5PHL 
@6)+ ]GCWN^6#R*-X$S45/*CC62RF?;;6MF/&VI0:9UH 
@5N*Q[!/#:IH0A4&? -/*W>NJM7X7,_^U5WA0;9C>IF$ 
@M2@1;65[J\44B_:>Q5>'>J.G,]>YG*6,,\3;\WN:=>< 
@3HK=LX;)Q2^Y?)G]Z+\MU]^FV_*2W&GLCP^ _7#$'0L 
@:X'XMU-C>HM4%[\83N#]* W^3#Q=:QL_=_)VI6\A=B, 
@_G,TEK@R%YD%IY&!9%'+-F5H3[,"<5._:@S_19?F1;P 
@&AD*RU6$)/"OM-&@<#DU9JY2X.%H8P(Y.9D!700YAD8 
@(X.:[ 6[Z3_ SH50VG(HPV>[70*L\,41SB95]%WG>=X 
@Z -<?KKO)GX>C1^HV0FDZ$)BZ9>"3$?$G?:^:XTJKM0 
@*&/K'-'@=5:<[56OJZ<'"AEO_VW@90#L38[8"F(? /< 
@[E24)$%V71\*3R#P]-;>&/6)E>,-(M#N"HX-!<:BC'( 
@V#PM+X/92(E,U+B+ FP]>DBL(>#?-'_7(G\[N]NZA]@ 
@?SYO<F9SKF3U[=TP'&!Z;L(<@"(*E";Y9_Q (OTT95\ 
@]"L^1&;0;\6_;&(V_,L;;TC%(48KFL<Q-,RVPD<.4;8 
@F;R_&R'6##(BV[=Y4'0#X[7T'(9R6>)<(P%PK9!+7X$ 
@D^RW;'=$,O2,-U5!Y VV'#T GLD4L'G]@.?,\QC/]E, 
@<. SE .]E(GB2_R#V/RB=(UY\FB%DQAG9Z-<B27(.H, 
@SN,UN1T'RB8?@5I6A2^H<XIE6D\[.C/R&PD)HJ!%(?8 
@&@[CJTVM36<15PQ1PG%W"2("$Q9Y-<1:N]JQ\.@W#?X 
@5AK\NN2ANRC#,SYN&G=<%ND2BNC__C@3 2UU*C?9CD@ 
@>MX"*8V"G<&;KF>IXU)R3?V[MS1\G].L4!;W.:%V7E@ 
@D?_=8YK9I:8L.WI6#:2P['GW;V<[%0?@J2W(\2#Z9 D 
@5"@T^5CGD8,_E$D+.1C9L!_0$$^SU3&-EA$H& !>Z#@ 
@9O#O1=1R1\8%FTT)$*$2M,O/*A[6%=&^Q;7M%]\VDYT 
@'-;1TP@HN24Z5@;H52#UNI)=WXDTW)RZ[+3C1[WR @< 
@N*4*(@0^F*@J;'J5%\7:TM$-0#+@K*;S=.>Q2'P+SF4 
@KP5$,9/%P$U_&T-DC@#'!625R71%$3<(0*4Y!%X'(C< 
@B]<+,:78S_(\7_9A#)#HD%3L"H-'K<$.5K>]L=!S^=8 
@M2;(;R/P$;!C:YZYNVJ'60V7 SDUT/0QBU!D*%,L.1D 
@:W+T0R8#>A]WA#(:I+]WT=A)U\Z/60:!RV_?'/H&.XX 
@UT1)1R>-I?O;H,&:]4%."5?5R=%%Z6#.,M.61Y-^[(0 
@-,C[<:8?NW<6R8X$1'\DT]!R^L=P@[=R4&9AWWL;Q-< 
@;S68:AU=]:_P?^'Q>0(O\MG& ;ATTM5\_8D0^Y-5D-$ 
@22J%II#XA1H*]C;,2H.\X72H:YY>'D3@CF8S7ZP*F2P 
@-LW^H"GQ-WA50E!AT<B61JE1Q<YXN^Q-2:S^%UHQ+5, 
@&POR';ZVS^/NM>^0ONG#0OK+@I.V6KVVO946 ]D6!_4 
@U_ROS6E8RP",$@[@%>/?,BD@U4?MA9Q[H%3K_(RY@00 
@P(7V8K/_EJOP:/N*>+T[-X>-^ )A5 P>R+A\#>N:/=< 
@1!B\*P;1G5\:G[XLOAM@3T$,2,H+&2=QG4!\8JJH6JD 
@S: 32Y9MGK"5>3VD7J>T*68B@G.R4NT,Q,+L0D/];V@ 
@])GRE3SX*^FP)-N*.RSK16/!ZTA>;%6@KTQ6%)E26J( 
@P62<1=!9ODBU"LJGFX(/K&ZITT"L53/RF#V>.M$XF1H 
@"C@".HR[@Q*-*!_? ZZIP I&-\_?3@Y\&%:I Q;CC[< 
@D98NW7,'X?_M.(Y&?91>5.NF1'!1"'C^B,)B82&Q@#4 
@7)IFYL390-NIDYFP;6;=?T585';N@8 8XXY?]0CO34D 
@=N6SS3*W3D4"I$9#+[IO]<\.YW6%$_?2=IA*IPIF&*T 
@3F!EZ KG&[*"YQ)4>XWM=!1 5NEBS';"("LEK1BC#1P 
@$OEZUE0#1'&L=W=?I2<K >YP*OLOOD3FI)!"P^?@/RT 
@5,:1]2'B[S47,1C4^Q ;4*$P4U\H5S_Y;R$U5MB1PJD 
@#S/B@)I!$QE0J[?']IP*[*HW-?>/&1]9^8I[II2X4Q4 
@I96(H3_!@QY1,_(CNB9(+&^36M!@QVF/&M5YSC@;G6\ 
@=D:]<2*>E7D"^-<WVP)M%NX"\W=1OKO1CP4Q*JA74CH 
@<>EQL+-;S AHX#=J\T= Y)C&SDN:Z-W?*BT=KJV-J]T 
@J=P=,F=MH%F!9-*&WTPJ1.W57FT$2LS1^:?C(Q<KUF  
@HNRS8?Z!MND\2[1!B\=3_'V9//"6LD*'UH=![_T\P:( 
@]NT&!B/>3IP)J@VV4%B&J5\_6P  =)_VFMW4[/(=^JX 
@U(*-18+)"&VHCMLF6Q,HQM=)OTETD.Z%6HM([M8_7+T 
@7ZP8/7M9JAE86['BZC<EH<XQ&_ .=:8I/L[XS?>@N?P 
@H7D/N99;[[^VNAI+KW)V,MC4X4?>BC3DS2\0/^RV>/$ 
@7FB7!Q3.\Z;_U5KQ>4#=R,./8M+\2T]W*KP$?BG=-"L 
@_42"/+A*,@[V156#JSI 3,_KP))*!K)AMUS;W&9 B<H 
@ K0]L@+)S%(K_'X2>,QY\Y88Y:U!H1FB&QD8Q_E_5?@ 
@,6VS._G<S>,K<GH:R % X#C[Q>&2Q<WOS:_LD]+I)E\ 
@Y_:@ZR(X//_77!%UZ*'EFM(P" <!<9%P 0'D?]IM@=$ 
@T\[:,_.,#D'"T>J*V^B0=3@<8]/(1]$-L2LQC.3'WFP 
@&6QLJQPR"/(3YG2YZT>ZFZ )_V2D=RKD2U^$:VDBWAL 
@B :\ "TA-'2"1F3[APPA(%4NN_<1?S11V2'*2  6X;L 
@4NU"F9DV)+.# X>3]-@]?=MCKYPNO<.=I)6(L!+QW \ 
@<3N$>EE +U^_T#;-1TG+5!C;F+QC!?"2O'\(.<UK=A4 
@.O/]1Y9WW!&Y2!@M](/72BN8DWO#XYR ZM@<8.B+F'( 
@3T'>&:N]'(3OEJ^R-W3G;$()/(Y8LH2.4F)Y:%O!Y$8 
@U".O*;4D^Z24?!U;#L)+:8Y2%P<RY>UW7OJ77,=&,D  
@-[ODVH=7-W';H(1I9VM_$LG#W*:VBQTW.,OW\ 8!O X 
@M+4WX4Y1L=_[Q09PF2S;Y(3LZM^P^CYT.:0>#.)U/@X 
@YN"'ILDD#7?![SK <!4->Q%/A((!:_:%0,E[MCT),+4 
@\J!$E3B;P@<!E1YM9/U^V+B-'''ST>6H/*$8O30KQC< 
@H8>,9.D2-W*VI!=+M'XX&^44W,":3P;;EKIE'YJJ/L  
@!LF'W'6$,44$B^G2P.95X)*?4<P0$(U7D3]$.>'!R(( 
@C7A[I.CQ;L< ?ZO*%'[49@4*$4-D0$VBKWWZS,PXS?( 
@[/7"^)A/'Y$T_7(>+;N89:^S%)#8CZ1+[Y=;L>;.K_  
@T:6]TI7]B9MZ,D\PM>%YA:O"5;!Y"V8<3I3ZNRK6'4  
@GLC$FOT7;0)5ROTL-$+QV+G\("<,5B^;K7U/J6D'N)H 
@'N ]Y8:_]L1PRMEOZ2CD0"1ZR+OU2M8S!GILFY1\$YL 
@,U\?5XY?+QRYU;6$UGL]W_'(KNQB\?-#3X&>B.LCF7< 
@QK5;*"B*"@$7 "U]"/+[O*X<?V"K0.UST;#"4ZAQ0TH 
@$Z<87[<'\2U%R*&=^S.E%;<W 6O3PU)]0 BO4^,2]6( 
@G50&NL;BA9*ST<FO6#_5,R-[M^61YCH6?!@M*:05N*\ 
@LLVO%C ](XD9E13CPG.?MLNBJZKZXC9M(S[-JS7?K_$ 
@"4)!+[X(3^GT19GMUSY538Y-DW_EQKX.[G7T*O_$V', 
@M?08>UI1V<JLS)=E+!@3RMLK2MIR7/DD:%=@SI*BTU0 
@%.>*)$WP+7FX=]!N9^O%)#"+OAUIV[% MR2T1WQNJ70 
@K>L'"MFW;O2+^@D6\R)^ 2E0@SL_"XT%Q1ZI!=49"\0 
@(U&IM?_=MYNX4I.N@@8 KQT_!GB:>^<RSD ).0B(HT  
@1@I_?G,NUX5N*3&Q^+I<][*WO5Q#.Q(*.ZVB=I17]P\ 
@^5JS!ASZ)''ZZ^AWX-/Q7'+I$:.5V8PDDV?GC:$ZD.D 
@>3MCL7@BV*E5W)YO^ ;:HB-@ 3$9#Q0$=:YX+L_?*1@ 
@78AC)[KC?1EG1?4\])F.NY(OHELWF%GG,B.U91J56%T 
@MATL0ZO7>40A&\EK]F*CQR>^M2F5WU)\PQIPI/^^(*$ 
@J4I:M%M'*T5>9O$5#+HYED-J>440?X)VR=>L*<ETW#H 
@YD/2/BRLS:M.BILJ4'04##KT2X2(J&)OLLWFY-'@*)\ 
@.3[6Z&_?;C[)*BSSFTP%BPM&&GICO10^Y\5_TI%5YCL 
@/*%0ZIYQ43W\9(FN*'(Q?1ERI/BR6_4D,]O<\NXVP_\ 
@"TI'T,[$*7+N,2)LM8,KROJ,!*.=@_/P8HF<N0(9NAP 
@63$8600?U.#2#'!(=9T/(<_P?FTP8:MBR8)U;O7J.VD 
@B^;K"U[N=A-5M@RZ _P5Q.>GPY*+%:R_OBU;PD_$S&X 
@53XI086/ A&EN5Z.QLJ" PREF)E^%&K+"4&CD&#TIY$ 
@FV06_W- <;8O!(L(*'S\@(;RGF]N+RPU/8*MH@WJ^/, 
@\C5S'0>DXHHSZ/Y!YC[[KLW?2B"2\\2JR:+!L-TY$$P 
@!@+S6,EIEOP7HF=BP>8H]_0JM72)Y=)')]&7N''O'8, 
0&: K#Z(_^S%';;9G5K.CIP  
`pragma protect end_protected
