// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Oo8ksNf4lApjzEvlHpJLys45EsrgBtPyXbMwFViZhq64Wffahod1cZyt65BurDMU5wP6Dvbu/aad
wl5l7NbOCehejfLTV2BfPVxG/MKf4IP3e2UGe3CtabIU04+GUcQuaDETugw4K+pSP4+i+Ir3wvm1
tjYr3x9aZrbRdjETntTqoORcmF5zXLYVs3vjSb3VJkxvaxylT98jljVzZA/W/nU0oIGUo2qOhZxi
zpIiXonWWDbBOuqawh9rH74oOfZllG3Bbo9Mfh0a1khJbftD4VUjhFInFjK4qlIQn5lEa1ar5wBg
htT6dsoPsHFLpLjpvN7V0t9BLSvzmQUXU/hxsA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11392)
AaA63ommbGmL5nfTiDvyC+7Qxlhdy9b3t+ekESYMmnjiJDBxxXRvqK0iQFlLWm1ZnnSQBlh/PZAL
WkLwGXPNQnldNKwrMJNxEuI9XFtBaYEczst/pN3oFb7xyinjm/EjwJKyly3lJt/NsbXbl/dA4LWQ
GC8wKbUS66uGbVlwJQD0cqvGRacLRpl+It1FL6eV6KXQE8bJlAD+eeu0+gld4u1P1oEAZIxCkma8
IAYV7omUA+GpV+qDFT3fwQmCmNrIsVZtHb50sUG3tqQZ2HbWQcjLZz01fuN/JZrc1T3Bbp3dQH36
jCsKpm3BbqvBWQt5Rjvm6v4jHyPPx3HaPA2Xf/eM3XNMg/hlNVxsMars54PX3QXmQ3HLX2Qugm0Q
qRL+nmcLMnM0XyU42xEsWhpYs6FWf8svyVWPUb4cxgy8Vrw8KFL2E4Ut4sVVT3FfrSUjV9MVi6ts
MvFfaBsHN8n25vm4sY3E4ZoEmM68E49azrCvoIuOfdLKiz+wW7JNOEhVnASWPiTnEL9/avQ06+0l
XhqaM06wMfdxrR591rBFPdoWw/pmtcfB9E1Nq3HumaH7QiK8Eo8fZ/b0IGd2RhSOifE8b7ijiuMO
359pfMJn0vUWFDYCtxCS6IxMz5aXoI/q9Egkbu3Ok2F/nDaPiuhICV/uuCxMwoTwsIeFxxKEIty5
8V1Wb/9ZoeiEvZ90B6KibqsPyNX6x2Mvbec1SL2ejptwk0LEDDe64Hq9jZYvtOORr4rb+8yuym/W
lZrpDtiBEH3+be4Nc98UdgxGy5qDdcnPQ1miSOuebX1v2uiWaRVs1T3gMMCJRoUAu0tRyjUriSW7
q8vZkvyeGljAzEW/1auoxi3HBY+QJW/czYubx2PqgrIdiicGKthY+NLoT/KVM9Hz4azhjaEXBSkt
qfCKIC0cIe/7xpfu9LtBI5L7LeGTDFlrWqPjaRM3LdCrt+YJsbIlBlB4EecsNaS7pWI1e4/jhLud
oqSbO3QB4xozUS9ju3cskEm03MrQLcZiPL0PNoey/TwnhbSdvB2iyJ2sV1EGW5MuP8y4lLPU2Gz9
nFcCEeOTL4zQZCR3+RuCI/rz7Kuc9U7DXYFED2Tho2lNgs3bzDWBiJ3dyvqdhkhH48cJnP0oZgCt
XF8br6j5XY0WgJAJFvrG0ioszmaB7+bA7VcgL8ZHiWQAuOHZ1Sb2RUkldifNwuQ/VoYknt0UVqKc
bZ4SLlarmVquKTFZ9oKlii+YS8oHeLva9LYdemkgj0tnsYFjKxkjYtbjZvqHYQJpz3B4nsRjOwFo
hLsOc9AytVlCJryBS/9avIX1+qF747DiHMBnKwdvrK3U6Hxv/q+Co3lEQEdF3RWLNZoWRZxvk79I
fYv2CUDK6pW2RHoHtvGm/msJOVNugeTE9dTCR7M6Pgt3LltFZDlQyHJSUKcaiY3z7pNuUvbbe5D0
ZOFSMYspofA8AOzTTpIrmH1f/hC4dS7cmOOIBc8vMFTxm1FHs+S1d0CcKgc9RxoYrr8CJdoFK+BB
nPt8rtOFaratbjpYkcZ7UOxEDpfe/2HN7GwlIIcck8Ac8K1koxswdPnxIAnKd//WoDVIpNStJrQe
1SxH1ydI26USEjBKWNYlGv0iIwvNrSEmFtPsj5DcI56rUotJ0Sz2Ol15UzwtEoX5k8E82Uj1AaSF
tj/X0GzDoHJ+XMW64JMSroX6zQnvVpFErwKlPYZYcXWMjBlTaQR4xvWHGiVbVAskSCSKl1pGHven
15TNWdWk4crFVEKCDXrjncRWBzJCZ70XBYj+RuL7hxKW+2hKKxbmwzx6nf/m4uiNg+8aZQcqi8Rv
U5lkHW3/KIqVmAFB5rAJM9J+pd/EN/0uunf0RGqCmxgyTCwrbgqO1zxyewQNATRSJlJsfseb9kva
kYY87tiu7RxeWf7oNxMPejd4qsApbEOVG2sCb+Y+aXPbxYKkxxItC7CJOyYkt9WevE3XWC73YaXf
ro6RTq09oMzDFgkLjdjlXL5DjIGQdTtyZJ+5FwRZwbCgJY31Gcsp5VX5s/LaU8bqoXe95wP4skwf
AQMhmV7kbT6N2hFnAw3nwOVFWtEwcUHNGSwDBE5dn9a4OXF0jpC6dOHGyC9Zs/ZwjP/GHhMeraIx
DzqSDKWGnAV+6f2LzjexiMmsF2nXp2l2+xSw2CmtQbxPfIPxVxgMw54GR1V7SUxJKrrlrEky020G
SH+0qr9q5DTlFn07kciNQ6wOIbtylmVMwI+0G2rYNV1rNR+7TgVBi5NhzasB7EQyIe70aGWFb+Kb
fDCWQJa/icvnwjnMdVTegCrbTFiH6PiaK1U2Z/LBa7vFj9+UgLzaWc31jWs64IbzUfm5tVfV/qY3
IMoy+1JdmKgtSYHrn3SYmx52ad8xeK9BOFK3dAxFhoFnQT2pbaVnv0+5TyMoVdIbj7YUJi6TrnhV
p2ILONb4wDgfE3+rLUbbdFrfj70+BnpeDWwrOz4tH+F6l6CPUQWpSdn9VY8AnBy+JK/Ev2GGFJZb
qvIqsdOfSCvqPzMPOKXKPhWhXDU6Skfq9WC/z8MZ7N99AEwJVcVWUHF5ChWJ9SB7GsWJNJTX1gpp
IB9CTqtyWXRD/xq7bDJ9pzNlxWCmMet/RF9viIVxqeA2lsYg8ofMhDnMl12qHVOgIovnf+ZQBIeX
bH2wFIXuwhkp7HgAxR3tlt17Nrl8nzGQiFjb38J2/temJBeEZtIhPmAbKj3i2Lsxn+yLk8DeWOJ+
fDpABXN2cv/QdUITouMHGEGAmfM9wPLqc8Z52YgHqRSskD5GFG4DjzBq9X1CXss0HQor/CpEIHDT
XGSQpnW75Isu7bekpfNcut1cvlfTintM9cekJjco8sLIHAdFI+J5JKKGMpKScRwr6rHyExDDCidf
2A2hkPfwDSol9jbsyK8pyxLkaAS8oo0416dPUX9D8p8HlsPUck6a0D3hbDMnlRa6P2yQvrgm/Oj3
/m/sRX/gZUMTY/JsiQp1gHcxmjkTgGhNfOxZfDJGjnkU24+s7UJuBPbok2LZxVXEqbw+weRiYrxm
SOfm/obhb/69qWDMNuAYqg+xGPwQBx8zzvv/tewaYWtradxt6+7hoqivxP0PcIdbce8sOGfPr1uH
/cscVLaqDejgbO5i9e4EdYUImFfRWCYG7RqHrv7bPChiYWn8onUqPd5NAv4HAPokh8Lj7rj8ZKoL
kWFhc4Nul37ZemYBle0Im5V0oldvIUkPqnFc45aKp/MwxGFAf2b/AS2zLG9XQWX3RaUcA5ei6nLF
w7Ahy1fK75y+lmmilpmBMBzLrN5ZFfWD0MS/tp+VQE3i0bFiqYhwA0dKo2c4H4UgQPOiseldFrFu
5CjxeirC578OBWOcKI9pvgFrF14eN838FQ+Jn4n3UF9tTVZDFGJxbvewgedmhj+F6l8YagChIXV4
RuJoUrZl5xoRv9PwyM2qRN8g96WqLtzLCBYSJzqu9oC6oOWtXgGLJd+z7ZWjwNv3j5MAwLpO3+5U
sAMC//1vcz9eafCs1s2335tfmaX8exhOePaFEjMMIvBiCPUnwY5M//nR3rhpjvEcMbuKT2iHotjC
qMa0VDO0V9nM8Jb84XBiVGibslXBvbtWYi4GqZgoh7L/NBAZe1oSTbvUwR7J5rNDAiDHlCdHlY7Z
GC4YdSxFRZ5eMbc4l1yEeMC8HDJVOWHsbU280fkpU+Mtiu5+gOykn0+XHzRQcbzt3cAlulJ7+MAY
YMrNWJrS9OBUZ7z6i589RbWL2t28Ykgun9e3uppz392jrsQ0NR43/kL1AprIeOV5KCylkeDQ06yN
8C76KnX9GBIC0Wc2GwUXISyAomeWSNx75DCy+optoxH7hVOTWyfg83GOWsT+L5yDXrBn56zE5UPj
YC9LgfOYVs89Gkz+ThCWrab5Ogk4XsEsc2kMoX/GzK8as1O2voPRMfXPMhHf4rjR3BKV9JUGIZVJ
w8wRJZYhnkl/hZWRgrMkO1Kp9mOPK0v4AQQbNkVml30zZjMbh1pbo+u5kr0+ufdBkKDa+fZQo4bP
cqv6oD8E/xm9H+IX1KnvuOQrtz/PFujXBWKiMnOD/wKlExR760++FIpX2WggaxvhSwrhNXZOIDRW
DDX7BUlhk0jUTUq2AWF0QdVMugSEOZfuio3wqC6zj379/X+X7eItb8U1HsEZUu46lTS+/ckmfXf9
ImeyxqnoGDZNYOwyAi//t16G9peObvwPxzP8Y7sFTSMO8nKTErY5PDn0pQrdT0PSUdIDktEn7NF3
xUkuu1tL4ObK8jMN0W1SChcefnQ1hO48tS3Flx8IgH/cDLn4d0U1QdsF/JEfoKXiCGwbO9MpIpNQ
4E5lWDVqeV9AuIVH4X/xIGTXDce3ohAASHYWtf5kmRDMn0VTull/UZqcPVXLKCBrrxd6975Fkein
0HusoaZKHgehqUVfMexeZ3mqY04Qzsxi97UXClyYI4HpeK+pKH6eP6lWoAdO5rqaojP+DNeEGj+x
XyjM3tS4PI1hve7fc3Th5LW6Z8zXDTDf7fODEX3f51QzqwNosaleTjwa4Fi6xebgapf03NBk4K5v
ZQXD28uaisQ1vfhrs/4HDxe5p4f+Xi0gMnJwOLCwRp0j9xdOtGq21Xxw5NeBHNg7DkFHaL2Ylu8F
kP2cSkYCFWnBg1jvbs3hemBj6XnEeBKP9A0IUm1lfJ1lZNZGu9v/QNY7OwjzmPzEBG1N8p43pxJQ
YdpEjg+AZq6msQvJF1kwYDJJbhjWi+lHbH6/W/5cWIoJqRpKaJ0T3aKZJv+Qs7MnquCIDbitypK+
MJXsJdLWyfTjDWrCjoVsT65tvLNKugh2pfBANJWKOSyTMY3kPS9sDm1mtHyrCDMPMBFSZxF8d1aa
AJXq4JRXeWO54ku18tH6fWyQw9GVb/0G4TKsuZkahr0ucHrtKtcclkQ47qt9BedjxPmI+8RHYTK8
614a4VKh4mNE7GgEcbxH6tle1cLrqFdf4HwlzVfq4sSlDIYmATCu767P9BqIFvsZXp9zWkyz4J7M
qxm/M46HSqvKGzjxD2hFOh0CKDRAe/uedC76vFIRRRist9fIt0QBPygEEniWOxUa9R6lYnBPpWps
BEF8rEkO0GOaewZkXWtGvr+j6ufCvNgHNYHDK0gcIND09a9L+1WA+6v4iQ2yEpCkHdOzCRWFeLL8
Z8Rq3DtXctlrisUHXxYKox4mg0IaG4ch7rwrtmVi0TlBAzY6hEIKr6iufDC1FBTRhwVm8BNZgsXp
QkpQVOtT0jI4bcHY3CDYcgr68sjqRVcB1ADr+YFNESKK7Unh95tB+/Hf14gOZj+OCbL0naKSi83x
qI/YdEsQzVIjdZhtCUbJIFnxJ08EU6p0000vJO1VEPeoEynuMqLB/ikNV+7SvcjRwfWW8F4oSJew
K990YJRpW7wK00ie/DJ95GZAXPckgm3vZ/C4RFsPfZdcRA0k78Cpr96Hq36QawVpWqoAGAKZtDOP
I2/nR5YrH1j7hqEIerFzBd/gMV1NxJESpiQtXCi3rAqxDofto5vbdPyhgV8uVgFkcH616yJg9z10
jzJorEpdrSBqcUKNk5Y9owkgJ8Mr1xjPEy0k/ofunQcuxF8nAK69Z6BLJDjQ/f7TTBV9eASt0uX4
1+Muk4P0lSVZcfsljA0CzwxbRmaUBYRtYE4kPlXoW6u+vu19zSACoux3s87YetJGpRNJjd33Q8Jb
drCIJ6fh1EJdweGVM2abt5c6O+Uvu7h/qVHmyt5Sq6A6EAlCdwgqm4uDXXs5zUwavMzpdL13/qBP
uc//ZRKh1KeAyhEOd1gtgkF1ToWkD0dxctmrK1MWh175MSuYyYXjd7V8r15vGgPunbT5lpDUnZxV
8f9JHJLdKH8Pt6MoXzA4bGRtWF6GPNXCS8wzrB0CCrOv3R4KS5e5grf2s7U5q2bLynMmmFGwP6nF
iZwTBzldx+JLbBOBrSTffVl1hH/Ma3nPYgsnq7AzJUZ00Jgbu0l65wxfbAMgsdJdmTnkCr2Qd+3O
l7RcXN2ff3hHNntMmT1AFe5q+xbpDNMBaHo6CzRm+hzt5o64Og86slliV/sMA4Z2xgejqkE2s1N6
DYV1qYJuhIBRKZ0sQpQmfZO0SkTFopLI+HNj3qpPtBd4/nTMsv61yBJ5/BJLHoP7dSNdPag8kEy2
dQB5zax3l9Oe7UnjcExlkmDnA9PrSIPP0u6Qlzj9CFH9jSj0Eh++joZYyWBeK10SYa/k+A+0zHrx
AGa/e7YH8YPj/7q4WKEny9JkAkZUWdM6qy7O0KlCedpcLf2vc7m7CwqHTbvazKxwXu31MvS8cwNm
YLyrR7UvNF0ENGrxJJposDx6ji44k4g8zxcSlz1m8yAL1YLqAN17NbS0IOK0UUVb5C5YC/sGemUP
tdoDfiFpjFncEXPkEVt3oiaX1PsCb55R2McJ8UdI2+uGhrCfEcbj0rvLGKpyuixog3ZJg5MBgYmB
GK1Zc7huvv8kATuK4QOgJFJzShWPEcYjo5era7uyKC7LN6p+U6vHX7BEnOzbVtbVahR0YzZweZK4
VYiNgkfx58nkWl0VNru2DXFUnIR6Axe9i5yr5aCJmOA0cbQubIlcx23sdfFVwddgY3bGhsQFu3mS
TWHjaZi1ppm272vMzTcu9qePP0u7eNmpiF1CDbw7zROvh+RcpQCJiJMkVe3ZmBfRUiYtCr9qlDvl
RKzM68nHujmLZG4c7OdKJmtHy5JDwAlcRx/CE5acx3iyGnx0lRSLnpiJRx2p0SQvuR8m0SyJbuFZ
ihPDr0t3iST90kOB6Iwdz1G6woAioViF69E5RUDNFWCv3o6+gkk/YwZOYOXcTBzCTSPc2VmUF0Jd
cosep9gsHRp1NM/sfKOPK7T37Eec9KgcvdfKYoqMfSg+MAZdwZqPfeFDgljU7Kz/lGoTFil/71TX
DGMjB+TjlqGCyPOH8EbdEvUzVoltOsmlzLttr5ZNZ0GKqH0nQqM8LYKhu2TS5vJBeJrT3H1Z/7Xq
4oqUxf8/H/Tv2wJXrggutBR/6upCb3E2F40ZRevragLK1tysoTjGPNcbQhHIMNmdLN8JN7p1z6JB
tD6xQE9btd1QpEudpQqDBvdVKBsq449eMrcW2HPX9L1yt0+pMX8y9LmO5JWLORFOLDmtxkRdyXhF
8ES8dHse/f5l8PckeFZKdLjedAS6LOxfBreVncYrzun3x6l8C2zwaPuqFOGuMhw7G7hHd3Sgowgk
lzxo5qwAgBVfwtmBtcuzQzIHrshp7DotNaav6LG5Hr0RgaB6TZzY7Ky+GhZPh9/OWVbJ/chjyJEm
Cm8PsK5yRItOkkGudEmwDXGhud2LmMzJR6DW85fpV+kYYHCnnE70Fk4KyRgUAFXytQSR++iIu/Q/
UYpby08XBQL+QylLzj4zKAxdKwcUbo0T5YHtptbApHmSUA0olhntuSmchapIFz15YQOrtJbGdvKu
V9aD8OxDHNztnDZCaF9Kj9ZupWC02v6HwnXBJxaxC2D/D8gl6KXUxQ7zThyYnGdRdRXcSTqNuNOk
AoklIIkR3v+W/kZDiCwE1f/7h0uPEcBztFWbJHu67olZ/+Gdj2T91VwMebN1Lgo7PrKY/lhn9F1o
vQigCPKVazeV4ZO820cQ/sxXCl19OHN45vbuyRbmHEAU82URgO97G2V8ThofTCiDy/UkQq3BYluF
NOH9lHvKZyZy1/6zXEZjwXf9X1Diht4EgQ9ntpwSODIUmsGdNsIiqjUTOHB3AnOLDcAVI8fKAgt3
ZiyoaPljCSDMHu31MMyxdXr8UFdltRHiDJP/+PoNbwCHq42sSN1RBFGUEwh/d2PNoVcvt+cGzwqw
xSLNW5/azO20bMobbdGYWPEC2olnEUV31j7Ujrj9c/sSgtR4pk+eXtJ2a7ITuuL4kwgR5kpaiDeL
KU9lG0lgxccVpr3zleRfDqxIELJvSKpUQ9EQ3+tNziHkmx56mt+Np3SVxWzwsHuyL5o3q/qhuW0p
vSaBpPVHeSDJEdN8Gmyzx9OOzhDYOYaXj2HSZsw6w6IGNuOyKB4KP33dyHrD+D8WZI1wzfhEOKoC
LV53WHsAhYnnY2o55zy4is/Eoa6Ktjq4lQO8jsAVsdcr6vEd4z74gaDtauSIHlkhwTwIvSzHchZo
rbLNu/gblj4qnOo4lI4i4/DOuw1fbL5YyEnIpxYV9ESPCcdU74788QrmN2vdUR+I2WIeZmnc9nFB
6ucS1/GJWGaYrWjXqxQCOArkDgftbzHTu1F8RfoS7D8/3eaO66Foib60xGrh3IaalkzheXXDr1Tc
T9umoTXYvo0Yr+Z0T+Wbu4TENs9E1856ZGczH/Rozjw3CKAyWqxvgR9neSug9SPhR3QbyWLW6zuo
LfNk8rFLP0mhAsyL2U2pXgIVY3dTtNSKb+0PraN5IuUn5hve2rVOysdXZDpAuM94jkhkFNSwW8Q9
hjIrWxVgQY/wYPHp0o02xxKCEm1G7b9yCUXbD0RRArBv3500Y/eyCFh6MOFTCoSC5wX27VUaVNTm
mAh5NGsrG+ro3ym6a6TMcq/Zp4BH5ZbNkXCpD3ZhBihrREhifMY27f/1P29hEiF7RvnNK7TqDZbP
c4KWpsJkiiJsLNq0BgT6q8Y+NvF4zVjDlk9ScrAKl9iu9hCP2vnGNbj6VThtdGneoEDVu8JlRG31
BdsMM07SKNPEdu+xhvwXA+xdQrBmo0js9R5ZOBElOw5KuSrJMztYLh+FGW2ei1yDEWSlyY3RmYYS
gEptroGOQvaa+tk5QYV0XVpilyMksArJHhTVZAJ6FXINDt+R/8uax/dEKEPs+9UGQR+xz0VPtSyW
J/IeosNjfiHTOKvJrVBgopBCrsmxbeY68mGgOb1WdsE3IMFbb5Lru3zoQGWdQCHafBsBlDnkcpcF
WIXUGN0S1Nz6k9S2MD+2zVBwJ0aFuIEJOIqv9t96YF9Y4PLKhgcpqmLc7UjnaqPQUI+DJES0Q11e
9qqJhgtYbq6GTGXB5TtMWyvopp0798T9cF0XCp66QL7ypnszZ1WsDF19qE5vlmH9z6XFhG6vDIQ8
vj0nIWcv3I4M/R+PSMRE16wSCvqCjZDT1CUa2plBBg7s4i6k8cl1k9zTWgFU/yoHwKHxmTzu1Ey/
CUMMG8+P+3wkNz0WX5ETbCKCclXk+crBMZoHVDyedYhrZYq4AZwt3CGUjxUht4O3Yc57RIW/ae91
JKWUIPCU0/rJaUDVfyYVOWYdUTZY6B5xWZVjccsW1xSgZ2oWMvGa1rjmrH9PpY1d1Ww4ulIhiU5S
7tEdfZuujgfdEANMcsjLloohqUB2U1dqYeXenyFLGc9q1R5q9pLMn7mF2D/4H7hlv+HXYnZf2etW
ZwoCmcXR+/4hlUL3Auvsu3un/uXd9w3dzSWxTF7NdZti2gd5WBy9s0EORnufGM8FNgm6gCHP6GMG
u8+LdkTlVa8RROsdDxjVkrOaqaWvYohv6/dbpBP+SYTk9LgfPPB+SVshyxa2LqbLv/hU2YejQ2rA
XTWLIXdUYBezOpn2t//DWUu28m+LvlJsVqRYpTHj+7IafS+jWdDt0jYRrSh5vx/vHqvW+YANOQhk
09mrPpkh/tV9GW3bKjU+AlMpwGdo2Rv3A53RsgadkucjsejMqhGLgQJZPbBseaCCFKmHT8U3qqze
W6/W6gh08MFQBJdDzaIHD/KUOOHa02c6schAjRtZprG9jatw4c1fj7kSBIoKtfPtGiXtlke3T5/V
fiwAPOxZrK8w1t/vJYb2GDql9Spfy6YYh7Wbo3D7yxSYnyeuhSFAQyF73mjbW13cYMdTdu4ZiPPm
zxGyUr/3F1w3OHP5pUq5dO0J7EjTVY0AP7c2VjSSydRjHsPzabGlD+LCFdYJNzwMUzgKCT/1PwGP
YyAlS9jS1GvkhC//PGVCMoDzu4GlVNZpZvKE3vXDvIxHzBWhfMZYsY9pCOTdwQR73XifoknV955J
Ns0dxSM+GSb8zeKSFzBbEtfFQSVnFiDUVNZ39YQj01tR5ynx/p1vWOF3yKQWrspmGGbKsVkUh9p0
cAEhZW3xFZqTJT4dOVd77bAMWj/MBgu0BUEtQwxh5Pq5y/7Q2f7OK2DL9M3TFzO/icI/5ovnUYvW
fVueqUMbCniu5mQtupUNIa1EUXTbyw+6+IxrIBFvtOv3XIFb4WweK+/m+c6xm9DQ5tq+8zkDWWV7
LB6c9TXsx5fafNLFnRzSf7W5gAn08WrEiLwlpsFex6rZXf+U/arn6kIzX8FGriFe4NP34CAa18TE
4PAj65NK6LvNoTifwt7bBXP/LVTnNqHMMT6r4RP2Cb1SMKFSJ8i68Vn6T08P0nvch8Qik3wyBp2l
6miDQqE7hUrHpEL6K1v4gKdsRg8qmuP+H6W7Pg38eUoO/ui5sem7a4SMyIZSkzBEsowujIgnCF/b
YAUuYQyBpX9T4K9YeGruGv7kc1fklccEdz220LV42ELT7mpoPrOmbwuMizgEbNEuyj4wXceHBpUA
5qd2xd/siDbeehIwTA9vtK3CGFQq84q0yJ/aewiSieIITlBXmMa+vFilRtCLWK7RMdsIG0TLTvq6
3CUA9+Zb5CJmJ83z1c/MTpha3Ndy/XiORHjrYeq6Fq/eugM5Aop6rHR+ESj++eEioCW7W+qhABbw
joV56n+D6SYWpdasP3clyY/RMycCW84H+uNgjmHXFm3CJh7j0SrWJDWFz5K4r5zVFLBRjSSj8bow
8TseEp0Rf/+YRg+0gbWO0TsOeEOF3k+NbUxMyzpGohLoCiCX43TcvR4PAd9pCW0tDtnxqOXlvKdx
q/DJt5ptZh7A98MGvnNt4F/flecsAZRqJ+hjpTnLZszVQRjhkuNyDSkmepnDoV2SVB8hkNNfFf7Y
DZ2uKleAljByqVMmAfzEkAKzJp4D09CWG6H90cx0LM3IZvJrk4wQy73WCoXjnUPou79f9GvtkYsf
u3EWtu+w55xFQOBYJof2wmVUpIkzuRaEftv5UtEu2fWU10HIM8nrB6qJR/PXExndv2kZC4kI4ug2
2bWyfVBTxku6MyQwavydvZ81b1mmQSzCtJ01TXOcKyGqRsykE/T1Kih4gfbRPzIgCkr31qCh2dRh
sluLIgspkqLiBLazaxjCvK08Q1A8QR4sd8u9LXvrbUpEbL/edLlnVAAncyv5hNxT5Hj6HptbbJrZ
wYuvzNdhS2fNY+uFsFyJ7cHSzB4BYYY+C53Ok0DKJ312udi5/ay5L51f+LxrjLctzce8DZ45nE5+
GHXm1W7TO0yVXq1nEvknbGKBVsoqUpU75eavNiXn79ISI5jNh3Wvh7W/p6DZn88C9AOlDzxAt5q3
8mEOQXuBZ1IPy67iO40xJZp2GHe0AUHgTtT5i/hCzZJ1bphTrNze6FH1YKS3c4WA3IJvtwzLnzHa
M2gsokEY3Y9saBQZHNlKuytdNcK4vzRsFRjJJ81ICFY6UEo6ekjbNmZnhzDbRwcFweYUHgnc25AN
1iF93304HVzINMCYd1s/GKKQnDaf4AI7/JI/A56nN1q7T+gQlAR8tqOJNIWvh4ejrwyTTVGVISDj
WOlVTsredV83Hx/zhkOB6ZtkEQin6ZQBPGmOzQ2eexjPF5hIfYOwaiWFfM44uwzPuVj65FkxXU3p
2gJemL4Wj09jQdvz5Ee64frm5VO2r07R8/6c0K9Q0BhuOBHrN+kjcVeUGRUgIceEzRSPHsLmINuO
YUpLNKth761PCeAkG6TKfVMFeKWj+SW1rInM43zFTAFmhR1pavfGryC8d2MmfQFWlQgaUm3Ktn18
nA6W+N2wi9spotg411z4x3B5XfeaIYPE5H46yeBJtR0pMnsk91jwmKwU3xLA9MPqTUpyK7wxguxk
C5lq9Z7bY1Ch+BF7qEZZQLeAzQXdIWgA9Heq6dx9m09eZdg3+ihq7mteJZ7a1DEsEOyN96I9LpRj
t8lHyWcNBvtqaP9xL+kFlGWeQmx9MW9nPgxIRCN0XCLCoqRn5ncmnvb0g7OJYxCOUq/rhp8FwCC8
PxSDeYMCcEJC6lVa2DGxmVcN0CwgXjqdfPZhOrkHVS7P2VkY0Dpfj06XVDJsHeoDTjrptlpRGBRO
C/BiqjIH0pYY5phzwLZYRfyRlsWP3vccfMT9Zx8aihexxQN16zKJ5FojgFdutiYQT17/ACQFn3kp
MWR/FOKz8ewDumwj/q4Q3+02y8jLrGnQzJZv9WiwjF9iHxgZkXwQygDP+83sJnna5Kgo49+JjzlU
6qFAGAYzxSIJ+J9OSxBQq/OX9pyBs+x2WjyQZHdh7nfLol07LGeoijmme7TWkzpuwtLPp1wHVhga
81mN5nWlQDDdEeLjLAmGFVU9R9tuh0zhKkmW43nj6816C1zG/OLvoh46l64DuX0aMP9VG5O+IQIi
ZI5MNZ8O9M53UxE9+/0ifYZRZvgLWilM50lXcJPkZhQNoYnMfMDUhb7H0JtiHRUFtIFVFapFHwHD
0g9MJRSQRXLwSEl88Pl9+/ncg6KpcO7oE5uIPu1suZU3L9dZkgWjvVmg/W94oogESmGx8wR5GqLi
dIVSD6jHKDUj0HkxxUWZe6WiU/OW4XNhFxbq4E8nthSDG69UKWOZw91OOCS/AR/cWUDpu/wu2rK8
P7l43mCI2O1UUfTUyoKJJ50adyJ0DF5qEct5qzO3C2tBG21CLISonYzXmB2ke/kQ4NjQKD6K5Itg
ywvCE295G1FxBySTcTXG8noASRcl80OBHoAXnPk+OaKOUwcNlnfaWP1SWVP1DtCJlLX0/Mx+MhkZ
OmFAjuTTNy3CO62gH8nzHvTsBurMNY2kvYi68cZuEYSFM+tGLbmkXu6fBalOENSvJTgtGEiNGNUG
yMjsiXkBBPEHrvweDy616ju1cP6R/wOqV+DgoZQhD56v0/7AHPCveY0zyvChaqveG4mLae+lcpIw
EoV2Xlbq69PsaL5Y/72xPYeQm5l1iDPb6MFa6c0B/GsPbCODMFGsMQRXBMfCVyZ/EDf5HpP8kLqn
+yo58NDz0DMrIBkRuhN9MSl16eCe9OdOHdZ3tin3LRRk8rdrb9jZfT56pUkHyHHkeJqALqkKjEh1
vt/jDykNK0aOuORj5T77I+u+0DYPduBNNuTMMUqNUM41zcF33/p+ivtKmdBWYps+qb5ky8SllBsC
K6IEpVZYIFyRNYFYqPvOgeCppOo+Tc8Ez/Ynx52AT8lAHZXPuOs5aD6VTNp2xWm9ZjTcv1euFaMv
EHowmBNDPvX4P8K/+3pyU1vM1syX6YXiDUe8/j9Tz21+kERXnOTA0m3MSXCkMJso2S/r6QBNnyjI
/YZSwtpx3ziybIY8SjPLTeewbTwVWpEeWg7pH7Y8ju96cI8LD9JJVoUa/I5rhPP6RypTOc/gpluJ
Sy4Hm9MXodrEyBoYPSIFiO6sAulvGTlVigdc8SkhaVbs3aP8Me6+0YQXXHnJaEpXXzbhvuTKkx73
st/ZxdKP1ZuKcOgyjt9pNsmtHI2oQmauNrsAhZQ1/u10FmrKM2scRdCGMx2yyyYKAnvE8csr28xr
ox6SZSmzSZGNKmaMMvh0901sATqw+CFZaqFOS8+4BYhvDtMOhALz04m1z/WVZXlQX4Z0QofVfHaN
6vFZXgHf82XTDSdQghc+PVOPDW85NdUUhEpV0xwPpvgxSzphIJC9vqdz7dTirWojJOrM07Thu2hp
r9L/DCeTsBGa4RwLDsO/6cKsGJNJ9zUmW9Vykilk2+Me7bsQhz9G9NndkObjVIjv6FZQe7+Ymbwe
+l0bJbzYJtJdI062RNcOSv2msfSAIUkF5WvJzuQsqIa1yWcPazbLOiTIEjD83TEKUuU2dtWESiMI
eVZArTCV2H+EsvsTRsQEQ4acvKXH/YjT58yPeCNA4rHE+Uuh/dnXUP3xRuJeEc3+7dOJKs9KCkxB
mWO3mZl3p9qE2rGc9LJok0n8bWyY2uU5UjqBlKkWD62bfLOY+z1hsXrpl8H8Z1mCOxzIBXjwgEmo
rj64kMYlQVS5vi7+aNetrSvSM/IFYmH+G7VZrkgVG4aRALYzLL9pLPpJxnEIA2Fivjdzy4QQMD3B
Ke8iSXZvnCvVM8bt3vO78AoAavEFkm0vl+p8gUXNpLJc07/505Uc2aV2wDWI4E0UlDrvTi6SYJfd
wB//dA7fjkCR7UXqKkrwsl29PfEbF51yGcmhfDLcuejuGOBNaacln46zZAunGSvHtnzh5uUobswO
3CSgT6NWqbNsAluBkgxVPBRCpLpy07vkfg5daHzrnukgstdvpeLrJyUECtuXxjepWQQM5Lm8NYxA
l/bZaQC8vhExr49QhO63R5m5FYYNWUDA2Lu1l+0oWP/pAAKEEJIgPDrQmP/GiwKArX6v77ENJ0ZZ
Na5FqwfrzaynNuFaZSXb7U8VMOjuBY7ol/K1LIzzSKt78qe92KMpDLwqYx1mq96hYDTnFGM9VWgt
AtOcHBqsdhk5l0Adjjhs0rBEljjUTc1JRfsgRw3qqQE0wNDLjpXGpTu0UtQdYyCrrXaG2PR4kBcb
z0gmrWA6I+saU+Oxsx4FYekMrHam7/PxQSRlKFeqNmuRC0qKUDlO2wb0faLGXZBrqiGOCoU0Wqm0
lXFmX9jmdVNH7oB7beMY7G0s8p9CeSMG2RsUUWyP4iSl8b31aigQ8G5lLSSt1MmVBAtuku08G63r
mhzeq92bZX77M7NaFTqP3UGJHbRzR6OLB+ti0ZqWNZog8/oSNov2Y5Fakp10u3cltQ5BjgMQWfPs
QiPLbpPoPx5L5JhZlCrRtmLpLrWAjdVG2UfhHpcYroc0HDiGhq0A2dG9DbovEzIcWxdms5GpCW0I
AIQEObVIdgZLcpSR6vxthMIdyQOSQdTx7Ned3IghSG8u9lrloOLQVVR/ZS0XooizShtWhRFSOWni
2kJPl6znw6KKS014BjAeHsnj3JWyzo1P723EY6HO5pkmvzZh0clV9CKPyFvsImbKSi4C0r5DbnFp
jgAo+SCWrRWHEv1TkxpokCkzsfZ91PTBb3W641Yzb9UbVfNAsT2Wx+OdrIak8R+y9o0psRoMXnwD
CXrOfveH0H1ELc/d2iwKuAF09ogKshA1fYrX7oWJ/QXMf5oIQpDJFifoz4IlzLE8cMKucauvH7Tf
1BO9K8W20B/p/BtIxyXXJxiPaaZwq1OI+bJL2gPIS/p1rpHaNdNgaotTHUUwWoZWEA==
`pragma protect end_protected
