// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zz8sp3NcbyiPf8UEYoahop0SkDY9HGr4sGeVuu3O881ZVwYFjW3XtSuzJpXDrvG7
6hzg6hxbYkflV/PINw652ECqnqbW0q3+vh27Lim1zq3gpBBqNCO1XF1SZKmTb0zt
iwJbQPZWdsry0Z1vln7pfVxJFqBQsBed15APLSAuswE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3344)
+pXY0tfVvBSJbYpIOj3rcrMn7w7bS19PSMWyEqsDensaCnU1pUL92SHfl2sjhegU
5kiKhuxv8MXXyeWrnXCX9mQaMCODMcwBtNmHcaalKI6Idt2b2ilG86MqqCwlFhWE
QgxGMBSo7koXcs8ydN8Q9q6wzayZower4RAYQXfC7C1XNM6Lzh5ykHiI3CZcQ2uR
7Lc0b29vWsrL+LhL1vIfKtWTSUIjwdZ9DCve6chzza5RgXbYwyUS5/ZgYAg9/ZwG
B6QUhW7VgDOJ9C6LUMf1XfuGMmZ9URYYkpSJyXO8sVrE98l+Bk+C2Y38lzsu0gnd
beaeg/HdsZ79mISQecp98SYhwSA0hwW6pYItmfasOadLb+5b4Fqt2XA/XuZJoHbk
A7DhsUoB3JeG5D+JzTyurt/NIcXF5N0Xjizyhye3M6mbpsi0YSxPG3qEbd/cZ4VV
4n/PGVmoaq7kdoPG4hhKMbXuUjEPalc9+AgOdbZf0AipqudTeE6otUoXeDAv87Yw
aPn3JGoIjD0X5iy38WzQyVFgt5g5l17hkpSHD5qIaxnFObyqQ4oa/PkDtIdA0a1T
kt1YrzN67+g6R+LQy174dtKiq2xZXGoC4h4CwXC3QkiqX6TZuDKvXfR+XC+nIOh+
t1I1fO2i6OyqmkLxCRrgB8b1sgVq1CL4HfrLF+5THsvD7dK6jyERQRO1emDgzziV
+GzKFg2YYQE/Nf7t188P08JpCq/u6MUz85Ut5gEfiTyb0rKpDmPkz0ny937xwa2e
JgH/fDPr09E3K18atSNT4PdG6eEb8Vjs+MeldXs8Z+3Pl3YyL/XPKluPxQ7vorFB
oYRztxqBOMqys9qRQmUIDWriUcd6F6sIxHOyQ1pM9gJZiZJgnXcaUoGNmMql7tjU
zvuvNnCB5wpcnu7OUdL8ZCDqaw/xQWQdjriK/QhseKn7LELD/zh/HWfzvXUA8sQ/
D+2pHU1/uoZ9J7t0lwfkXHgcj90QotV1GEE5zaPm/DKpn0qa+t/0cQe5f41t/Q0i
MvP9JtME9NZZa83OqqYLe3C6qMtfQrx/ymy9OgefIX+lu2tKuppvWsp9Ff3usToY
JW0JoYnSNq/jwXqs3nlPerWFCsDAajBjlRzc0qoOvXU9p6FhpV4BJQu75GwN2KBX
Sq3GAjrOUoaG84MeZ88x7D9qExiIdF6TgPIEcM30ATLe4oe5XjAVb0L8fGUptLkw
UcpijfSYyk69vNkM5vdb+C6mNHPho6rfKlkr1WigaVmYUkIy/dpKWf8+QMeu+ytj
nRn9dwRK/qFY82avhq/VBojSCvgCpKwHnYe9xE5DkzlLI2FpyMMooLk4Yh2xvoIw
+DefjSbc+BOXz2e7q4+1zohDFpBrgYl+bJuRolMLC1nMupIn2DxLIDcYODBqGDPl
uYzTW5YD/hvSAgt17YNXPZJwBOmEqV9czzI0n+yZINwsUTlLcG7xMaQ65a9JvtpL
2378tx6Ye1ExzFkmutq77fxRr8y4RnFdQpOcQk01wsMRDZn9id/XniwTFiUmAREo
LInPZFo4eOZSXBmgtdhJ+vl505XGv5Cusve7A6qMDSGlmfN51Ku9bTH7hph2LOZT
08yHbX5EbBGzrmL4u6KYEqef9V2uTXDnnzu/4P5/3blURY7MJGNvWv+k7u2Op7DV
Uj6UsGmlDSQgXWhX/VqaIXtTJp35oE4zQ1P65f1/J6JguuWxpYjwr7Vt6KjkTuQ/
DL6GVh97lcDhd42PtZUEVMzZ+GyJoj3JywLL/VxuVcCL5Rr7ZWXxLG+I0p8OXIi2
qfU8nzVBsMeWR5CyRMIhe9mO7M6TmeONGMqqDUdjoxirYiPnf5YEpy45MIRXD8TM
zFxVGxshxSiLWM3oMRl09t3dpouIy/Q8HVTAjzULVsIOH186a/cscAAaC5ME+PLI
u2yhwSg+eW+UUmOzAyJAgaZe6R+gzgfGiRxKF4LsrTs9DtsW46bEpoi3TFpcoOnO
oBnIGlFXL/nXrkvdjeoo+7w9LTzh6RxTqkVw6xGhMNcWIdAPNFblM3PfIBNdZq9L
Hr3AtcZIPn1Eb0dgYDHpWYWrNfr8x2hm1rHINJ7vFW9UwxEO0dSVV1JbL34REUDN
AOYQ6FgiIVauPLH5aBfdJKShNU4Nnps/nPzNOOC+NjmFXO7Tx8UVjSQxoZujte+O
kZc/tZylLf6WZn3Gga/QbEcJLt7YS+96wCRIJ25TwMjDirgLNLuc3JV3qZZloWs+
hL6Kg+D26RS85TPlOi5cR8SyI/nOLQ3gKz1Y4v1aobCUKQRqjHgHNYsljA7v7RL+
L89Bcac2dyCogTsluQLCz0SnOYjv1bNEWURwHKv7mRwd5rawGbGLZugNBtl0uTGA
c7HiLqbzaqOvUYJpr0rYVhb58ScbhWpEd/DI+GtXdVPYObpf9fYb5202Qo/VzaCh
nQzd4flgqvlqXJtmKsnkataXgmM6ZB/geVSaOVzWz4C0A4iPVkriN8WecisYehba
9q20RFvgXZX7OWofyY//IW3DfnWYopD6JXZRCSEn9PD4EZVnRl54Uxd+BT7AOVyt
3lzaCt23OVmyugg7R+0ufcpaDN8M/nhF9jnuT09ekx4oZZ/nitPhEtymuw7NGihH
LqsOpPLlr2YGwUVBYNwtlZYLRQpf61DeAGbuPUa++aR1c5TV6n8moDShbiFoMObg
BOO+e8l6nXkqX5qOdLeh0NhJoihLS6uOuB/dUrVyq+xOgJ5ObjqKZ/lZGuKFcmi5
6g484fye3Gi+SrJGmuZW3xz8k1wmgZhELNi4WLyooMKQVt9UwG9SdplwefEi4G0G
Vsa4rA241q9R7RkJ1HN029OVC4xeyv+n11lPW9DpXAonllBqDw8IHjk+20fyGZGM
uMCCcZZdBRbvK6Su+tCGVUqShONXY7nhwA3/X6RUeCwjztOoEoYstghPiag1LRUP
57tAuFE7yk5foXsfq4bfY2rhhiCYJLTDO0QFQiuPJbluzidE/qRjkfEblhmZmPpQ
0yjnRgJTyqEUpHLRw6Naj+A2wlB4CeI1FdSvomk6yfDD2Z3BCH4kaTO+RnMWFoK8
6yPp4nhBOSNEsVZYNnRp8EEg0LN79/Nk/t1nX7siWfa7fD5ZcnruB/wamPk4mW9B
8AqrQTsH0MSLAtAOkVkxBNZLUNdHyeyBz6lt+yb4LujlyiAmzElPsVoDkRde/gWG
Kr8ZhDaz+HZomGfpaXtv+zhvOaEnukDRR8EFZ+Ck5nuJKYfmAE5XJ3AupBOgLSnu
T4rU/iJu0rviRdiohIegFVJ8Lh+2RU4Gry6TCq6LbuMK3l1ONOy65vc4YLYmadEy
JxKfGzqKGwcaemQaE0O1eC50pNITX9IRv9B+XiBKEQl1SgQMHfGnVct5gb3tnAhJ
S8ewNwXmKPKSa0X+JQffixN5DiFeS2svN/p22ukBkzjXTL6DSjfv5krfZP5q8pnf
LrvSKiu+VCjlnpCzmUUcyDC7oUNzesujb5MIIpyYUqTd6gDquMI5csMM3SNmLP1L
9oJI6mmqLebHXXL6jMyV8OwBvx5UKDfZMu2lckrV1jfn7xEUVU+xB6ZTQW+93XQJ
4KA9MkkVt9TMNRwV19ltwypwHkjlKwzaiM5rhEa0Pa4RTkVSwoUgIsVoWse4zjVB
/q4DzIsrvbyUO+IedqCIw7ZUfSALmrOHKiBS5CqpXKSguNB2tl2SYD9A3C7tL2M7
puvpnoFLKu+x/igIO1OBYBGkOjqm9COV0lXRA/ocqcupeM+BmPJ87g+Jf+r35rsQ
6nkZfdCLGOumSxoTxUVLp/tGJJ9Mg+zcV94BMHm+kxHZ2408noOMIoB/sseORVMr
kJXKT1CNZaJTqRAFUK95+5ZWtTInHGadcWx5QBr2jcZtV23Ensk3IVOFQrJBFctv
EiID17nFku1CAqUe6NARgSONv1LQTjPImDlaA/tTmLxULHvoZ9a7HTeDezXaqOS1
gCIFTw2yCI8SSIe6NPM7Nq39h0VoSvk76SKoqAcS9m12qDPomJQiU6A4as+7J4wA
J0VGMp8F7ig95uIelC77CyAQRDOkhmyPGVqActyxFqOes3nFZ29LdtwQXfw843+E
wFcHundl5qoSmvQ15cY5RR0kCgC/EZyBMAZ7pmh+fvJvAZuPVw2ZqpyYqAi+P5Fh
PXA9ZOYh4X/NazL7H3yfC3avMINj5TEn8pGqlsKa26jkuqBWED708NQaYSM/hfZV
EWOo5SG2MBSTEaUG3w/TsnWImbANePFOmg7l/vdNPft71syijlZLz1nMU9K6tozc
odBzsV5Jmi8AhFBaQm+5J2/4nARIIKGOvfQyOcJcmm+qHxrYQtoF0M0300DKlt5k
YgboGrKCbA/VEAcJAFnLCFYnNBON1fPn6AVkqEY/Y3HIMdiNGHpZyDx290B6IOhv
Qv4bTp5YVLvoA1Y2kqP+Uce+3Q949FX/F4mi4yxXaWs=
`pragma protect end_protected
