// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1B0hLiBSMFtxXVgDbLHtiRVw65PyYdHg5PT+erb5G78HOvEEWqjqSKdNLY0Cud3vztVaDf1vCeEw
G7H1XDoBA2JUVgD5GgBsTWKWGYoWkyYjoJAZWVxmomDErPKt4VELciN3+yADFgqqyP5l0V3hbUpo
PFQIAIuDr/9VZMbC9aUSKm54xEgZ7xDo3Cz72PO+okrZdK3JBSePPVGC6BtjVlSa8msYeKH0stn7
VQEfzqnt3Xqhn2jvpY/mtzyw0sdev5D1hH2ANP4FM3yLL0RKYaPNTx7cr/HYwj3/OQ39nMRMzgYC
Obkf32FV4FtaQEzlLzBqh9GKY4rxJyVloFgLZA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13456)
zVQiEpHbL2b2JgdM3qebpR3/cNE6BKLxA92B+MEHbO3+V+vSQv4xnj1ortIujCYrq96Nz9HBh470
wnk4Nmkb5oTjRnfD08bfcahe0eFO1jfqa2QCS8F22v3HyTCcEm8+A4UJiOz1lS+vbUiH5sx+esbr
bCfRcSK8ojkGMw1+fpwuXZ4QkqtGQTtKSJoMtcblAcJxUWpgtGN4Zx1Sd7QcG0qTSXad/VB9gau6
Ut+1sLj6fz6sgLUdgoPaKXEIppRODX+5fj6EwCJPzTXbu3KfWxk1tt7YwDWuZba0IyLBZ2+ZKFe4
PJ0AuliX7Z8SxMJSagU7NUsocC9MLNyI/2miVfsc3Kv9GQ3SFCYNpDlVfDcMMUTOCNX/ycAxYDOG
XMu/44NgXXzWjlL9s0ebrLG9izh97zVfEV0DNaImXKAvMlu4Jka+WL4xbZ8TQj/FYkLjwhL+X/Lf
fSVbvADQevxJiX9Z7tF4OEmdFA4mafbJACMZoC3icjacNJIxhEm/6wyyWzEkIyVzk34C0t1bYDdz
i3r7BX4fV50C2EO9C2HUGtKuYcSBnEf8Y7ia/NcKmxgAVxCzwwkkBRrLhpz/lKgf/vhESEnNibqJ
kmXuAl7YWGbdb+PyUXPcti4Fc/v58LD/gjHnGAIIU4VYT07MuVK69vJXRBg2v7WnKRoT/d8PHMUV
QFH8kDlTb5A4AB1qpmsvn5Rq0bz1XH9WkGdBHdEC9fcoTTpWS3Us6r3kX/ZMvvwPZUJ1d/1nBTtF
QjqK2vm5+Lzq4p+zoW6WghXYTAg6E/+Di5ZFGqb+YsGj1IulfVoe1yQxZHHgj2IfJuY+FDsI7Jan
CufiMMVawWKDhucOPCIi04LHoCN4oSwEn+ZD2/c74IeLonzg1dajtV/CYECDZObjUmLeP97wfFCD
/kmaXni3gzBwJKlUwEWmifwPmkurbSAMc2VOiO6ROTq2YSdVOgY0TbaYxVmgYm6eF+I05n/4eUhx
evt7/z371AqkH+MKxJngv76GH4n2cgqREe06v4zM/SV4zsQ/IxAGAzOaMy8EtsxzUkU2HmuARlx2
yShK05ebUR7FaigrknEPxifTnKyP4yBnyZYCOEpi28ZjC4C9PSYsHItAntiG4u3kTlqgHYzDamZj
emmWHLZj0rmNAxS5n/6v6vSGmU+62CjK4msodBiTA/6/5OtwF/+UMa2uNQa4uwO3VIgnA0QwGPkO
7NUjWWL+JyoBlGzLPYBao1KaWTgDk6yHE1cUQzCcm7VoFGLJeD6Ldo/Q9/sZp+yrL/rFGl+NAzyu
UXq1qql4YNAkFvhxGvqHKxYzlsU7NPh9WzeI0P9RW5WeMI97+w8F/fOA91iMpMOTuOc7QS3XXi5V
sZpqBQ9YA8ONCtUGBX5cJzo3TRoNL4vaQ4LGkDH38MvhBOVTtIJ28QVRbySZnJwezm4CfOqvA7Ir
EEm7QL8cD4EBVTDVMtVwA4G+BBayqUY9Fvl1WaCFbRi8nPh2t4+dYaCARXqaTQNqGg4KEl32fHE7
Dyev8ici0Gzk+F2F09vvWOmKQAsg0e7EHkGvV8aNy+ocXV1+e/Pe9kLjWOXOSB8iYmkRYW0rkSod
KFzMIXhbSgtGcGJseFiTZarVNXrvcxU3yi6io4fJ96l6jvi+hHkYuBJHnxYslxkmIEX2gEfd8oGm
zMS5AIDn6hlHaHvhANvY88OmcmjsSeganOgF8zK5hDW+YOyfKkWeZDpSoM4OqI2dSgwFjnOQ4/8t
A+IFDqIjL1q/F594ypDvGG33O8KI6AUv5oGJgHJetfRxPmaOj2i5etogumBaMtQPxD6+WOdLFB+5
I2EIg2kzcJqxa1yey2zq8JkVb/t/JI2HoaJ7QB/Ocfvs5Et4YxLsagTN+BNEDY4xaql2w6dog6F8
AjCtbsw7lE1hkDrtJBTlPoXfDdpVt6t7oGawklKbsr3pz7NAMK0Q/jrjjzVuv+7zCptwOnxZ6KJE
OpzM5auUDOuOFXm2T8wrvVWTJSbuYLs9ZcIl0U2MFM8UFMdfpd/12hpLEcz0/sWh1cBdf5DwTi2D
6mrdsNxrgMaEgOUyIEDDDbwKcj6TpJ1EU5V8LMNviWS/ItSXnHKBya+pkst+UbaHtjuV5OqVBccL
hvp8zlGt2pYH4TSOJbsENoToAzPvn3NtAMYxqMk3zNDZJnJUAYt1SR7DfeB1T83Mb5g2uBYcOcjj
g0ku2ujKsDwXR9Jmk9lVLQUo4tCOMKHTkh9He4bGxxV/pt5ZUX+ossAk2Ywpy5SGwYRH6/5NI93z
XZH3NaoqHknC+4tk/1r+vayMw6NOIHKpzF7avlnWAlWCkosi00svJR22DzU3rN49gBS5vJTb+Ux3
Chp003QpI+A3NxpnJsAH4+UbCNG1nY3kegCfe5YbwkqecMRHUG+XnuxYsxP30CZjXSxEyZtK5V87
QuPdWIHyxUI9tufWSlBm5Xw6Zpg7gEk9s913UyKhAFIxZ5TmUFjHFfg19OGghCn7AmzsjsjZUmGa
JI4R3Hk8ofbcxHC769nWWP2YGFbcgM/dYnKkiNYfQzBRxB4jFtPieUhuf8Zt5JlPPMLz/atdduFh
MP8bpjXsRWLfI8Evgk8p/eVqe960iSgSo459k+Z7qDEKpTk0HZv/LMHGLtVoKwflXnQj5NTFtl4X
LK+jMbVRITsHepOIWq1aci4ydnBDBDQSADr+hUcIH3lv9LYksYjjNb3FePhQLs/XLoTdqtah/hTu
ZYq3MuWuBG2IePQah7SRwMaojlHHepnNOA9kDoOQ4vGS98I6FpA7hTLHAauV0dUjJhmD8wfRd+Wj
GrTeR88GDtoK41SbP6V/9iCEpxWZaDNeohsA9qbgftda3ZBQ26bskxI4+mls4BGYMU311rwPye2r
kjbQSvnScmmUcGsBLhcTIbO4RTl9DW8d5ZrwV3rNgAdAGwG+K90BPix9vwMD+pc5alWdqZs1miEY
SuOqz36X3uqOe1TZDtf+6tzG5lgFN1eKpSEIdQc5VaHGpxmZiYOQ079JzwphD/FfP2vsKfefwuHD
27KImSQxOgR8ng+VKRDQMNe32yZx6MPOijTbTUDBEogLkEk6OCweIz2yYgFQEGheLzRDnOggHUIV
HFPvfBHJwXBN2P2ndG+Z1/AbP93NrdCUwopiHHbJsAYx3/2HSMUJ7Ye/4VD53ew5v9nHaBAF565v
lNdpN9i2v7jSMbiCd5M/epmrOrHq55JnVjITq5HSj6iTJ0usb2LAusN3tvEomq6teF4qf5Anod4g
v8Z6+FxSrJKpOGAu95oaoPs4tPiFi63CjXL28cx2oi928YNNf1pmoDw9wP2MHPf3ksT6/5Letnsm
M7K+6NTpcx+GLbllyZcnyo4lAHvjNo1gKQz8msUn7rL27p2H8Xl2hhrgFsdBhwsYiu6WnK6jxLJ+
5v+0yuQS+5pblN6ohhD3b9bbapTaGn5ZLdeZXEJxHTiUxi4hvtTvWZle4EZQ3gufnR3ElR3PYnhI
+54h17IiWk7BsyQ/hIJ7IoMxzMRKUawA2VWfK/cdh0YUmBTMq/UJu2kbDYgi2xtTTtr9/MwgPc66
qWeuZq4vsEWuOyp+lABXHSxX3/UJxV1SHzypiWZOmhFjPXMhlmUWcX7Xmdbj8DHOujSp6/Wyb+VN
BUnBLYOS3F4lpNHaV6a8l3tmeWhhF9FuAf7KsQNQrNfyq2DCSnAp6N/GO2Keuk4dqi5yqqycrFzX
12LY+VBk5CxfVMn3SbPWOEAHKq9bRjE1R+d/Ft1T+ebDdgjylTrozuWvreIYvUQwpaqhAdgGAaqu
xeOKhf1IfcuE/rWfxNVf/POBCjPs1JTZwV5a+//zmBDW7O4U7c1xRmOddBhsRZvkTu3ITKtzuXws
24sJC3pLko/xifHExLUwjlp8uLlEUadjKzXsJTwarZrvNGUiRA2268iKiNbu3zthYp49yGmriD9v
nDEGiGOl49pmbh+3G6VyxbjXy1IJ/OgsCJIlmnR2CH3IV+VtLVhUSn4KAwzkIQfNpXfy7peWNdhU
0nZpsJSYgcP7mJC1pIxjxGiISTJe/TTuK+B2Fgzbpqv12BmGLioLf45pubH5e8GfVlsrUf7l9Aa7
YO61VN/0ErjhmGhF/nB4WPZFS5pL8nb+T4sn08sXcu2rcPFYor95SIFSwuPmotciwuJhyhnvPO20
lg66huy/rBWiv3C7LDs1NKfeGgHu+J5TaazHVFKBuoxm/wjCt6gSe/1SBG5KSauDQ+jjeFi2sQ+C
a1qwvndVSMmky1eV2TpZgvA6V8UgyAHc/7+GzJIe+0HiZmsdXScZFYFAFFxCY5hYfGRGdqP5i1zq
khu+CsX+em4lEUhrwLRlzy1T3fGmUFkXnaN3n5HFRVU3bF1KgKGvX83+S6gHSR8BHU7D5mbzEgMP
0oCJbuFA4K6Uqz/UX1h5OeY/2RuFhUcEzlhbZZXZzDE9HNLIeVdUKVpaDWFLcs+glfebERppLAO2
PHHUbKPnNWSztIdxM4JTeU100NPRoIb/7fIFZLAjcvKY8Vs2j/MkkzfEyRWh+DGIVjjYq9OzK+Ff
h36D58tS444GnOyprYKzn33wKeAsFmIO9HydjQZzYN6bqGsMwDYmKKiJtMglNxTW23oNpTZxfVD0
7W60VRhxVs1rmDAbKmC/WH+Z74cHAF0VVQlKhCknu7ieu9/PTl3/0D7RS1YuclupqxDj+8Q6hUy/
Vi0w8/ReoTZ1JejpRPdL7SdwEWm+rxu/qusZtFuHAff/jEijkBfXjMvhdApkChAC1UyfoAZM98x0
1ie5DCEE4AAOQlD55wQ8IB2/je8Swf73AKKM9g1ZGyvPqfDOB6Bz2w0np9+K7k3VKx8O7gPTr63O
rZo/frPIxvG7s1+fUX8Vf73jbZfDlz4hDGFP1GYEZOpHezlJjf2IvgzGWzqgQwPoyepHsSXP8U6U
hrkwrdYIR0yHcNtIgeAKJf78ROQv/V+c62T7DS3N/++JK7T4EEnTqUi6iutsYmq9gMYRzHaj2n1f
mNEZikX7e5Fh8Agi4kngzTbtPOGdUc9lZ4zpe/CfI/ZXG7k3K2JKLxlgn+y0XgH9U6317Nc85yA1
HW/KU2+dDTOpUJPua8pBRIWJucVQILrUyoDzBp4qEGFKeJQXXmfTAFC2IqB/E1F4wMEqcx08PFfZ
rJJ1KW59ExMwFPqc7tBQsWtIeJDodEje53bZEGADz3WKjnM9c3aHIDFJNHbzIEO1PVWQjgXBkNAN
dAMKQgjRbvFtQBdfgJzIaJ/SqqzvQYqa72tjlHA3li9sV8woOOCzuERpuOQ0TmaYoSRDoL3458OA
7zUtV+EBXu9FDu6QpoSFZY2FDu2e6N7LxNnMHXtQEyMWhI89WymP2CPg1BP9/KxrEk+xIjCoEU/f
58pusptqEJDgQc3M88Hxycg8bgltO1gG3amJEalR8EXYuB5rAM9VgMX3q2n5wmJmQoYtdMWwqkVg
Euh41855DPIZVxXxoCj2zp9UoM3xuBZOCZT02qeZQFmIaTJDYa1DljjlswDvo1J7eDC0bBsmduGz
qhWxcA3Wyaq6nSQnjFy50kY6CAAmzWaCsg9EyuosWB8b5nuUht2vs7ghCh9BhwYrkc8EKGbjygTT
2s79GFgtYu1VKDZmIA6r0I+1RHyIbVU+8UkwMG8SKICmceoizCbmpxDCjcY1mEM2fS3WyqxBpxAx
vHYjyXaqSyiK3q2UL9hcdUNC1+bkGvtjTSAXMlSO4gDzWqv/y/z5yCNn0ur1tJ2zxkr69DiVAJ1v
NwL61XwLhivYkr8sn++K2OsOCwR7VRE9GLrSRUvZnTDL+ShXizSo8UaUe5nmyWTEDPyMDja/vTYx
r+rVCzMgrHHkGgO9D65+fxK0/qnGp5MeQwAfW1XNsrZgKJRJXrTQIZdY+GCmGjOKEmhKMzUI+htP
GDoSk4P+K/01PVvTHh1MsSASKY/IgIfChBRmM0wk39hclo8geZ2jYkyye7hsOnFPBazFmOGC1nuI
JHwR3wwU+y9kxM57LcR2ZPhqNeyg3t6KomxiRhfQ9OOFf4Aokt8qRj/YkMN5jwreIlRtAcY6SUFp
8rFy33rLPUrkWXWCKRPRf/68Hs8DZxVpxrdYQUGp826t6RPI1tIPVUYfKP3Uniyjnc5wrbuX+ioP
Le409pRtOluhGPMIK81CHJIhSapGqDEt/HWYOaMzuKtdGOHsULQ8Fa+u81VIYAlDIEAMnsVITUke
ltZBPK9+vyy9rdFu01EPHPFDz9efVOoUP71fAFhFyC422f72JcyndWrgsQS5YzAkL3Z3ZawCvW0j
mi6rtio7f2tkGN2BMghmHLe/u/lr9RtG4jchbzYj9ZHP6KD5cKQRDsrXRXm6TV2Ea1Pk4U0SPbs+
jW6wzEOEx0RoWb7NHlLo1T3p1U28uiWDD85691STYYwSUH/4QCzPviCy2XBGLH6VUoKaYWP7AmgC
vtAKG+BRs8e7SuVqLjr9dXz58EsJnuHLQ9VxIGMRpUKGmwDosgOjNiSAFxiYwljnO2e/nql71Xr0
aBZ5JS4OFdLBq+NzC7kGM09dOIaYZcW5g12f7Exa9pyg+FA6ZkBQRLVA/J1GIanb4ZXY//lzOU/v
El9KYGy8jaqBlpJM7Mg8R9EzoWYRsFrYge416MxxbTtPiGKezNisr/ix2tJJx2RsEwmSCbgZM/Ay
r9IJ8GDMUj5wzjLe4kXX4bJOfl5U4tBzxQiDeO6Vq/YMPghRQgkNuYUqasjrkd9b0GueyBRTFbAU
4RR75CTTfxxrAxevq4fY8IVhkLvZdxPP86/we4sWN49M+KN/YdhU1TNywyIhhrUv/g9ZMWtO+H1A
+WyfxS33f944wbyEw3WACavJP+W+b50Pt8dPZsTq9w1lJ9f3UHPMAMctM6ms1OLNwPoE7U4VQ/nw
WWRYzNkNS9RKhU+SIM/nYH7KqAh3tjdU20m8Y9LG06yd8zpEwDYxYjtYPNKCV0eTFXi1V0vQ3WHc
B+eaAC/Mb5FbdEPo2+b82fnaubOkBZtGAdkkgfhbvYcX8xDtsOy6UuD8VP2MKvqCle16l6heFscZ
C3ayexnf935//qFHS5BDyPRjwPpaR6p0RDpJl2Wq5UmarZmUnfLpVYsQkHetPeGmP8B4ji8D6NhT
qNuuODfPD3IuDm+xkqqbIOd4TD1+CRZZXeLF/Lka+VT4Xd1/Fbh3wHPmK3UfcLks+DA/rU6aIUWj
5KfyFPXMENZCRs1V6Etj/0duyMtdvX6KhKHGUQCqq6MRA/S7NaWSGSPYWCvvcCg5hdZhS2j4SzKP
qhFwQxhGc7bwfdXPKBzaUmQdVROJMKneYalZoW1hLtSPDS/P5k2VcYJR9oGFrzau9b8IObVvEdhR
YyE2mjL65s+czHIGyDFiPYCnaklju+blH+7OHeUq64SqTjwo3aTbcpNkqYj2/RfYenUrprkTziOd
vWDN3r1E1OEN+aO3TyAe6bObR2/jFK2N7+Y5x4dkPeVWlcYMHoPxyxW7a7r0STNW18ID1zQfqIde
sEoqRq38NLB6LkhLdyzR+4qBMNZfOc4yfoJRfk3FWZiZzBSnotVUDyzVmCGOFf7ba1+Wmkvtboyl
0sSHPSaZOnhbzfLvLGYrXpcBwKPF2mr3TgoGZ9IE+X2+A69kviIKwxkKknPfrCNw5xQLThgRVl6v
bd5hL5L+ePR9hglOP1fyA5XWLZI+cbFFtukdbovHAS8acVd4bTNoAkhsr1+niulqBOnaCW9l90Pn
Fq0oeaA955kPeSsl5k29iUkbJpgHIb3FIXySO81dNJJROVa11EvoKXbnweFk0FsxPRwJBHcUuukd
NAAV+XwBXGq7nsBpjHZhTkgJTs3WgNVerVdVZrUopJXkMJIOnEq1SEXiVugL2FZlJWnl5f+3/S2n
8sR6FjTKS4puuDS48eVBlsryTNNDPHK5xN+2rhLGFnWRCM1iarB5xY2qCf3vcrlaFZUG3j5TrRAE
5FK1HrwGBA6HIbQ0l85AXFJdtpR9WeTYy52KmzYcgG3fCgHHWzik9ToHBvI/Xz3uNfWbLfhfTVW3
USAgSOy61AXwfoI/8NLcRh1+YabSj7WqPVxjiv2Lzr7LggAGiD6scTwYpAN0/tBSjR/LTEEnbFNA
qqKoiziSny1weiJIDM4iGhs6GdaiRezsML5dN5WOtysDG/481ldOWJ2r6bTQJGYnZQD3GVITTF/O
AcmGDoiVxYQ6Bgov2fbQ1zf2Tw28kQ8k2uQyLdqaavv4EImkd6bSVNJTu+im6Bi2ggiEkUW2QDIe
ZV5Cy5OJ2LWjMeeGau3Vv4Qte+2rViSN33SlARREYTGxx1smk0jf0sFID+c8GMmwNpOLmxZcp3Nj
O0Z/NWjM3rfh9QBDTlaR3cGzxMNGhFS2hBSp571vrt3ExbhPYwRrY4O7aRrodVsLU+ExKP1sojEJ
Ep4NhGPlEQXtaQjGCtI9S1kssU/QFLhS3WSiS857kvlueiKl9nDfVfLmuVv3p0PL1BCp0vSwNJhK
18C/gi32+v4ZnQLVmBzwTxKpALy/NrWmYcWL9JHdPTr7xaoqN/REmMPdRXw6qJQ9C977WAi0Z9AA
h8Wn73vIwVIvRT+epO3+MsqkuDf8pOhsNdTVjeHVOoRyElXZvyNzFvxYZLOlSweiOgS0tYKjRlZ+
UIthQDGeeZOpvT7SeWlcvAdPMqN1bq+xKHHpxQ/vePl8fmI0qK1BuKjBsBNAmLdXGoji+Xifh2nh
TyjicICG6ZilOEQY0y3Ma7DbF6IwDuMNDTbAl3fPsLWHzP+vugjj1CbtSD/QM1HrrJ0wCJ1Em3B/
qDqY9w/OyuNWT6gn9Ne2Uc9G3qCaDT5uTkrEW88G/KJIVykSaAsVfFPmLP9df4uSmf/vaKxGA3vE
hgAcvUIbi1WZQPCfutI4N4NYjQu2s1Nt3cLs66KG8s3q/9neHRkAfAZkQhqo0otbYm4TpvCPS4Je
YALQy/jILa2IxmKz9WH9qej8A1VrCuiVhu4jogfZZiQoi8ahEwqu1IznfNHXnkQYv9g/VVHyigNh
7+vPLOLvdSHfWlQWUFkM8xxFcXALnQ8j+zaV2r3UcC0YcgY+T4rlKoAXY4yICz9cm1JTfum05xwI
3BD3FCR+AGEZmHvcwNeXmjT/4pRnwBc3/tZS165CamCz7AoHvmdt22rEA8Hzg6ha6wcxbvK0lUjC
VUPq8Zn1PyTerBs6d/Q4fiB8ExQHSgjxCYCJzrfwqktvM5PmjndCdaYKucbWG7R0upMgiw8D2mDd
P8ojlkNcTtrjCBnPrIEb4zznlqvazjJrzwbZlpSaAbRwryv54pXhwnN/T3peIu6yvDakvjgKvRPq
AaWKnqc40px5XU9cyuvZ5ZrEmF1lsNCujeswUjYNOIhPsYoTb8sfvm7ZFN5DLPlgbcimLIw3FHu1
Z63MHAL9EAqS2+gitm2mU+YVZfBiHo2Gui24fGsHuQA3ro3oM2utC3sooMyXJvhFJCPeiApekbKX
G5n/DBWkAyYDsgv0cHszwZzgZ4Dx1zaf5Ak/5cRxrkH0K8oQ5efK2ZvvCEz4fy7ZTE82GexQKG23
CX5EVvexP7hbvhwWNbtcA0xLTjZxLUsYaNCmtglMPLjfEvE/9ci9v+mpQvQoI0e7KoIp80QNyp4Y
XstBVqCOYvt5SP14CcMcjiGItLmYPYvzgcQFpAid18FZ1jUyBY2xeYUBOyrOcl3yhwFeXXRl0Eb5
r6mWTwCax2LMCuE52Lz5o5bD1+tfdtmc4SHFZkVn3uBcII8S7okAAOTOzgNF3Cc7NsoJj9BKrQDo
wyeH27qRoxRTdIleVf7mpSkeaQOzBoUynC4m4TImc92faClPKF1IygOjMgj+ZuIX4Ph/IhA9vQrk
fnngeoJnyHYjjJZ59rLVwxkfdXcsVLY4nQj5RuyzdMBMXyVRanchwUvibyBl1VVc1NqtGqiEOGpU
hFOVpICYv4MtQPWDzX3xl7sVL+GSIRIgY6n6yEXZjW/iGHT4FCpXDNDdGO1YjSf4fBbmSb0u9+o5
yeEjffeu1xENubESc+VRUJKmFHjmpPxyBoBGounK6OXzzpGSvkMZK2jLkUQzy85tDsaK8sscm7H0
I+aGT0mO72vt4+94v4wTLhbkWLOt9rO6zSss2GTD1ZisUfZcVvhT7iIAbzr2rd5qj1oKpNx2rLTH
Kv/jP/Kz/jc0Lzw3emWguGy09lW3qfzWFcEbC4CfLsymSYjOvMlwWdhK+0g3yL/H3piEj8hEJH4D
0VAKF2f+xGtL2noT1l+jiXuLgjTMLl3QWnsboEpweWImzPwMLkeC6ao+uRosoFDHDZ70uqe6mykG
qaErDTtTnb/dDmMrBPfMtbLjov5EsmWb0u1V0yVWfkK9eQ6joV2VQyzeaVbdq4LcIfk3U9c6oAnh
b54iZhPXUztorgTSA/NN2rPGqD7xiaIjidaWqs4cmmFlC9nWJIp9qyM1kTqWD3FaOChCuOiiUunB
MA6Wu26CYIz9ztjRjvKiy3ao8c0Otua1OQepXcpOya0CqrYcBu6X0oovwtV+fDarsSVcuvYztYVi
e31mZ9Cgnp8nyW97meZrbcqxI90oQ/RqitL3v0vtfDcSP2UkCOaAzUYbzVeL1g7aRJ4J+VhmpbfJ
60muKMyynbIyKotbr7yCSUknFT5z0iG+GcRHE59jbl0mSaAKUCRBJBVz07E3S2bb0FSM8vDiupBL
NaMceD8peM4H5X51PYa0wkFie7CMuCjsDIEKX2qESweeZVrVcT0jI8KVBsDhwWGn5DFoHMo/8MNM
loTjY/BIkDQkamYPP5FWMdiy7kHcFnvPuFGFimOuTC4LVFfX0q8gOpeBkkI7T4N5o0WtfRfzga2p
1YJCEH4FMOJ3G6OARcPcBDgBr/PjMO28TT3r6d3HMtX66vY6VXiOPgsebvUz2f2rVo4yQIeEBig1
zvvXl+nrXNRklMmLk0ufxd48M7a9QEqWDgZR7KH1jmj4zam/dCJOBpHjnp/RKxe99heOmPDfR3Ay
7RFELXH55JCTbn4lri9PvGSpJpZ3j9pbMt+xCstnsVl6cde1tWpm5YCuHgve74n+7HcFAq0/YHBG
/En/N5yeSYUpalucwUMHgP2vZvqqWQ3f/cbw3A8lHStChYt9K4TsGy1CtiqP6z1B0qeAZQQm6y6G
TB2klr9lTxSgcHpndUd5zOQCky5oJgzchxxk4roe0aEn9bMI2sFm5SYNyvBCls0kpljk8vtTWWUM
mX5FR9cYVs8HJPsVV4slFvmfjJj4pTx1jj5G5yGY0piGJIKNKS7Nffq4/JN7+uIcNlY3iW6BQh0W
0EwhW4tS/Vp3uf5c7hwrMAh4YZ1Q7OdwfRHgqDFDToMijqi7SLa7HrXo491cb1eODD5hZWYziRoL
eLL3rWkxYjRYUhjGzI8wweqtQsXDtURrflyQGY/rNOkV/zafeoL9PWq8iNpg6t8EJbauBIOfhDYZ
Z/j0JIaf6rR6L6btls93uCvgENnLCDO5x55iCDII4/qvpKiOtJLZDRJaF4SHCAG+hC3lmsmRPgl9
BwB2tGdWXyAX7WwwFUZm4sLuIQjK3WWoU6N81751ACcMf0k6uqf7uG3uI2wQ5RjS3sYDqyPd48oV
EEZd2zxoz07t87RtoUB/7pTSb9w8kd2TNJA+sounki76maqKHo2mf1q3wl90upOzvIcAtM+4QTBR
xLnLicQVnrjsQETWiRKXL0TwO/blh1t6o9tMLBXjuH5cMWqlreaD7+yZkEWVOGac+gDSjRvGF4/U
ZUY+Fw3mOCDqd6Tofd3oVNrMJ8OyPRD9cyjC6IZM9+hQkdjy++CE07qiClUvWtmtR0veURVE90xV
HX0eS69Ip/5SZ/S8obYaJ8QoJPx6urx5sWovEhZLAO+bym55PBbBCDOsyYJOEZhR8C6inUXjYizl
n040+fRE8EWJ/hCgq3qp9TwC6LR+N+FQ6NhcJXL0Oaf5FmOmGVAPfw6rLBb56i/NaOOrQvc7KGBY
aUvF54bQ1gIVzeOfnv6U6+cX968H/ZO36iWJ5DdZ2yKNa4fssErhRqItN2WF/fHYjQfQra/jlD/q
u1PaU6oQE8W7y6QeblRTjL0TKnBav32iOeKQ6Yz35in3zIYtCVAl7OtBdj41hElbeOZwOm2V1jAJ
Gqg/Prz//o8NvJX4okQcVf4d0uQkV9xvbrylX+kTDF3yTcoUtMnOYgpRd/Jql3UhDdVNy5m4XE4D
mmkuq7nCU4VS87Mb2lFyfucxUMotUu0E0SFAhfPBoRx+dSfMaE8ojy9p6wW/oc/rZyn/ikeuEXOk
HgR/JigObOSwBSMvhCf10jDSOS5Qiby2vudIcCvSqt1rb1D+ujzWYQefNpyEamhYdCnEV3eYrKNU
5q9h7DNDMTqdmvIVW21Gf3vRQB2IHvytX87JomcjeRKpDKwUPEV/+issx2PNKUFioWtur6OLptGa
EAKSwyyzQoHE8MNsKPXY6SiAXy/F+M/Wh6tfmerB5j4ZL4qBPNNBlcSWwY/m1ysSBQWHNF7rhgV9
7aThB/zB7SDnw0lsbUBsQkP6oU/PPIFKwPZdKJsue1bDfKYXlHyW3lAQy/WfkoMoBYa39P/tPqTu
f3y9q0ISgPU94YrFUfv7vy8nhoa+jJhV+8dEca+48WoKx4DiY9Tgxs1wj5WXj9QI6v9zHImgpaxG
/n4zp3fO6MHjejg9ZGPbZ1EqmyAhFFV5B3QHopKVTmELVWheBRgX2n4Y4+bcAQEWXb331qFsws8O
Jcy5qX+vWX15AK1dDOgTYrQv7PaENtarjJK4S9APb+qJ26utxxhq7AnooWXug2dgqL8x5xcLoxoi
qFWj0XNSsC3crEgpBZb2yem+LP98BuPNwhajGzQDqMMlMo7WqSXWAEpKVqCq/6MpdIjCBQK3pcjR
rF/W2vPcGsgHMaYvfcpWclGio/Bn7DYn/0QLu4rTKssbni8zIwpQOvVpe6bATxsYjhGAKlPsrGjz
qxBAEVj6/J3rab+L3TfeF3F46eCafN9I6+L7I8+UYkTMV9xHzTxWQYvcqJMrtkP8xfAXZoqGpYir
4NPL2+l98vC1uuuTFMJgPWOhL2Bd9duf0EdD7pAnQcr4cuGRcQxyPtgyUgSUfnxWnTFukX1gbIv4
hf5PU5LiPBlMWH2YSEoHBLkIvGUh/p2VILMRxai8K44EOICeZZVKLeKczmZP0Em27eZqis0n/N+f
ezTihE1OrAAPrhJ1hKhZr15ZVjf75gh5ERHpyZJmS04DUNDVIVqNrRgeLg/pGr/ZaBlVXTkrS+nP
35PELOaZDr7saZjucMK/LXj/HtQjlfsOENVbAHKdBj4vFb6gvuUFbffj/KIEMjcWyqsOO4J2Njsc
Gt55ZE2KQKeuUUG3Z6J3qn+EMnwBsmHk6faOtaaN1cMd1GxTwkymHvr3R5clZeNLOLu0tFBLeetU
0PMRTha7GH71qlRQdiXgxoJjJTdDSHM/hOFYvBkHsPHf8RgDq9u+9Ywt2aUpudiNMpsYYlQ40bQY
UAJrBaMJu9LS+KBqC4bp/dC1vkXoh76t/s3O4WQPzEy9Dl32nHeTuMwMHQm+q9FJbn8xIHlpnDcK
jpTQyQo9ZQ4/v9gQzH9V1KlD8BE8+Cw5Z5RFuQJ8LlgG5i+eyLuTftIV5osAC0HvP5TlC2tBPrKl
6Gvrjp9dg7i6oI0zdDbFpvtyoOSwnlLBIY671miKakbGiecDtqdQIris05EGFccCy2nFRLNTRH95
uJLBR4JcDujx3J0FWqcjIjhVMi04HEeClKEKFYhO4mpE5btyQN0s/qHstOe4khYR4ekvfeRq3W+x
bBaayJI4tgVUlVAEcxpHp2VNXOCs6UNZNo1UFz7nH68+G9oJPPqYEgeLoIOLAOedjjXjuaKL3Bny
W3S/1F42G1OCvZX2J6uusQqyIYyNTDzKUoazPe46LHyhk2O7bkHiEDn6EQGp6y8F3ei8dYa20VvF
S2lwm8ppZmHFu9DqsB0iG2HLkCOUP5G4U1voBdLvxfXSDOSVPLVyRKgyI/RK1HeidyIFVDtzeCIv
FdarIMGQ+/SSA15IhF36qKXehcj1168f/bXlWLDGCrSMZhaZ3ISwqzQG0tHo6jCXuGhmxcXbnRLH
cG7V3SOSp8WMvlyuge/rNWovTiIUvD5HzRAEAooc4Zj/raKMzdYQjxPYPp90gwlUgSRDhnPQbIa2
8xhDe1CycbsSIIuspRPXLTRJhgSYBe7Pr/SaTyDYJh40u97ChgntYH+5xaULyVLC+aTByMpjugyT
WBaME7HHrdz/Icz0KucXbhb/ldIENczil8ULG+T4kjf2GbaQJgTFGXrwsiaAOjb2VU70kmNrUm3O
2AGg71OjjbDBdXtPV2/IXmmPE8VuNU2CDpOEfPiTkNe0zdqnJLs3+t+mu90U3Hv8ObqFQ4HNZ+4Z
43L41/oQLlMstishe95gM5orntR/JksOwWo0s23sKC3RRhQuTOZddfITdIrFT/m4JFPJ1U9cHFkc
unAvH74j5m8dzyzd3wdej3sth4ZXTMxEhH6/5EJwE4+hKdxSWQWrg4K8NGlQESqt9fEem3dndbPC
3P5TbFaIWDKUeQjCzsbwDhtfVVNPw8k/NiYspjs2If9WkbR5XLC4GoxZPpCrdXeuRkXSVoKqWggh
HwvA5Xxlp1P/hI2hZGOd0dwSYQrb6eJyMdYSaGHIh8lZC9cI+6B7yUHFlp8LyGCLW8g1StsBXlpp
XQ342og2hPhFPV3cgUoVO4Uz3U+KAwnEfzV7y/lAxO4/cf49R/t5qc01VVB4Z+Gxo7UtY8oac7+N
oN2gLuL0HcjDmAKJAUoFcTmNTjQ3NZFSWV0GmQeYmVPPNQMra+LASvDq4Nokx0/eWpsWhY3bZXkJ
JHm2k+kgzp5+wkeEQoG9JkqRAYjaQm5BPvMBajQh7CpX9ni+aoedNPzmTCbBErZwp5CbXyRUdb4c
OC4f6+vZRl1yx6GnGmL6/CQFDcRipaBNZ4GOU6ZTT6Tw09ZhaEw/v8yVUin1Pny2YZSLNq1myjPy
vPJ04Tr13SBiFCKsgrQTT++24TqrRol8CweOvM89pFkABaQBcg/VHJC/2k2WhLrUhzYHkAaFMFIt
weGuQeTsJXf4+YVrkHNQVOgCmd/UE6Lqx4AGauOUtIItZTLZELP2ZJmedT+ZIHZVNLEjQqYTbb1H
pIaRIQ2eZfmZiAoivjmum+024AkF2QFd2UWeCe5b4w4gqGVxr4yjLoch8EPYmyGlFJu8Zx/XgXWH
/7MMbnp4W+N3pzesjuUhqwn8MsWvPntmgIApHd08Icx7nP/S+dIaHzCV6WHa0bDvgD0Rt8nCqCgi
kWfrl6fPK2pn9t7/iIHQJmkhffNly4Lv+hKxee+mYlX+n34/TopEkW5MGP6ocZmdimmnKAtkL5b3
qcl/O2GqnkWPQucUVqxj/gTEAw0XHGyyFbiVtJ0ikPcoqlxcMyoPBsm42u5XYF49NIvpX7iZEhv5
/+kc0H1197P1QrK7e6C81GO1JXVmRFr2ZSUjY0Ve3wrA4ALmjM50GG8aL0pGzQ4qMSWcXHoXyC6K
r5iwueQ+BbioRYKSHpPtviyKgL5aXZOv0Sj0bTDvhap8ZYMdIwVuzmT8b/kot21qQiUrjvpq7WMt
viG0u/AwJGiI0phhgJ+bszz9t+YtGRNcZJPRmcy8aUEcXYdBj10aZ19HpNyUYQVp5cOlkxqRuThf
x/KLyhrS2bBZZBQbCKfAaotuS9NPNVdaWjtlI7L6jxpYcCNoMMOdyFIcIlsWN0qO23TlIGba2UBD
lFGgcv+Ba2W1WTYd4BUQ3zEigxlqlvIYqVjuMQJ1on3sRrIS4pwenxRvmVYWgNx+x+lIBlQpjR17
jJwOW+essyOc9kOnoc2crdHqJrbL2QiR2r3m5DsO9dNHUGCtJtbj3Str1YyG42y1JxMBaf2FQ0m0
ki+G/0pK5WaY5MfP4bACqzq18x4eEX6lMLz1HsFB9QSPLbopjZFJY0y8vxprgwSqxSNHiUFXCP3b
SH/DlA7yfK4YSDgrlexe2pfeTE3vgJrXdSweZT7ncNY5Ue75Bt5zi0EGGuAGW37P9BK2q/RorF/U
DiwQ5ohVMlzCcP+yfLFHyXzLSSoQxEdJVx2e9B7lpwzliU3PnSx8TzrfsWdQJEsa6oKzsuKMe9nF
iI0y/RpzjDpagN/sYSJ58qOgC0XPsol8xh6Kv2fYW2xR99rKUo6Hy4D9T1G9PHVfN4RNV6sFuDN4
GJJTP4/6U/DeXLfgIxCb1WtB9GzuTk1VQd6sry/xhUtNi/kImyP6MhKqHb9f0Hl/lukC3u/VYu/2
xY4BZ7QmZscIjwn0t13NKI2NXzPdPiOznAVEb0FqXD9d3Nx5F+1apJGIuJT1iN9zvs6KVhE1ctVV
Kq3wNgugG9q1HC+5LMX/XWAYedGhTaxe+HQobMuqY5cfD2CPkWrcLoJf5XBskr8yhLQ80JT+XCqj
488YV5tUVGeABC+Fc3dKPIfnna8xk4cQI4Wod2IgZ1QAsZr3Ehht5wHWDp0JeydvUr9unGXErwMT
UMt8+AIXSfnjGb5X7ESKtAkc3HvjXVCjoir2yyia8XeVDX4X9Q3VQfUCnKH7dOgTFCzXFXmXzAvk
By+6DG/DebQAxqF4pA5qWbUMyRRwJ1n0mhhRME2f38SU/imaQN0XP5mX1zIsD/spLfEm3Kn6RinM
1tOGIWfSchHH8WxK/o6EX4YB/EKf9IlmSTcgnKty8JZaWiwxwxod+xXJcbTvNbDpBiHRWJYUpOCo
TKhFNAmO0tJNUym0IRWCcWdvXu4V8azmfBOQgp0Dn70gVHz+6T9249Zt3MBe/wVhIREIRPheBRNf
wIzZTsOhag8r4iXOkHA2EPSu22lBZ7HrYi4IlmoiFSCOEgrqxcQq5ydMEaDOW3KcNCI/lqR44R1t
g1+j5RcWoA0QciOOH7bkbI02cLjx6J0XVfK4dwrdMpqa2bE1PXQe5T8BKGlMOk4RM7jVGkSzbyAS
HNcREMUXf0LBA6Why7lhXc+Cmrwy6a3nzUznzEE9YjNlszmLApACV/sSlZkqjoS6PC/ypXiUvhom
YNjoEYO0SQeEt/N7dCOg+lz2a7SRNJhmbik8yUKg5CZVbsqMChaLepM2vOokaM7DQIJ4/LC4zO8P
aCMgceyixLNJEpDds6ONI1nTvdOkt1OILgDIJxc/ACn6HRyDr7DvBpXja2aGcJYc6qiuNr8UG0A7
Pq3OzZP+0WBs7HEICr4VCdoBMolnlSHNTJMzRPblJCwig1mO4kXccZzv58YseSBXVHFEUCIhjCi5
qQD7Os5CAARhDr+qAacSBUxZeeGDH7N4WfJ+qt/MpT9ueJxyT95gCsuUvGjz8Z2/6jtoE8h6EA2r
UWdj6OyZsQ3+tRzEgEKGfH5DZce4Y74BxlrgDALTM4tIBXSkFuUZ82vLzEx4MOlv9dsYBuEpZIIV
4GrJh75IGy/Yh+Rm0w/Gzlnl02VzZCtJbi5XJxu+9WUvjC6+Pnc3xa0NaKQNdp4J3ps5wORIBGww
MyZnoay7HJ/lopI8weaA0ROXztaS9zLgpVEtZWNgZXiDSMPUUEcYKfTKu2aTBnhIcIyf853s4Z5t
Dv481DYZqUlxhxqcg4NbWidHrla0IB+mZrHKKCNo7zQ0I8Z0h2axe7qHwkJOP/cJUyCiz94vZwqI
i/P/BceX6IELt81fb1gMysgCaJG/2bLrL4FWmHt5DrH0OZNllt4I2KAM0UIN5/aKd8IVtyZBKk9Y
NW8X3r4z9hc85MDLVcoFmnU5O2Qn64si67AzWGtBb1QKbSWPaOxCb9u4ZS9himyQHDcMwxsB+SK6
foao48pTt8kp/e7BNjfsjmic2Cy8YtGz68oV2Dd0zTW9l+OjokMEu2O4ztq14olBY2RRAtf1NcaK
3otjHg==
`pragma protect end_protected
