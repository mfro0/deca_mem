// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IFaXK4ZaVbGK1ABoAHNhjEh8h3EiMneVrb0WczAXtRBw0lmzNIlAjOzqdazq20zb
BzXaaZRLHNN/QO8HLcLTq+n2cdFy5Xp9f/SLGP9RCKkdolrD2nVp79o52kz8lIQH
ZYscG/kehM0EbJO/T7RnRLRTYT0wDJsEaCwZEX1OS14=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18864)
mnIxLEG8evpYtUT40m5E7p2TkTeVG7XhuTwP8PPrHnXeFA6UZCrwQl1yBM8I7hld
8od6aMHNOLeGjiRoc6ER5sJH1Y59bLkqQGRZZrQZusluTNNR1XaSqefxow396Qvi
Ga9O+w/d1i1JgXSDEUPjxz6sffdidu977tWqpnq+TOW71s7OXFOP8od5er9WaSJy
VGA0dWNkkrIZJcyb6p7Rqwn9OpbmXQjbS7O1OqY2OaYSkE9W+Zoc2VGKCuV7mSze
Cvt9nn0S8fFY1mUj3tGo4c94nZfrqdwzpV9fdbCXipIL9rTB0mwmYSjZldWhoV2I
iWld1GKdpxIfThb6dNso5lEGX16jYO6LdFUzW4AZ6hTbjyM3uA2GMQe2/R3VV4bt
KaAHX1m3uC2Y6xQWXuUrKU5+Pq8aiPEHsC8XMlXMxDpDClvjrgotob2TZhRhkzVy
xB6bovnMGd1tawtvtH+AJvkDwC6q4BYb16CMdjE3kiNS5dLjzgHysKOvLlzdBRkD
AfZJ1uZMwADfg8ql/fzfADrPJh5kSQYDN1mDQ9UMdz3p2rW8wnhYQQNnAb8ZEV7f
dCgsRbjPzL0BrxbCjgh+D6J1f3+EYg2avTAVB45w4aLSboZW6Dr+7p+neQRIEdbU
dc5hs3nSKK9z0eJCHL+lLh2zSDVlWMKpnU07XG+mWA65QyGNeh6ucbl9p0ntK+n9
QlwtF1ioBvjw1AsKMWIs3dLVGpjJulHZL6ZpbJGJRabE3czfPq6285OGTotZBW2v
caXz6/WEXuwV5VfCGRr9cbgKl8BAcE4htKyiTvEstF05y1Af3gOX9PARhTZemfkc
T/3bApR3EqRsGM+0EZVVHKY9OrhHoNwpUV3O0sA/AiTyZZEH8ZjiAZVC+yekiuem
AOj6IXgSAebD3Y0kb61tRNHO69WMjQ3kL3LspUgkqt09E+KUM83vQXAoPF/dYast
DfGmXnzRmet32yz/t4wILDqdHI3nf/2GGRRNuHPMoFVFfi/UGbGQgBOO2jr+cAvT
+sNTAQgHbCTpCWleLhovU/cpWHFPQl4sZJcQRLjQyQ7CwpLKOom+8LkrpUHCk9uU
kFBleMvEmDrRCh9FEZ2bznEKR+rUNa1I3RxRxFgxlx5uM3lKgnJwz0SQwPa44dg0
F8DchuI3Dh8YdMZTChwoIRk3RVv3Z1/De1kaF261fDfJQqRxcU1+nFk3uUhVwr4X
1gqv2WKgM9dgFcNicNywJOo29imyj/1julDcPSLI7VNhNtPWmNb95qDTWefBljBV
nqlAgM8nPHNRrHJTpqR/mtkbewQKBoeQmqJ+++CjUz+dgzjTCox0WEP5QefPkwKY
sb5Kpqqc6MrUhVyYohFDrHNUzTX82tvhNcdXrj7ecnj48xyGzv8ir4h476LTypJN
nBQE1D1ws/nDaIV50bYlza5Ot22Wr2e55aJfm0TW2QktopreN7dCfMnO1p7X9x6t
HcUdJZUOSkCtFFBTUceSZw2v60s3jS932Jsj3bUOglsH+imlhTMA1W8HU4vhQsXD
AOh+s0SqygED7e/I9m2WC3DEtztXKctftBvPvXuAMeE3dFrcbHktCnL5VYol51Jn
Qd4Pl5gEGN3ImQ0wXflyuEEss4cLBO6PDcfDEYVNRYuQcqMR0F69ypcjRXPRjkWD
hkOSr5HH3YNhrAhRwHcc11p+p4t25KroYhK9jeIU27FrNQbxPP79ciro5QU8SpMP
uAeLnuaDCxWg5yE5xpS3HuaTBo2OkSt8GNiyOF/8pu8tJgAc+Bge5thdNKmEuDgt
p5CtLQJ4TbXxnI7bupYKkw3Acfgey8utxQK6R527koVrd3jq2F88QvTp6PD9nKI5
/dhtoRp0iRGV5o0W4ryiaxcx3IWBvSBBjPdRHCiC+kj8rmJbc6PF2oo0Xz6sIDOg
af/5+IJeYJSsaayNMdGEjv/sPngfKtTka8bcwdVC/Z3uJGoiWZUrxs0RlLZxRSPF
gNaFYayS4tQN2phk80ZWVu9D2O4rGWxCFuw7n2N07qfBaemK1m8sfBiIStDZW7cJ
4SLfU2P1eQe1rdohlH/PcLOmXoyPCSZ1N+auZffnF2zU1TZTY9k3zVtjdJjj+p5V
/jV4hPqvmUxqU1Jhz42gpBoLfnmHlyBrJc5/nnWPeC49UO7lErObrVO7XdT5gurG
kcs+XZDDZGZo8ZHPBBA2mZ7rM1yDmOgrDhtv3h5YmuheHdBlq4HmsdiWgeQgpfl8
av3Gev9L/K6+7TAAYtCkh0+9bnFPnZJKtfZ82p1TEDHV5qYYSvCPFwAwmlEAgjkK
sUHuCmQzBuqHeLINt5sRu8zOg0/+PADiQOl31HHqUGYZmaLQvseei9zDEcjXqp/c
E74F5tfzfWPn/TFLIiNibwFXRB8qLlkishO5glbjWF2nfN0GAq+wd6/zAZ88x65i
l7JLxSWwtteSOhG9wXtSV+sptNabjA1VqGPkylaU/1/opSbcXbbPoifUDPhtl5+l
7DNclCVORnrBOqAvGZkPNvonARBKf//G1C/OJ60+mHnEnokCCQk+9deEcUc/oJvX
wLh72lhEQ/2gU5t3/De6R4fdxUmd7n7p1MpKPpdnd5v2ZyMPuXIhs1EvKMCQFP2/
SNh66H38P0uP595tsOthvXb9dW3SkDNrFWoxKar6QcbXAAUOy6m1Xt4CZGhTkM7g
9LksA6uyHjj53WwFrrSMGZGe1//mVTCwvhUyh7SPxw6UEZo1DRk7uvbDl4XbrBre
+uelqm4KP0o2JmAnugYL/Oi2MKpJXFWsEoeiJ/LrHPS6234YIOWio5RubyNITSAD
0Z0SKgdzTHx45hO0QYH/ZNrOfS2tcmYSBfBi3/m1J2irOWCOHAac9aE3VVL60JG2
5EV2B03wwmkOmqoiB8MojZTn/tqr6gPUQUKK7WB/wyp5th6AYW2MKSQAQmd5NVyS
aprCgbL8/SjWBCJc56DhxkpiRBGbGqz9SIOaDuQbvL4wiovdaY6+v0kWlgWwc8s9
DS04YltBHTRuhcAXPnbewlVycfdondsk6g2qHZ/41nl4hqwETEpYlDLnSk+Hb7m3
hTvjiR+5f4PXVgw3Z3HMlRRUFBUEdsd+RYjdI2jJs1j+yb1DzszHBubVnR4hYsUJ
H7Z1d3nHKnzoboJV+L4QhwQl2LpCs8KifsuRJZVjP3o62h21UVHhkgGmXiGbqyK5
TZ1CINHSmLKfCXhNGpxXbACtYp3QWsvB7xBXkfjrN4c6rmfHD3c5iuSsFZUJzW4P
mqaAvDHukr8+x+YgBylqWyNNZllbu+k73BcREJ1zt/AQvArna4ZGGBOdAnZqFnM4
gVocSI07DDqnO6I+yQMpIxRhE+4R7wzAvNkWdj2+b87i/6IJNwENgpz9TPOGtsDL
EKVn2z8zc7fFAR/K2jukwpEzY+KoYbHDwMLePxTQhhkJckN0IAfGwjE2ag2mNXrp
tNS7XqASJyjU4IC98FnvvQDXrhMTNKLMswjDMpbfvWUMiGno/1Fy+U5JkykwEanG
De+wzjYP9u7X0K9ruq/2ebW0Q9bSdEtfIR4jpQT277jlqd2Z+6EsJaBVfr3Qg5Fr
XFhQwQDJRPopMJ9Fpx+L3GaiY4wwvy2LVAgaF49YG00Lypsj0j4dreS1JuYcxYzX
qDZqWa/Lvi904JiYX3qcX3LrCdXvQ2ISQsb+ssJW82jG9vkQNsSH6Wi37buJAkst
P4qV6cbYtfwWaBqPL37cBUvL8OklqJt/jZVazIKRM0e3c2XERFnTggeqCMOw7qUZ
dNOCj0p8w/ep2HheYGQ1s06mjae8fgwM8Ezh6zJcJhYPpG157cjMlRWEY8U/cjSk
zOYbGUvBqycezLtLAo6dx8U2VdZnfVAG9QH4xua/fagAXwB+R1E/B+Msldp8nUJA
j1blWe1VHv3bXRCkV7Xx/1YqUFDwLq+NHfr1fyYtcHeOut4QmYEvqWthRtzUkBwP
oveNvSPMbW0k/c2R0cc1X8T6UNLjOBv4o2Es3a4i9MWLEgRbtlrWXfvnBUB4JPv1
SOhWwabETLxsKyPZEQhE0OVHn9VgilTcPydQi4GvghGEjLPGC59+PiNhzjSPfysM
Soo7ZlUhUGajZ87mBQ4qeLtekVXT0e0hDNpIvsdQm3Ou2+xr3sHC0AlfIIcN3q7P
j7baQm8FDQXfUpeLIZViZbOkm0pstMQYKTu2twoLV2cVnb8hoq7rKmGb7DXyuroW
brPz+VQTrULjWr47AvXBFhLWiPE/5lqaZsgLfKtXlFZBQLB1NwuQpzewWtJNZWOZ
vv5KrQeKGSvrV4SlBi+7KyDh0XPAGdftZic03NCjsZnsTFlxwFgOFXCJYdmY65zC
z76JhhmMnVMYeu47wmVesBYiCmrGSwRHLg0Jd3ywi150zAeaxqj9zYkr8bGj12Nr
y0Ak2Hna/dSh2RLgX7BdqWVfcxoQBQbClEkTOveUDsWdyT4EjXcC2I5E1L7AvsQp
FOmi9zQq+4Ln0VlHGg7AAeDkaydLkMqEi8dcdq/OkjTrsHIkpzVXd2Cs5a9Npuue
STsBsWYBPl/SWPusWU9/nWC2oscw2BEKE90NNLhXC8toVGDUe3RLHVSnHcKvthng
PRMHS2qw8TgV5O6lcf0dvf0qETIRdlIx7uPgXWLJrHQjdDJ7Am1lyZaRoXJCR1t6
vQWvwpGAM5TojXntdgSfcUts3ci4c1IEQvji/tUh5j4VQoAHpcEn0fnYZ9IrWSp2
VOFvJaAnlwBGgEm1JJLV3pRbsctXsN6cHtRco8aB+QIYxhFBTJtBNZ9G1PwY1AJf
MaxBBFny40RRpj6eUarP7a1aFy9TuW5UMEX1GSek6WrB2MKaXySOAzLw21RhlDrN
M8wsrCl0vagc6cG4lSz4j9pye/lKVg75X/nO4Z1FLJItLhA9TbIGFvavgZgcaBXL
P7KDOx9JMPl1wx4fwKgTvOdGNT2Y4AcBx+ets+t+4TKhHFm32sDwz+jTcgLHmTYp
RYSAG4XPCNSSKOwyVVqKch5Vh2mipin170M9ijzb4DyEzDkwVyK8BBGIjdnKUHgr
GH+beqOVBsKUqQgT502i0LuV95TOxdZN5oKeSmIhqV6DL1ubC7nkON2PZ2xvVNBV
qgFoUNmISLkgF3MhIb1G/68S+O3pVqOE9WCbo4BaCVxiKB3HQwZF6U6Yo9JAWXS8
gCH6SNgLRr/qmCDvltc1LD2CBdn8Nm1LZ6tYcVl/kCDpzqAkQv4Aq80zWXjtdTaS
xsLoJVkpN5AJ2fLBmVcIt/tP6Vg8TGS1Qk2dWjcnwUwWbK6kpajGuxfjXbNaiQ/8
hJJliWmt+NLehSLivaDuwOzxsMgBZPcXXjT/4okXQCDnWRGsTxXGbAtlnBoErFbl
KgCTt/i5dVRK+JUC2dQHxAuSctMKY4gQEJ/Gjw/OQ3NXmHlJq9pYOJjJ36KBjcZl
RCH4JGH9LHlv20g4JSunQ2a7A13pJOJiuXQuKXBe8E47STF9p4S/fFYiWILeoSgw
hpSanUPFTzDfs0lokyoOT8sDgo2vATjfxKP9qG7mNmQCuWtkGfcZrJCG2/h0EUDI
AnhUQIBsJYIWTebFBBbQ6J4jCnFajkWin8Rf/uJiJm6+wzw19uYPwTciVODH6/UV
5UJWY2OWkFd1AhxclSQfTKc+FeghSEFx+vOtuhlwlMyfvsRUQVp5xo0JC+PR1fZp
p5G02oGY81s5fQHjTZ6MW3QijBW2x+FnnT2x+pEXuoGYMg258oMgGs8cKOcu7rcv
0X5KahXg0NywNE9MPQLm2i3V3qD0vVoVizyKvZr8AzjwYpablVfJDXmhBwsQJi2/
iIU22tHFrP/1MsjDGYennqAyauRlCOUcU13bvRVbtKXBGaK1q3YWV+HM7SoH9Dxm
+rqWJjxAKWTdn+okC+sj6CrISGvkB/GKWkzr6bocqRUnWs3wBulaVEK+pLPNDJET
lB3pptfnEIqzNRYOrsgxdlc0ijN1QIOK1/xEBlunEjdLA385wEPuqtdeXb6IAfEd
sJBtZ58J791VEWAeGlO8RvY9MfPGayiRlxmwmcknyEtzuoJUHh1fjq+K+gSQA6N4
KjqtJTALcIWZmknsMsWqAezrQhFmbmYMl/s3Y/YRDtlEjxT/H4oTxKg0n62qoRuv
uudqUTUi6o6pdgVKBO7s/gZBpc5uzE4J99akygELIKgiFbam+6WAFaZWjDDQYjKB
L4fssQXeZb4v2B6uzmEzsyFXaNwjc7gK94Ae/YTosuKt3v9cIG20Ob+mYjilpPD/
6txixNm91LfOqy2mbj/SdYnnhwsWLvSwO0CjHHVWyB4nTs7pDIOAokAiy1+W8BUs
SefA6wkvJjODI9I1j8xCEKpjeU3haQsRn9hmVceKeswjfESIz4JnL5Vu/P6o4INx
gKv+mO+HaQ7UQlE5YkAiWCc9j5zASOA3x5a3lihEffA8tBfwVkLCJQWA7X9b9dDQ
9WueJZwGNmczWyc/i47o18XAeWgpJeO2tLRrq6MEjf74P0kBd39aUdqHkrsaagUl
04tEXksnZdkrzfdAlArR7U20wR3znHS7fgQd6QJ2edTIy6P2+WuUeY0aGkPBGm9i
Kbw+ARNBIpDkLpu9qL3TzMDBTneo4TlUy04b4yhW1qKxBE29R0Pz+1V+uNKLIO4g
BC2OFR+gUcYTt9wCpqJgtzdSN83DEJz8MoT9kNE0+ABpPO2CQHDNLDzWrbKBfDsi
Rd2On+hMsRBxw9WL1VzzRq3HO+vxlU9DYH8RtYEj6IN7HfnMD/V6Jz2XYcsnqte8
52dvjFM02msNEjUPWTXmXgvuj5U/EMvbUoFzFSa6XKwisL9RvAQPUAsVmEu93Oxd
dnMkKuTd+jojtok/Sv3rovNE1F1CaHgSrPcMW/bamtTbEVupfTqXJUqjtUrioP+v
urD4PcSPcaGskPJV38HxBC/6ott9GvW2lmqDyB2T56MLuMKtsya8ECkPYxeeYdYS
qlQGTRprz00bOUcMn00IXV0UChGRokjU+GT5nwdzoAPBRF9eztUnb+PTdIr7u2wz
emRmUeg7eNNzs/+BY+N55bhVG5pNWTftaBOVhDq24kRpoFuEG4vVRAJQ1eqijXRw
5XVZWmetPa7I8/j4Qp0uaiXEeMBCL3myBwZgIgedHt1ufYpznReoqb2Ye7xjz8hY
Aw/pHBXLKuu1N9MJWYgPgoUsATiaB+bNGRvnKQw4HG5OX/sRTM9SMqkxwkia2d9Z
7DE1/zlE5L1XyuPeA5maiNJTGwwf1brwk3Rx+aQAqi+BIN08Ps6nVk1ePTEzW2dB
lZfoDIhkklHXfedZAWdIxxSIBRKtJyDGa5rENGwDjk5/zr6Z0wxqZG9kVbfNkDLL
ze1LtAoUhbXkkerOcfvpnIduBzozo0KVc98VDre5JEk3PdTV64q0bB0AM6dxe0Fb
vTTzS/D3qmYJziuz8Z2BhbPhCS4DjvtRGt0MhHRS7xMGTP+HrcJKHC/jkxLBtwdr
VJ/zpB6nKZKSXqtc0olbirglZJ6Hq0CVm9tT/N9KZNoI88TRa5ABTwoxr/qnvGzo
CZxjBkeQnEus+o5/lSIycKiFsDPuWD80OMjQCO9zyh3sY1SkPZBamxDWvZ4K2gHt
qUWBcy2ic1Md5PaHpPDL1eyqCz/6uHCWFHSuE8CYWL4ihyHj2KsCb5uEpI5UMH2D
1nqbsbj/X6qLrE2H74UcvJvZgYlc8yTqvmnPBFVWzyhMnX6u1D1pzGvTZo5dWxci
C7nJjULyL7EWgghtPi9xFxXahN/JZ4G/7T5ev9xO3g+Du0ZkSn97REq0gCV8Le3x
mZqqMQIIa8bA0695UkD5G4JGBkb3plnX8IOw2JU4EbcXmRgcEzmIM2NEhz32UAT4
Zf91wst7C8bq0BJt+aMjz+lGoPXKswPHVPuqD083aEr//zGVMqhBy7PG5C0Kxx13
WdJmRykJlrwDtDZM2/8tlqzKhzp4r9GwU3ThrC2VRSz2ekD3gxrvhVRhPuRhnetD
1/gqYLwe+NUB0hb2d4e8EPme6WMd/oGJS6F3ykO164/ymMd+QtZEGa73mEL/8mch
b1VjHCvd/o3SMiZIb472XVNO0XKHVj+VvkYzgWFfYVwzL3Rtml3cGL1ZwtJVgdgQ
aNWUC1yVKnhHzB37dk/SA9M0wuQc1m+aVVX3LPFnADeYG/70HKL3Xv4yKF8yiSIH
edfINDHupaEM1bznJzfpKIurBeXNJ3bhOVIzpfceZM+oZfmmgBfeVX+3UPgrJT5c
33KLZZKxiDuTqvgKI0m0UlWAdEV0fy4lUKSDS4DAN4afkv/Lz3CwD/ShddFFUcWB
Ls0vj9PQR1mF0Bsxvrd14oARm29pFWe/T0rOZ2F+pwWuCqxaMIlzC+DxyEyWbWQB
dVQVbMt+y5r18++Sr2anUg1HspzeYiiMPKpq6vzoMKLM2WjSzV9ttODmzLpdxedh
59uc0GaW0haNbGUkZROuFROLPw0lfgU5C5bZl2pW4+LcrCwZUtldjn7ML3+XWbrQ
kKHzuoTdSwPd2Vhwpk6t2xQ5p/WqWsC/YiGEXPWN+e+31Al13zSMUruBNyLw/Gx3
ZLTrYBDQ7l0zGytUOnaEtVIZJBB34MhGGzk4hgCp8esvP9+Xh1CPX5mF4DugvmAW
j8Sh9JtiqU1zoa7SdVPrsS/v3CZCf2DAZn64GdMP0bxwoA7y7qNThoEjsffQjfhY
gAKqxlwmDIH179dnUpqTBn9RJiu+pMPVexZHfTHVBPP0xb2G1b0FIEhc/Y75mCv7
5IM6eQ6+pu8WCA8b8626tE6VN+UH7p+Lf7FiZPXy8N2AOfG6ornc1V3ZNpwKXP1+
fRPnjFFSK3kmmGi9vIoI33sw8jyu595C7eYxu4s5QD7Q3ch2VAwsk8Zp23W7uiwa
vbd622l+qI3w8CpUdwSBUrsmrONUXHgLyjNp3kHDEialzQ+scE6WncrYZYKBqi71
28lMftzA6j25fA1ZHnDQpNDzmvPd5qbU8aT1wKK7M23WA7DkP3f8vI6AY6iZPZBP
bjTA74yqRjbnlUBVRl0HyRxBj6/gtGOCcDiy6S4cHRa9kg0WnvppeMFCj+Q+LdGm
cFirJeiqbg8FXwFeGFLoY5EcUzSheWhEU4wPdkevX0OH3fjUN2ZGBAuX6nJ481w3
JMEhZgBF+r5ZnY17bhDt35pVoTku75frVKfziQ8mY9yg9sRgoXEK7UgXEe68qmuv
/B/U2/e7/hYq8X5CBUAI4fIBXJ5ABL0+2HGlunt+isksa+2SnaHamrs0ByX/Lycg
aRTr5+lFmZ494lcSeLXY5uCkmoWsgHMrNN7Z+f2Hz6cSNYQv5aaOsG4qnyLtMwEs
V3Bg/95NWyXksUHMs1+Khr5Kq3bapxCpyIdwjsNrK2CL5PNPe518vQB22ls4VZ5G
gpVeNPdezcn+lG3Rqn+5vwizTYFw0kDQpSDggr2iboowAKV5WHoqtBsh4VrLYAJa
uQ+Qm6P7wK+e2cNm5J8LmXf9wut9B2RYCzETXvHgewL0+fjxSK0iOqApF+OEMHMI
CE3y9YpTo1gsQrC76uf/XPyzOFcGGnq9UUwWaBWU8jYL6eAKoMUfceCcKCHnkDIY
4nK+WUyulFXN/bFDHJAEWjaLJqccrHRf8+M+BQ7OviXoOOZVKmeAURo7PLEOtz7y
tn3LzxASkWBOYbFictgwS6g+TtIhMHqZsxsiRsEk4Zv8v+tiMG0NxEkgVXRLWrCk
dqWhpXhYTeu6Ir4Cm89gD/6h+bDSJ+WzQ/xIIsIdC7Gv2Tp1eJ19yZE/9AMEcxmQ
HINj0TH+G90Q0VljrRWYQuT48/HpVRiBi5fdmpv/7B/Tp5lAixvZ02SX0IH/NzWs
jv9v4+2U+dPx45ahUvFtQTbU2nVctL26wqifWgAVSjIzfohNPqFWPNpz7G22KWmP
XKikQHu/npRjEiH5/VNmv3XaErA1gJqKCM98JoDVi6lfz442EkTDm37iGfGno9ew
/TDs3kC88eMNU/1QAFkHcJZgF1YmvV4YYNwgEAjvrKXnXAOupFATff5/kr5iQVkR
qnocA2FxGiOKfkbz69CpqSEbqzeRdZRsycGG69vcVLHKrWXHpe7dsbvrUCz5yu5b
S/TGkPUyY3Hw0BXINpdF7KOxeyUAdMTt//AqZbysDZrIadkfEb85sIzzrfl1FaBV
HGEIg18MjglH9Y9AO4jukIkvBUTL1Y09dreudUQSLL6tL6ZBIpsFKJNkFajSiMW4
4hwQnMGTT1M0dnn/QSM4WjDUf3PDcRz2St+j7ww0J/eiZ/nNBTdpN4pTMFRWPlK3
pnlnYUgSTcrU6+VXreFVBDorSCW8zTThW7aFXn0fa39Blksl88CfGKNmwUA4w2bY
kjTqUxignZpSgbCYBP70hERFeFXvzUfOgto64JK+G4ElrDKl7lIgVb3qOoIIls6w
jBa9zUm1hvZfYU7b3l31JkYBnMUjsEXKNh3sM3mywcpmCTYSOaGoiTUVojn0rgaB
tFv+308fvWhRyMh4ja3qYjExfiKeuihQBsXLzLRM1Yt5qmEPjuzdH0E7IN1KV3X9
3rEzdRPy2zWYPYodJMEu0lcyX7cI5cFqAF7lWF1tMoG7d2SDbkpBqnhUEFsiHFt4
7+kqv9dTOB2JMNfYp+tZApHhPeE3lrXOiORluW/mqhzMqCJSG1gj2svPqzQVoOuA
KIYS3+OsQiBHOI9vlvV/VPly8VPunOaeYjPJrcDvOGyIGIf2wR3SCCMx5xW165Ve
OrjK0AuL8z5GTmR+pkPd/dqn8gwUXFc1httz27lNHZCW2mE+M0LWJkR/6pRqydiA
qWf9cBzK2W0ClX0/vJqi4Rr0A0dgiBOn8an2kC8jZgZ68ZgC8pMc7fjNDiSysIF2
6qKV+d4VKcS3QhSIXMsTARdCdve6wY6BHSfX0lzMADeoXYGXwrRxs+cE3Kr0CYOP
PTtDMAcZGQBnXx3beZbo+olfybPT9NzqyGoCApLVJ/AC2fU4KB7djD8Q12sH0Bm/
mXdqP8AoI9OA8LUISZCz705ovoK0ua4Q7pTzVXx0gicoksqF7JyBaD52KEzZOi0E
thE8CmGuBFC81hzos+EYJIlG3o8re/AIfvo0dVx1Sn1kUF5V62gLBT0L4HydU1al
jSRbgZhtSEIfL+UlymYYNeEIwkmauqBYBaH4xqhywqTFnjXuIfAsr97L33TjwjB1
+W1uC9hZKAiwIsGtsacGRGzSIrkdBDbDJzZF0JxmLTt6hwta7iBsMcAPww0kCeJa
7B2/xNo8YoHD0AGILq6cLzgExWKN2tXJZciZL0tFVLI0ZIX9zjRhN9KMpGmYW0Xf
IW0/wdV6TA4AlrzxK9Z4J0FYuTEkGGEq/kjwVMfdRKGeVHXonz2T3Ud9YLIvFUew
qZF6GPkmdl/JDDo4xVSujySGbWqx1FX/vusJst82houQuIiPzX0T+Wrn+zMPs8u1
4YiDx5kj0y0qXqjU9FRmJmFaDThO7fcfVJhqqBLnB7mghoeiatDsNJ2mrdTvL+sQ
ppLlvJ+eMZpdEiibzrlLjPfkM/MYIfpbN2jUHDsIyvC+quGOnWPT5EYBxz1azj6v
nFT43fFCevYmpXhz2vwTqdHHInS/2kVS3NCMXvIwN6CjPkXTrzOgR2uLsy9WEHYT
gb/mXwL0qiK9yb7+6V0W7uRWyyoYij2KckJ5F8JbEyNJQx52QdbARI+vVbXHEKa0
UughBQPNiEiU6BVVtrhdR8q9GPduuZaDRMcogQFm+1HZMNOj39G5ckdDxPH8aaaO
Au7VsggkAYXBRb73oI0gizNIkxJloSQN44QjjjMOMvfMzkfiPPw8zf9VaqJtcksE
nbZZgE4QoHROjTdmh8TXWMIqQedAF9CSxuB8jkJZU+C1ftKYwX++2tBQVfNMK+1j
lcpeejSfD6xjKLLiWDUdrZF4QbCwP2lmDqmrS42Mbx2rn7Y3pu5nJiH43WA2YPIX
wNzsuyktFHGescLLXOUSbERT+WtbCvE9RcRTx2NRVIZ9zX0vhxAOtgmXjgYHqZGs
MVTbk5HRGTqNfAUcWcDfYB2cOBBaXlDVKAgaIkpPYWWgg2I4YozsTuZbCGUl2no1
EmDqMpUcl4rlQn0nwjDuhL0AXsklvV6HeBFD70FyHE+0FxDucwp3UKd/Mat9lHHU
Ps0Fh4edznBwc4wm/5XR6I2JLFSU+b+OoaAMmf1ra+exEC4nuUgaM4zl4y+eIpox
xiAo44I6uWTWmfF+biWtb5fizGnJ/Hc22KI+Lpr5dWH9U3sspsXinWeepoV5NNHj
uhuSuCTHZeDK76AxXAQlZO3xeBrptJfr50lgkUWoChEsCYaQ53a/aTeBBYpUGWPm
AwEzkEybxAWstesZKxYgDhzmEQLMy4IKk3UGTHwk+vNBhzayGbfhbsGYa6GIuPsx
OVaj3/jQvA8Lc4LgclJs86w9VBNyRUOS5AUnEIVe/iPLR6NjkdumOiB3BJdjVSLl
3zbLEm/cEQj5a2QE4aqpWtVBstrRJYuqdVMOzVAg3aBhyz0tKw0e3zYykQ/T/B1l
J8Na94UBbz8VeLqn73IMNnBGFAyk/g184dApwZtxHbfMHPFcILj/K6WfR0ut+UsW
LFv5lM5VyorpHy2P5j0SITpuWMtxQyP4gcJ4jiJ37FHzxSfjqP6KHrQG7URlU1zu
o7BQcp6tqRa9R58I256Y3/q2x8DKVjc7m25WiDZYC+GgwnbvzvgcizkycBJfYJ/9
zZSJW+q/59AiQeZWY3l5IT7LcdwyAZMNaIxw9QmsdZiaupfU2Uj6uaOSGwxFV2HK
sYyi0NESktzQrEbow6YLOGRTDQ3r3dKvFObGM/8tneE82ErBPV+mdt/y5jRa/Lyk
5APZuyqrtHAhcMt7wO/EfJ37lUL99ioVO28beG0DkT7VgnZrJWULYCn4mcLwHk8K
StS9rbEWAnG4cn4uUIuhGw/KhWb2DkTTOa3PAMHdDTRo3Spmz4w5gU+pzsULrWw7
LnzssckITt9jLzA4FitEwVLhBkIfUiw8Argpc1k0vcJv9OlkZGlD2fpcVIMjnOgg
z3XVspxragVOCqbbudjJLeIE8huhyEJuC44inZMS1lSnGGML0tB7eUD7JmQWfhPc
nnrPBG+qhCsQnHMBJdPBT50gwuS/5KuFOfU8sUsDv7nKYI8zcANh0w6xtqh4e6t8
KswclExgCxa5lX9jTm1fnLbVw1RKVeDAx67b/xCrTLWI0KPzrBLR/VMQfeac/xGy
WM1wjGpj+TDvw1BzcrNAIBCtfmRmFRZDvPoxuriGNpSOeex4aYVh6BZ/JdeHqH+y
bkwtopM14sFbR1/u0zBpAGXdb4R1V423TnduBigwemmfSrWctO/znZNTMBwQiiPs
xEx3z+bPAX4o6nZxr9dQriXUep5bIYrmy9TxRuWMF6qFF8Rfu/xNNHMpKcek3EuX
wJgmwDKUZ5dlTchEinalqI4cGSunU+S46aKVCrNcST3ZxQorMaD9Unn3fDZYHUqP
ZgoUaY4IgowzpsH0mh0GXNVuxWWfmdxr3f5072Fv8nFwaPR3UG4Yux4l6HWbwLtx
2h4/Mf02u4+zYP5sOCbbgxOaTKWLEiaPuSdPdYLEUw08YxSdy2TwatUv5eZl39j3
ojggK3X+0S/FvCXN9eY5xOW7U6l9MY5t5g0Zq1BSkj5eU1TqLCVA8BXpqsJtxGpz
EPF7y8jgMpG3rBFggQoGmhbbZG+v369h3OogkZGOJ0JxfYTrtdjkXpKGqjpUQUPf
Wv/fqrrZW5tEBBTuJj3NaGT+Zco4y1qjuvgiFLMaIBl/efUmfdvhgfum6zB7VWi8
aMTUCnG+aJ1mCBzmJmkE9Hg57P1Xrxj/M4dXMsvBhy/HmW7gKaJySLsE8JxRv7o/
8J8wd2UULJl9QvMu5YC/+z6JV2xkuRacyDnsFKAKaLnkna88T6pHKA+KNL22bFZn
aqzS946Me2PmdurAzL9DAqHclLnsrQq3a+42t6YwngJuyCFq19O2859TOTQfHcYJ
7WKENZ1GqZ1jeKmmOXH66EO6QAr3USr1KJfhbIISje6B6UlACadDOf5kofjJwe4l
n5aNgpJa3LqkZtDLSN574LA+xAR7fuzn/dzFWNRU8pWvpU9M24a7/ruWS+qRATxe
1d/EukArScZDavzA1Fo8DNeXP7u0fZWp+CvSvi45IfAgay6v8Dv3/+zeLuFMjyzW
a0HVFx+Y0jTJhyOGo4XhPWcfnVsKxtJFX16V0wDzFDr3NaBKTtG6JJS26xofGkBp
t/ddv3F00oQOordr0k4xGj5GcChq4HSOHhoetRWoVzf9RfpXJY+ZlAfjeeUuY4Di
Mk+usfEiiWjG+FmXZ8zQeQrk9NDMkyUEhiOMDX0NeFFiPiFU3//WwwVYz2DnJvHA
G8vJ9qi7vMx1AjOLTHMhhJlMNhOxoWwE3rUV1iYUM6Utx6jFtllNzhISvlZZml4k
zByqQaoojmD9AaBYS3NEdPq6/v5idAFZTRMa7VWa2pY/i8TlaiR3wxpLbbU3ARes
pe8PNPPp996c2ZTEkqdKQkjLW9uiWI8x/I7sTM1wS1SNJYA09SDBCVBkec/FNnY0
OBbYfSq19VtPve99Ygb3v5dLCvnl5QX1qQTlQ+w5ltAIsDHLHSHvvaEHAmB+KakO
sHAlXWfLDw58qlWrMrGGshNKHvjGsMIlkdAqousk3vAl+Xs8RsvEYW8s9kBf4eBs
VGRtuw92ZJsV4WVDnr0s/kEERvdcOgfn71gvSeClwvdyDKOapGD30OQauwgXcZnL
sNAAT/UbRc1sh/5wS3hM1N9HqTktHCvXEuaPWRKDADW41UTkeL0Z79W3BDCaXmW0
y3LmW6nRmG99j57hrTRAm9k7copeOsyG+ATSWZc2HwoRWamFTRj7KNWennOBPjAb
H/ELyAQVddC3JWN3EZy1MrYOWkmmrsU0SnNpMvckrpAsNOgPYJ+LNh8dRnRZklKn
nqFUI/jWv7xdazO3VPk3vpXeKAeXmW8hle7sV/ASwvSFYxjx7kUzs8L0O7DPx7yi
mpf4oy+dR9lNlTlRHZc8BH2Vz2tXesEug1DFN+n0Zp3cWN/UHK6hcVPKsKyTsyFO
GJJbJKggs2SHrEIyWotgZqPgih+lz/Lr0pIS60r8RMfh91pp4AfyUIRBqzJ4Iitk
1TUQFAPQhkoANEbIdc2HF7Nwy73phITmj6WGINCwX/u6w/Q5z9c/ZIkfKLfxxuY4
3UR6VKIbYIaQz3VkM9OMjUReOvCXyzotCCE5VFEdPQqXGZby2JxFgwbQGXHsIxiK
4qQTNjbc0m6205nReX4EwDOs9mZeSN7XDmShzRM+fHyPllYyVSmCRU9HliU0ZdI1
5nhZwZlqrqjx9ymIInTpeBi4NVFXkaes0JkRob/roGvVwBvXCcgMA2HNq3rhaIf/
HbAWTmKtXk0LzLpwtTb3OLgXEJ1x/guMeOUnGHqWNumf9ylCs0qMRf4bpsMCLUe4
BxBVjMrHaYXWPgplUsg8waxER9kCG64QRUUaNTJf0zvXcy+unhnHzj/6crEM7hhZ
ia65o43Ng7pqljSk+KKshhmDuWPndPEF7PuRhDoWNblBkb0wcMHZv4LYz4D65y8C
heUTW6aPRTo++YbgwJqD7icMR/qBuTXMZ8/+CU2rgsU886rSAqeAcyFpgukHr9U0
X0oNmEiHdbSpiowX7dWmwXjB1COmmin4wLG2EuTBOP6elu9NhIsOlsQuhP3CxKEN
3h2Z05sI8k19klXc6wTv1QzivdrBNHjjVJKJOaI0Fo0JQqy8OBwuhBS7kW+S8C+m
VqEg+wCFUeHbuuznO40kYDKrVAAZR+JqWatFb3dkVoXJsdgv/6RxE+EW6RRN+v8j
A3QhgOTH4WwFMmgM/H8ld0bRmEKVK3gasGaCnIyk1VFjwPqCsZAz7nV2PfVdRue+
WYTiG676CDgDDPf9GgdVGbVyO2ST2Xpz2GBFnCKB+w0Sjo0nTvEA6bEWNyLLK/YH
2GfK0XA0SleJAGQA3vNRuTwYElTQzOqRbZS4pqki5JNuXNhRRPLRYtCiLB5VBV5E
n82AN2ubRpCcPoIeOamJVgCjDE/CXKXmi8RzfN/x65+Z8lQUXvLV6W6PxoeroFq9
tEdl2ynBwZC4RnZ9PFy1j/sygQivrQgjczXgeIsOK/mpdYwswLlqlk4RPbdsfRtq
wu7IpCdyioaRuV3yw9qNOVM5kwGEnv29szbdb2gKT/0uT6sK57NEM5Wy3Eee/LvX
R5G8bVin3nnm0lwl5HQXW3/iamLgIOcVSpqWOgKPCtv2ep/qxdoB2UitsntB8cv+
lVDAmLlhJxAdyrbU8EDiKbyhe+u08dAWpVo44YcXErh+Rh/csQf3YZG5rNEHzbXv
c/Axhtiq5IwSYlfswDCmQO7p4X9wTvOmB0w1Kc16fazfmOIdUwilxzhDmbV0fYm1
3n0O3D58QreQO9a5xvjgvEz3j4eTv5+iDWpnWaDYuaz5JZOgf3wdQrTgTEDS7bzP
oXTyHf/0jsLjA9O2QLK6SvRj8f+fggFG6CAhRQzwuDcPezmpY+ArWk9Xtf2+a30X
dKq20WM4ZS0PbAGaOHhPTS/Jf5PcvnOaJN1dMUUlhqYSr+5kLa60Z5SgNH25C48e
1CIiNNkGlF+OMgGghDolhvsIvP01GISEs9GtY5Id+SbqWwIrhGYhiVmFiE7WZnrM
4yCssQ9ua32e047I5VNM7RrxPoPWVf+27Y7QftVqSe20tYqG4jNnNXPXb6Id/A5a
6D4jbaB/6rqHj3T3O5j22LjQpKsH0HNZe87rq63e4V5FBz6XLlxbqP6BTQ3GPJGc
UlBVN6ilkENdG+bsh6Lc8YjLO9SBGjJEVadJEtMXp22zCr77NM9tI5X3qPoj+JE/
gGGrFczgz6AjeuCMhYk0b3WBBYXGYxx5HOa1zo/Gf93f33Wh0wwVbB6JJinPlF4H
ziDL2K4A4PGf84W1zJPlDX0VxHFT7cz+h68Oy6x6xqcBIGGNJG5DjJL80BH3YPwf
QGpFjvaUSrq+rvN5Q0+kMoG1OfqJG3gCRTQ/gHFvwifrFWoA3ZAKYm3+ATCHk94W
W/9vHGb33wpPUqLAovMb+VS0lvrA2S3SOYlazNqJKMjVmRSMXKKj5cky1vg1SkhP
qp97dn4oiMZDIWOzMuvD/vfUjXlt4RJbLKygNy1lL9o655w9FeWz9270agtFALWQ
AQeW+mwEtB1tg45hXYp9vi2BMR3/bJrtOSjgralkeFi2LxWuILO0ZPM+qQTC8dq3
HseE22vEO12/Eu2yhJUpcXhmLLelupTwxilvuGK2BGaPtS60fODCWoRXLzUXbqO3
CYemzh1ZNMuQ+Bg+l482rUHhiu971vRrQNFF5UW9jWnkQpw8eDM3nwy5Sx9mUi+L
Y9dnOBG05wBx03YG35zu/HPlCFInsOR7J5yXnChfWm+VuseB3feotSQIVsA90XSM
IPbp8AU2KIZTFruGvNJU8sTF7Z3d7jzA71B8+J7Mv71HtQVct4X+iQUwFqxx34sM
QIW+Ne1SalRc5X5ld0Cu1XAotr/cuG8IpFSjEtxVC1hssndRw2jiT0UeOruI+reN
71BGMVqhUUg5nZBo9Q93/drOSNABnAA2w8zTgCb5vS0cDFks5ZgC9t1TVrfSH4L7
qat59u2KMoV7TjJDWjhYmzBDZH8WG6fLUuksJE2Y1JECKpHEEh2Vy4rVjqwa85LF
BFsmOSDmAzgPRfoAxnOd3FBU8vtXQJrOeeVUTrLCMQAoMO2Z5by9oy8vZE363oYE
8yRRWsb7BhUd69b20plroViVEbBkedScMszqFR0M1gwRIkmNjgZjaZOdKFf7tLO0
1dJh7IicmUxYeyUQ6b+nNLzfBWsznLKGfUp74NmFoawZwBc3FNYD4UCp7EtnNaIv
jU1v4G25m9UReom6hG/P0AFte24dAfNIRIdw3VMufzG+bea8NTzyX7+EXcspdCRr
pr4DENLxNd1sM6CfKwQi8wURic7OptR59YXQO0d4Re6vG6yELt4sXhsPgLa56EKd
bTiTNyNOaYzRdGRVkoLFBySiTPG/V8AkDv9kLzpSZiUryXPCptUvy/p8AKaPv9QZ
1q3DG8vDWcqH6IWQ2YIrw9KtOXCvL3qQG7xJUas9WD+6FkO4zzNEpsPm6Vji23Mo
WfVMG1JAd5Ar+e/oSF5LCSQF4i2orDqR4mfTjIG6AVCTlzpXEqCCAM48GbkAgad/
fzEJjpdoSLLBLkaRemon4pCFt0pgXdOCT5TcBPDR/agDaUeSDrepqXHty4Bz+uDZ
XvDTtpGius3Ku47SPx3JLh1egtR/JggnfMLdXM6rZ0rrqcBlATJdJFZHc3gRI1+v
qNruosn4hMAOcMW9Gx34XXl87StbQ5XLzMRsIeb1thahufQExLb5V9AK6HerNxR/
Dj2jluHw6iUD+y4HssJRe7qqRszTRG4MraRnfs0/pjjT+pXamkrBCD/9eaD1dBpF
VJTWfTetc70bNAvvQdXIdYbiK9vnp+EjGKImyee1cbdCWbfw58waH7hnRT/7Qc7h
93SmZm6zOsVr/jfwxVx3GMpUVjYpoxjevU1fg4/2UCfdP60p+UE8mgBqueAJJg1G
G3TGNnQAVKRwIlDziV6T5gtaqp5OZ24wCq3ziA7dgsjkQg5j83Aq4smvkN+4oAnJ
AQtWm86vNhRkEqRgLgCKoMQ8C4mC+JpHFP5MutbX1HhQUcFg6i06rBFMVtZP0C1i
bFkTrsrpefigvrXqrcfTrLLCvPPtv/Jg0ODwTcMhNTd5yjo0NptHFi+tN8mqn/vE
EN1pPZsn4C01pNANgOC1V2WrgPpH35BE7TGokYyGqYmL3gTWlgylTfeDei/CnR4w
tihTk9tTW/O6jjaGS5+MpoptHBJpgiXEU/CnW76jrhW2bjI5zYTbaM9F/vZRB0gn
1yeVliPVYu+nM//IazyLBpPMbpmVk4luWdiPD8cTWbFLJVZBUuvymiUioDjLvkNa
9XobsX1GH5xJZy4ejtm9GOPK3XomrIMk9+mThvvMUZmnYGFCwKwDobL005bpq5Zq
erEmKayF+w8iHLUf1HBvbKhiiKA2eOCUjsXLi9sd6yyY8vbrQJO44VSmM/gi8dVX
9+fqYgtjyZ81BruENDkQcHo0/7LKk7VoCr0ft3aGPf6UhLlM7XBL+gnXKVrfhZWz
VnfK/E7Po4sveevvDAzJt53vgE55GJFQ+YiG7znIqEp+KiFaLZKOJYtv4hqSDJon
NI+bxFgsPM5Rh1/lFX91f2OVsGNaisvLf6paSwR+mcaKH2Gx7jksN0NJshOLKHze
dT+IqbLetvoC4YyQvMlraEK2iFu3AUfssjPlL0GgySCKGQT9OeF5Pe1qQBmhkcYn
Ztp8xF4NqPIjLUGv6U1DIraV24rrLiFSsf40Qx7IKdZLy3EpzvSgJQrFvPh4llLz
/A08z7rkq/4TZAccddvKT8da85vLHgjLdzVx4ResFIPCRgNTdGvYy7LH8KLjQBF0
J4lqky8J2OJ/YElKBJiHpdSyFUwM2CS3cdXxFHWhYS/R6uRmmBmEQtRFBl2rr9wT
GRKX4nkVnnUj165+8M+Y4PqlZPEECTyNSgxXYVbP1wahHKDx/P0CUnTL3kdOz/UZ
xqcnBeJ7keMPJ/77fpfMFgcWzLRR0YEoJDpocpHo1jRWi0SprVInXwG2crsIUpAm
Hb/xiu1FeiMDFRcCXbqpGjehDwpy7NEY+7qFFkh7IVYXeZG5m1IJS4mroYD1tqg4
x2jaElpz8vJ6UNyHhDsuAQykBMja+dgwdb0yPXetQjYlLApVGrXUsgg71igzKHQt
U5plOf1UCF5wCs2hhDAAgNjze1hoFHNQoIgFe9YjFA3i1Bnr19XE/WwhVOzb8PA/
uYB34wBzuUkSESeP9T5qxWwOFx+6Dy/iZ+TIl1sHb/5/U62LecZjSKsinh+w2eww
s2EjMKdggJpnMi/TTT8pLHRBDv+Pwco1ET/hEXD1CmCev8NnUGb3K5DovMiPXdQl
r2gaXQJ8WAcBXAevHkt92PQuqHJnIpWm7jDk8DW/5GVKF8HHveB2aMWHjTMmrXeW
3UFtkXWlUctTmm3RQ6vpQBmscSX0REqvbpqfY6C/XJE/L/GYt0HDMAxhr3n2pnWs
evFnS+cHbYOitSwJHFqteJhPngbKd8m26uqYYjNzJLcQedlaxd+r8YPE2zts7fuR
TUrakOZoel2G4UM7EUf1o1C6KUSlcxmRWT8iXKudzN/Aj/ZGWzo4Q1KCbFpPQP98
XEP2ty8D3gYeTrWZQ+Viey95K2Y9aArbB/U/JwMM4kDifFaa51iUWsAaHO6hBJTI
F3HMuD7usK/biSLAuYBdCXBJqJXQisJ+zekmwl2jrFkPiUF+gMKX23eV4Kh4AsKX
gREzde5JZnBfk1Hb5hKSaz5Dzd5DomqdnUu2uP5wWx2w453oQVoUMkZFxaFvqJTN
inFcqqrMpBo95HeiXwR2Gankltm0866MuItlEbQjNNPIEDTM4ME/ASA/JCxGiRDX
aKOIDEGs4ow2L/fgK5ckRPi5S2VYoEnJ9MWzI/5F3GIzNkcAEvoS68CMJxK8NNSU
e8ms2P3xRovZZJ+bP8GrNcJbyejt0xsIT/uvUkSJP/TKZsgcv5j0WElaKsEwE3t1
gZ73h0vSYhwf7fmdx0yZHnSloLo7AUecIrIvKYhPDWb6H1PKtH6nIj7pvlFYKf5e
lD5NopACwlDaxGF1P8Zw7oazqguTzCqBrVcuZSnLNjw1NcHJh5uJkEGAdE6fQ3Tc
9WXH8ngJKctYsCCF7jROLFfVlt/U/6+5DbAghmWPn17CtVOV8MnbLgGL5ER4huSB
N7iSKW6Kd4Z8EyKVxtxmobCZLX4xu4mwqZI0YFXWmnZi3989jPGR6yfNq1UuXhbP
/EgD7/RtBxwjgMdechN2q/UaRczCNirCWXY8n5+qpWuR/ooNml+w82bvmT1CMjm2
bImQSAmFDfAPIKoueRmnlOAZnXL0FkQ+be1ZlklgUpy25gP5UurowvRPSHRgKQYj
fCEb1Ol8zz3O0YDU0TzcDUE9/7jLgiUUTuPsd7FFDolRfaIILEZUBaZJpUyp2zT9
LqumjRFlkmr0kgF84LHmh1LovJqj1iIv6C5CWA3NJ5JOvf96gV72PmlazKQRRFBO
SwCmB+lgAdzvY2GENXzQ6at+zfLUrG0erAnJ1tqx54RfI6kiNygej98fPG4xteYw
nmkuRMqGrQQdEiDUa5BybvWKg+5HWtuhgo4tC7FTAxUM6Y7+hG6RrbnaQJODdJSt
JWS3QJmG25Yas/jtlIyiEi4SZkbT7ygO2gXjyOAJb7k0YlqJdxoHXK/m/k+qVJv4
QIUBBNx6TiLJaMTaC/DQi0kNeVU4ylILJXqumHA353jcXLSqm0W5uFAoPd3phMeX
7Majup5cRsI/yqni65U8xH7f51p6i8kzJoVQzfohVGREMXnHfBB6Oxh3YbP8sDz0
6029cI7wF2L0S4V7w6nK0OoTIS3DWLr50OH6Xi3ABz/COZART9sLCzWyWA7j2naE
Ui4FLxo71y8uOhUp1+8rvgv9y75K/37HoKbOoM3iRAbofOM3nZw3E0HSmv19Onoh
0VETdxOmPjpFe4BBOjSRqpIlpJxfUe5DREMmMtu6TIOqS9GXuGC/XBrcvFLibOMT
PIMa/KuQbCmPRfTa1DfFPzALLQEr3iGf+xJW/xZMR9C9oWrmwxhNvtKOnKik0UHe
a4y5+XjLji2iZDJkcyDQ7QTp/mG2aYoJgFqPjxJ8mPgFOWoJXqyj0yHyGByKk1lr
rJfhfSITiHt07YUH4WIoXlos8qHilmjcwv1gyzLQ190vpYHs21iPfUYv/sQqLo/n
JJZpoB3SrFKz+/CYsNlU41X5y81hAhRj88qsgAaSJbr/XNpsSMzz5F8Kmzslqy7d
u/3Gy2LQqreOiR0yxXsqwkyfqa5jicr12Ve2TiZryeFzgNmRUuogWH8bS0baxqRx
rD+DzXw2NTAuWhvqqxZRCICCOtf2i4yqcyYzOLq61rFMxDPQuT/qdgGL9mAvCluZ
FHhNEXLEYXVF+EW6vDFCf5A5qsm/GL6CvlZLNDBN14I/U0hA5VnVz2UANAfr7TXZ
Nhe1ITGeEwmxBrz+uj5U9bKun5a6xcYcOdc/QkjWEUaRhJicdQC7buq/+Ax5DiJP
uyW7ilmL2XraMh62XqtCiNw+btXdftNzV5woOSrj5D4LBQetSjYZ7V69McqCiEqU
mRXqWZxsplSe3jEyRhtC4O+JjsW2PKBD+u6DJKoLgh1v3Tb/CJu4aSvtouKdh+P3
ayzQjV0AKF5iLY/7Ek5vuIYB1ZRRU/xCv8W++chjKDnu01c7YwW5/jJZtJE9GGR8
rnl06lC71PTFLhn6l4uw6WEr+hfbQ7QkFHhG1cpnAiyFTzCyuY9wZHixa31tNJOI
CC9sXvrxRaWMf1KzJ7C6u29sDXlZp9oPSHDl+OjMsI6tjbS46L/IxYfP4BTdVBWH
hFKeVw4hVjEQOHdC7UJkazZoDbTRv75WGh5wRiafcI94iE6MPj5xc0Ei56DpHpcu
IDZCkJ45pJHD62rEuI/Hiv8kAL3xZNeL0qCuOBEjOTc9xigLqg2WVA3/DYAamZar
akfrEouxSdHnxthFuWPryuCImIi8Xj/bpshRsHsa3tOD64tId7QK8Imeyf6hJ0zv
iyDXjQAmB3I2P0u99zctooRxpYv203649I3qI/zjw5by3v7FhQzIoM6MidwDQjQF
u0dBoPExFfo5sL/N+TUR0fg56t/Fcld/+iAep9unObqUVJ6s6OhUp/OHQSEGoLCM
vZENgpPNievAnqJB230lyQx5r+AvUem7eOx4EMygOdELutaaU0FP4A9go9C7mYFk
ikKZxwye7Zd+t5WVG+s+YOWJSolC+5kN7HWMKXCIqfDAhxr+MhmzNIJrlw1pVOYR
HuqDtwIVGHsbYDlrYBvqR6pnNgOHDEazKAJK7wp1XyZNbN5ZhSyBryPwgkqaqpAx
69ytSmTnF4Tq1n/WOntlUYr1geBd3oQHwIMoybBxch+P+s0wEvWiJKCP6Ppb4kxy
tzmF0UsoLuXWfsHn4+Eyg5S63aAkIVQvt4AE3JBiIrrB/6J+5F4Af6QGJ1P9690a
JF3eomf0I8GrZnhYig0zXv5UCMI4bByDoHADAebeqH/AOhv/FpeIzcRAaS7st5qo
Us9VkfHTARMAc8f3jCENr33CNdWU+PbbdbrgW59t5ACM/sq4cFHbx644PqR6gLlf
+jBHmzBFWJNdCJqdbwhQ7PNdl4FNC1Gg5cNqeCV3fRdQSK/I6kOxiVLbTApLeU2v
Ogvlmd+lD/x+TxaL9OqxQrOPXYAXi103rrdCimjvXMwok0LfGjVf7fjGJK45zWpq
2Nmnxca7jkiXkHwZ51NTuaeH9IvZUv5caeRaXgul6dXEMC/WIjMxTP+0gXs3MPP9
7aRzAtF65B6/LjcZ/92QaTcCtU17SB1zhLfwTKCr7bCogbjrBJmuSDN9Xcg96bIE
GtiG/iPlER1+XARZm9yj7e5qNYf/jNDLHKRAKh6fQW5NDF1sQesxfRIBhhxyUDZr
7kCC1ulKYhvPWP6ddjUmwrmCFsQ/vBmOepj7vRULFexlQriARDbtYLQrLRNw7YaJ
Ltk2SL/WdxUqi+TGTeRqmt7asxGfCgIfdK8ZVqkCHLGj1mazzi+zKOmEhIYtJH0X
jazUP+x0U/wZ2aS3bhns12aNjDy9DpB6io4uIwpRjhObvBMdQwETpjsFrTIPsRwZ
HHJgWE24lZC+0EYaZHwlKRwBr+MHVzwDVbTxeNG0duGEx21cWuS9yiRu7Ia3t2KB
OJUjglROEB5bVHCNSX9tgr7FUPa+ry74yTpjTwfzpzP318+PmuwVlAiDSFkLdo59
ZjMfQwHHKK0qfZKt2ZRLMwjDlcQWxQ8BhR5eOaLiJINZaliFsKobnB3XtwKkyFL1
sPA+yh2c3KYNV21Szq9ohovmUjmRdyLWX9O1mI5nUbZ+NSsO1ZlCcu7uJzNTwniz
Ek/hOtUhGGmBP1jsZbd62FVXBjMRytXnEi5RTHuS7PzFDnKeVMVF/b9QDVJccFos
f1/ZydDH76ISPwINtL2R6O4jnYC0lYXKxFw0MaX31j1kCslBUyKmnTQYol+53dNm
S+BR+jzITpjaDTAjnrgW0WuDobUvyhSV1UEtC1zRm3xIg0rqQO/xAYWHiLG1gror
kgIEanwxM6Zv9PQFh7/N031EqWe9GWlEd3pEya0W1SrOgQvEBpjckzAKzSBxSpfm
IxGI/eAiHEySbh1xYKblauGk54V/y7SCLZdQHnDjGhOet0PxD+v88r1sMXkCkZrQ
Ym9AsSBsCOwiL6xn3fp81lelmXSIhSCJKbp7Ghe2Z71OACE58Z3CAkUnjc5atT9o
0zOnlkSw75qhp5nec5qlpwED9u3C+8aI7jz734Yz6D+zPXYdV7sCd9oxx1mQypaH
G02ZdD2eQFBtdk+f1ezZsieJywUQJ01vHXdmGrgHuBMAZu01P/4vqbM0rzKsjaig
B4Ilp5H8zq3YDg/KPsNfSTZMC6rSpfkjUK0mezE8dJlWJaiz7Pnyo4NvP256AoG1
v6vxdlVP3ZxHvq7SmzbY4LeM5dhAL/RkYatqukH2dAEJLQ4gON+L+u6oWn6rU+M6
Rhq64GZI2kVJ7jpCSRuBkHtiFXPiCWj/BJld+C/PrxWRGyZ6J+znA7MMGvD88p9j
dagVeDYOe35JNDx0gBLNof5BIi9hXTRajpobCSUW/hQ1JxgcjJibzxQmoRbHYC6Q
zgwZsEA8hAbILpA6A+cfQ0r/dIsMlulYEg5XF6sXHH3B/weyRTFUISiF/Cpz7yne
xmX1ES31GqZPazMbUokrU9/U9J69y2gG7Nzdp2KwX2pAj1TLDfOQTXzgtFc0xsyY
mvEcss37WpSDvGcf9OBPgdcKGtewm7VXqqMQvdCBXPp9cYyLgsHO5UC6bwbF9H5l
2/9f4b3ppmQ/4fiHsD4g+Ej7Ri83/JEYxCyyb4Qv+WmwVpMvjV9IDNCwTTj3GJqX
cm3shT6GEb4AO3e6OX0cmbd19f+/18ZpM4SdxYGW/Gl2+a2XNdPv1uJSSCCGIqXU
`pragma protect end_protected
