// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kksUNWWJTBs5v7h3r7P74w+fO7KN/wkjjPD7dzsCbpErRtoQYLHuLoVBrg7AUw2X
wvTNYd65i/+PIoNt96zRWUsGReo/Axz2+WKj7JuqbkGIyxmdi3XCFU771+HJHA+5
5lfo67hVOYHPaIQ4HpfqLHCXyS5X+DKJi247N1ugjQc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29488)
PGhV1DLJ4fTc5nyj8pD2/9uaEcbqH845Z02m7Fw9KUcFxVz7YUAxff6vBqscbge8
Lo6BnUc1yNuCfCYm9wNiQlrR/5xc2CKY1l+HYWXCWu+A/f/bg5fLjiuwRPlVLurn
6wYlNG+HHdG59S69BcdtU1M9886GFWygZbw62d2dfSxVe9rdKkUa7VllBfdiwPmV
/7yjlFKeiB4EWHIqRUcKzqq5yn3e7H0n24HSo5hiI6uKVeJcoABdwKqR1Z4RHZ/6
muj2sEnovjJAeiF7BLfE1ZYuxtEKF5YkjhHlbREN1Jk2W6D89yrgy+ZyE+OIgoxu
geLjCO7gK84RgEJqiZgzX84OohMzvKOTK2YwDPP3BStYXBRdXDFk1gak00XIKWvM
1wAZcTlYNm8SnrRpxTabi6pK4Z8z5o7g9Yh+rjf6HDUCBkkkl7gvEkjIG5G8kiX3
/nWH254zFo5ChnASu69687C/X7lbZxw3emb9YEwKSVn9KxModGHjVgGz9pVSxfm7
j2t6t65an4OYDMUgXwn0eJungaVzfOwNvkiksbyKbMybzdOquq/iZ7UFyYPdeFhk
mJC5i1K/A7XRGZ9RVMuj8/7M+Uj1Z1CH6C/vhQgZmHAQDhixX7VO/bDy5WDnmFIb
BYMaASdJRUi2VxGygoy/75DCm80iYT/JAVsvkgUkNwhBmBGW8rjlBqB9iaNtg851
bRlOtVzPG+btRZB/UjEBZQLBlxyXgxXRAjXdlpeZDZ5BbJIOLiS1m3hwohUztDcI
K/cEiuCgm7l04Ov7NpQc3U83K3FEUMEirA8aKVbnEL1oLjB043u9RUb3RHX0ohj6
duMN/HlbX/vCDDvl0ge65Viuc3nYchlH1lfAb/ACnyX4xbSNTzdYHf93Nf1DzPFa
DypWYQ2LDdrCw3ZaTq4d4bRwWU7IR+SGoQlJq6i78Ma0e05GsugDY3hd8TGEiCQf
bGiMSER0GRDsFUrz25aK3+cDhcDdP6SBm2NUINpAcpLJicBhuLuV9qVMcHq1tuod
eJX0qLxRfo9BCJd6bPQj0uPCfp5dXw817fTbhs8xaZEpTT9qqEyeje0ktKes/2l8
V2wbWaUi0nZRyTZzjMz+sxv/YMVCxQx/Acc/j05bDiyYeDIECKxWEtnvNoIBnGhP
l49wk2pNquxXj6AiFmZ6wVcIfk3Y9T2dvy0ZCln19Cg2oJ/toUfEc1qBnLHZG7co
Pbm1qcS9c+vZLxfH63XEzmJhLTPi1LOxGHJ2gVkWP9eLoajSjRAo9tlYlaocrHox
ApmOCCitivDIQn7NwEN/GMedST3PvId+qvkykl/24aL96w6pv+O54rtVha7p9S/0
ldczKSKftS5XbNuIpr9cEALoq9eMEp4wzPnuAcA0X8MdAhES7Is08vU75+5DleDw
3sZnBobMNtBHtvWmpHya8oyRv9TfoC3iXRPm+A/eQgQMzchqtnMSRP/muYWCBwnF
eN1sYdMUhXFtbZYn06enH3H4rxFdJP0n0eqDZI0wrzRzjpr+3qwu8B60/ueQARDy
spQ9T6mRcC14Jkym3KYWE9jJCBi3hpyobQKKCJ186ntD2NkDpJYAA1cV+hBhfZa5
3jMrQC6/ogKqy4Ndn/UIklG7u3agQ32YNYWAAmBuOs8lhAMrkRo24vxCZ2UKsite
sLWCQ1rtYt6UW9x6SCSwekE1hOb+y72ge2xlIhifTbgWoHvP0a3b9cemaw/uY7Q6
XgaUN1MgC6IFtf0MtdPynECK+Z8anN2dDfsc5qZaO/Ne9CvQm+Gr/RweIgLJ9Pra
eAXCuEu7WNA7ZPAQ6yMF/KhJqtM+Nm0+N//Mlq9lXxJrB1z8a3Qxzpyiih2FsAou
j4GQfZV4dA0rakDg2I0rhzbUeV4ntU/bBG4Buzm1aNSdS2rm4/t9ehz6SgiH+NaY
YgTOY1RVtoH1wDMqF3KSVWxvWCrKE28AQOlIy6srNrNUdbkvspcbaEdQ66PaXrj8
HOUl50adp9YYLm4FQLwJ0K2NvRDX4rtoUbdxLe1VwyraLytG/WjYf7Wu1tVYH5av
mBMx1CtS67pz0bE7SY8BYqjd23trDv8hVKMj/NCe9Cm/cHeJSmRc+9g4fCcu/ZHQ
754e5CeiWKc07d3M/FvZXQujodV6rC8QCMLjrENo/CX7YAHAwcp9bpJvmoT+Ifsx
/b5INmhpJZ8EE9umoJKjlavNqFpUXsXGwr8LFdEH9S2FeaU/iDMGiE8h4FeeP5LK
JkUSm7hTyGlHWT6LxKpjhW/6JZbNvtwoV9VxMxfn1XxYv4s3aEslx/PlsSwOd0HG
6yRQhxUXH3Ll85DJx5kVjrCfbMybU1BHW0yq9EYgT+XcAOt8LFIzmrzNmWAjLZiD
JzyQMDu7uQ3AIzViwZ39N/OTGRYkgCJ6fr6SNADaP4IJGPBObVY8qUYMYY6sOaER
27NpzHznn8OH7zncUltQwg1CbBDL+lQ10HU5qGQHmMNY++YLdNYFOVMtppncDjdg
fU7oNxyodJIkRR6tS3Kz1ObLZyCNQcfVMhEwng2LeLWsLeouToopiNSycTAtHYn5
+MsCBZMTCss3xb81W4kBLlBDKzv5w/WLkr/ySeq0XNiHgkA3WP3WetYuwlywdVqD
Ek/PuW8DjDnd+3g84bgu62YF9M/dlZw1jqcJHJT2Sy08jUW0dJhVwZVNS6x6QbTu
V2/GHCxiYjuPrYzad748bWZgwvkIpl/I/tr9hVZgdNfo9PqXViAOBHCs0UNQmlZR
f52pjL7VhRLHsfOgorKThNb8R1P1ZBicJ3HXCKr5Vp0P9KqKns/hUyxrgcdoZRIY
K955nIlOkPXwWHpX4zBVkpARtlIzXs0eZoUBz26tn2V+TF5Q89SZqS649ts2C2h+
ZbjOEh2aMwawR36KEdtekPBenkj9Zka3hacBGlr13sElmJrmUmJFNC9oGysFzdHD
tVHv1Y0mNDoe4rDcBJpJ2n+xG4abAlP73Z1F0ijmS8KVJ7M/bNF3e3qFJTykO79I
8B1mkYL719HEDVkDAnvvLbw8EN6PtoRViqvc4enZNRN60ZzXxU+hED2YgvLH7b30
kQAiwW306l2IDeNAOu2GqzlxdYf++2s+6QMsQaXrNKQBG0g/3ox01Er04DDIPkPR
IKz3EmN8hQCXpi3oupS1r4CnUVMTOjEyP9HEWhTKHzFNb1I8dzTR1ESDe+sVBB7Q
XE6LBJc/b6RFoO9oYJdPPmmtZRwF0ra5ZmLpdmcWQowyBb+hyNDFju9oQlobostu
8GuOxfu0slqSck3Jc45GOgYWzwMh30y1U/9J4zP3FbwvAdYJ7UujMcY26hUSGVRy
yhwv4ZC14aHUKTgv9N0xgQ0JuXadOQ/zuvJnYG1x8XE+Hb3zt5XWWq+h2VZUgpgI
/pwlWPA76k7S2rOek6BQK3TpoWB9PE63hvRJVEHZoTNC29XMJYqjd1z5RFT3vxjv
mKXV1F83zOoDFT3WgorsQj0lJXER3/LlI0w6IdrUVlCLKnPN52x4pMXx8TjS7+yf
vsNPHg6tosOFbVVqAIPKt+9azUQ+7RNbBs0TESo7XiyaRv0XYjdGkdThZeGFWgpk
RfDdz5i+zVkg/tHUGV3LjM5duAS0LkXMyoaPxlGOpud2xM6TiZZ/HNNFsvrHt+QZ
erXEUdKuKM61aPxYePYtRscOd6lN0QGMHRpFvy4U+ts6vEec8h4E2jfTa/5v7C5L
FVLPIFjICDhRuEURcFbviKyH7YaAqggx9CfyFKxg2ox7AtqK0iw2IFEocj0ZENBC
j0e/tglSp1olsY9EUQLr4HzF1bxowC9c0NHDR5DyRYZMMKXGf2aD/R6UJbPh7VWb
fdGtAMyRuv/Cb1BqCyy4kLDOQDioTl81Rj45rtrt4rofNvSYbAGKQ/RgzgSDXUd1
u9m526tX5bNAk0h6hxqArlsmMsCRNyzSKbp2i0KF1c23PyZIwjqhKkYPcwoN+RQ+
Pl5dgZpVOnafEBIWWCWOgH6VTKmuCNk3XwyptcZQB5orptIDCBbEYTRNE48SkAu2
mmm+k0qbYpBM61Yxhcl3+c60eM8zqbcObpBAUio9jEK5xkf21ijqhi6dQybnFKEr
sARQXlhUjczkUIScQTL8q3Ynm4OB2O8ir+XDQp550sTdQFzhos5TLsoE0qthwrqO
pupENnw6SSOu3j0bzyiqxtix48HpfuQmvcMEpTJ0pT44qL1sDTBm4WomuOjPfYeL
z9Jbi25mxxmRsS8ySLXv8Z3NPwfavs3CFJfa4LN/iKh5aE+tROZxNzm+ajwW/SR2
RxBdPii/6st8uK1oYkDd5/ghtZXGGUsVrxTDon3pe4i63wy7iMo9jykOOEjBn1xb
rnDtxsTWiR1C8M96DPoNysY3p/zmoRpKIy4vou1ypfpB8MSaGp91uBX96tYi337Z
22JONvmpn3O2wBHP/WLfFJxlKH+DHbbRipRV7pT3Wohtk7OSNv7QAkj/qmO+T18J
Qjm1tbX6DVKb/w25EN+Y9k96oK2fdW4SsY36JYlEGXgdGU/IMxjwOs4rX2MufwoQ
GMCgmlOQLo3lKOE0YNe9L4onbK0evmCT6bbjocjdyvn/b87UFEsibw6RNCp3xHVL
rOP+u1tGcVpDkbZp9+zczZKBcRvObb2rTzKWi4SicewQM0sBepdpt1Tf3O1V63yr
b3+Swe4lCXv4Ew4/sdwxeajNHJHxozHSNy3b2rcdXyZLPBN1PskxrZCHgoUC29RO
ituSOS/zZ+2nYBOUmPXSBav98nm0dy86POLTihWYVtjiEH4U6qq3XQ4PUJE1o9Ct
I0nv6DMEcA2Sa1BgS/mVky3/9C8wucQ6iZT60/jNMZpUD6hb3qNQwx1oAm8V+9Di
5QVtFwZFECxmhvOuFwH8/CyAC36N2+nxMTBSUfKWIFU3jTyGHhm3tWHO/1tmRAOQ
TRTZ+yrqPLhCSJ6VO3R0WqpgwfrzcgV5FOFohC+AeEpD02/KjBARn4BKULPGAFQo
hsC2CkPZMTjHowGRUxl7BcPLvCUdt30X/AnjO88WwRuNIbgAA4tY7/V0ymM/nPUX
bqHpmyGswUbIhWswIsVwiAjj72T+veTVPyOxOhVeaYwsLNZaOa4fxC5crX7lfJwC
tOlrNNkQAVQLUQaHOQ/2RjTMl7xfErlPG6V9pVCbesghdq+jKyWoWVTNtLhBRQG7
XFvnr58lZuF9muswPvKgHh//709SnXCa25MmmJ1PSRzppzfqePaTWEJZVKHBcMCu
UfW3JEMdwKVHGYXRxAoICzfkM16a91gjh6iI+6BAPl/C2UTheCEtd0Nlc8wknF8u
BV/ki6589oT01GqmdPfs6J6Twol2lA9wJwfPtpSHGC4O0Fu5fabGaaogD5xnlnUs
pLgj/NtmvvvQJHc+ND7TnNuPBiQbgTxF/43sfDsfcVHiEdxmsVa24HasfGr+w+WT
Blm2Xmwxq5OSHizVVkVIJl1NlHJkocHf9hYfkKApxySgseU0KB9TnpSo3Ay0T2qb
JNSt+592lQbjlQFuErvk4bVoFcZFD2N5G5xYnQTpyAQrnw4PHzdi4lFU8RJ5Jaum
yVUg0IyWN6iBsxLWb2xLeljvzbWmMPNzdMXQCl1DyLqAOQFPawOCG+8upivy6JIB
BhmNz+2SknXDRptcyn8wBKapVq8UZXi5cLXN1d8i8SfSZhSV+A+u3jT9V+iGHXJJ
1n3G+WufGROqdIJNwDQIC9ywEF1DMTzfsYZhznQX4BkeO7RjThW9+qtfIgF2gtW/
VqMs7IssBcDa55Z9PTWKRuSElodT5Muv8axwv7KdvNL0bsXVca4bOItcddrRSnRN
VlCQqA40ty6dsOPUFhzbTC+8SiXIaNdQ15m/FEkPv3jXjbamKzt/pcvKmFQ6dHr1
L37+oV3PR+g2Cio2GcZ8EwWbrCzZVDbbgWthCmzmtV3hHd0xHpxCxUmLS+OaEbbx
19AuyWsRQ2m0eKCYlrM2LbP6gCkUOaJCPL7zzHEghbGIufSIn7v9WfahIGgJH9/I
FyJ8iTByYX03ttlLUShN8vkicPwrq05VMnY2x7c5+dvjFIQesmTbn8ff5/HP3VRv
Iyig/6PEG4cDXSu8hBU9Y59LloAHo4zrW+MzSuy9HrR3AWwvHur7WR3n5OMh/jjC
UFOXCP1nqqMz1p5Q3NLaUpo+8yMKHrfC14xkPE1MNH3gid19kMITGvppH6mkIm9d
Vs84pYBTf1Sa5d1RvJajxLzKjUXW9Dup6l3aFfSMYM119BYBCtlx2IVjn/opxeBP
/7xUkFmK0GkqkffEc5y4ZdiUV7Pwjsi2G4Tn131gn/1VuCf+6IXNrjryTuB+mdUG
oN7BPOOHdSntoLI0vosp/UcRXbpZrwR6DcqbAQvIGvPPkFFZh6PkRO6i+WVjJQFz
gfxbtpWJ2/9xPzi0OJbFHx7STETRaYKvHz2AWlhJaPbN2vEdzJyfnl8LWKRymmsW
1DbnAP5wWBlHeWUFGkDpjBRYuBVbME4BxhB0ALimvpC4LqqxwrotV5HWZhgQNtwz
5ErOn0G4M3fZueEr0XzkCnpRBkWhRYMo4EK/emkSvm2S1r9dVC/xdbkaYc1yUvU9
PBJVbhdAE1E7YvGpUGhwXI+BaCsZ0/h3uF+Rf6TZdAGUIBn11UaKtT8w3dy9xJKa
CPdSOYiylTwhjwYCjL2NesI1Tc21qRvGveYBclr/ZkVDlBkUArRVrxkjeebqJzwv
Rwca975AM04pa9eRdIHJZLP4g5l1+cB0oabGOqquRPQ4U+oqxYtuMVGtDHdkULsZ
dA5FO5AgPdYtFGOKgOCIvIY2QAxkK0Ny6VGkv8cJJeWvRMFBsvMI8q+4mDsxdN2/
mHVDuqUCNuWemD6VO1AbA05+50s/61H0yoPuE4v+k9agIyT0Ba3FyvKmiqeHdflM
l9CsF2E4F1EZnnmyV7DFVDhqpSO99OsuRRuHKPV/2YEMAm9zO+MIVIxdV//imV1X
gANbx1/L0z2ZVet88I8uvHb94mCqjEM69KW0f5ZUo75S1pJwVio4rKWRnElP8dCL
IfZIiYIgkqsasRilNDuCiDQC7wOuBXFSLnjtkjpCwiZT2EZZt6w6RJaIS5f0VjQ5
5bIQz3hjo5PNI+D+ykkvPhHusgq2Q7pe1Vkxqw+iAR/ky34LEb+8oHXyw605TTv9
SIjn32wiWqu6srD8fCXE47zTC2DK0hvYanq5Ucp8xRJrS1vQ0zSNc/DrgsLztTLd
HjzYwl4ZgXryGr6wPY9GmjrMtTgsu51Mkldr7pTcIAW3qPM/KlBqHK2DVfEZqdjo
O6mK5SkaEjtPSVkEI7IAdQMJ+6x3nMC9sFzY6zFr6xcDWlErq1HrWJhNOZBGAltP
+9n8zuVVIPT4AJqZBdk0kc9fxargAUC26wAWooHwUQ+58lb0C4vEkGaA0ZCHsdlO
ah/0RIoh025wFXyvEHtgYCRKv9JBFNyAM2jdwazK7LE7wQUciLYfbsesYXbXOwZO
d/G8RxR5MhoVb7xR5sva5RCqssitGfWUpTJW9LKUjVZflzxOG+/EG5YWoIloRw91
8ATK7vmnwK6Jdf4wHvsYKPRVGiL+R9rL1NkllD37nh2XbsyUad5pH5dVwi28cfl4
x1dnVpOijYFvxIywsza7G74YvDsCIaDkjKQ4yQyHAJzf10iRcchCQ93jHkS6Weib
fH6oNUPDEJ4mJdkbgELSP1rDQWWnw95i62MiiMfBdr9irzn4+YyWIGSWTFJ81Tqh
G3dllSeLvxYpJr5NS63XpbUqfKk3GYs4bUpR1vSSNru8DM2Yn/XULHLALOPSn5Bc
3jCxSmhGu5/vmPf08iKtus8o2qTRlVTVnIwByq6sElp7uJKu+UWgDm2y09UDUgRD
0lej4wLpqOgyBn4z58OJw8Yc/nfZd50h3J6Tu+H9RlrtsmTGca7ew1h71LimYemx
NrwcJIhLBwCZ56wiZQOXc6inlpQRg+u5OLMLUfRDlqTCQlHzJFtQm9iegyLu354F
Gecc4RYErs7roJbVRiku0om0Fk+VO2Ei2whpx2X7vIdryJLceH1DMsnOpIFgmZYE
SmXs4nuxLnzm1aqUcixbxxCU5j2q9i9noP+B5tDcdnjx96iw3r+HxpN+lxKe4E4X
OrHPDm0aUjc9nWUus6PXrc++kWMVYQ+b3fmI6fFUT1E/EDdffjMNhVynIzFx1Xc4
CJlpAyc8TIDpPsmkNpEHAIGsarFjMt1vCMAALBWafTIAsb3wznyS527C6swEvkj5
UmG4Qlhf119OxuEGaE92+Q+JrqbRaHR4/0/qxppizOB8dwXlVFaU6N2kK9mU1FqT
7tzmBbc/3eME25IdeKpwdcPw4OXE8hR5DJyj7LjvWsu4hgXM8JHHx6uKWPG2I+CH
wak9K4wO7IjRLdmI34qWYh3KccSbjyzCigfJi7lXMEPcYwuGSanm1wBIRTO8unSd
Ftx2e9Ins/fddAR1FIkIPeZjdc8eMqAvKJPMJBeYvZLicbNCkOHMzDKEcq4GeCdg
fdbrWa8WcFDLBR7NNSk/ARPSLyQN2FwkYqw9+Rr0+jDaW/+Jq8Piq7ZzrHZteoWK
Ua+Xuvf6nkw80uGASlrl9CmykMOJqGnpB9tNAbcx6QndWCekUFw3xz7S0sQ0+qk+
PDiwBPJTdBKAuu430KR3i0M6kkuHtt9QCW4EHfDuaeaBVjmxuLh0eJEmmuAuv77M
eUT58Nw/dBh41etd1xbxB00VBO236dT42elAy4Xt92qgLdGueNLw2DBpTQrAO1QR
bQAQjauGdCEvYQjq3t557nA99OawkNlVvYYKR3ZiyDsiujEXhY46jKDQYcgDS9eK
WnDr3izkKpNYI1+zTlySJdgX719eHJdTgu8Ij0sBfF8Ov4tC60yCmK6E2E4V8/Pm
DX3wb0W9fAapRbewA7ssInWYcge0dgBiFIikoDYQQAmCvzP4j0KC0xIkw3epNn8F
X3InjICSEEI8I8r5HwNjxzoFeoo5eg5G+6yg+YnvkujEnDZSN7a6ohZoZkFL1Efe
VU41Rd1TjZ+L3uUZll1UmDZ+kHQo2lu0kRvJvPq7A0bzlcEIh+xKm4iLaQkAeggt
uTQOv+Dfpkd5ac0heESfBpCYsayK9YqPzYFaFgaLqPqllNsyQTS4KDzXKvu9+9PC
pqIY0vVmLM7mrnhD/Kvt/0GmMR9IPKv1ivhzzOmKVYNtLKreF2tdzvN7V6dBl4i/
jhVIhFv0vbwv5ocnmKly2X/SUYwz6lBPm6xdNsSF9QABuBgdpIxYjHpDstgAUnTR
FdZQ9wkAQkbLy2keR2icUKJZqWzXH/XQxgWFGyFxNX8nomz4Jdf2NMNyWVJnbURT
IWxe+FmoswR666U4/rGrsNn5djbfHEi1T0/QLQ2rBBP2S1b2nmFHg5y6Jue1FaQr
zeFFNlJB6PU4th7C3JATPjo25tWo4aZjuJAzoZ6iiMz1X4qZfr56Zp3iyJn9Ftgz
sPIavVG5b+hUA5xPK9cLoFKbSTuL8XUu9/z4/GlkiP5uSqis1h7sXiH/WmEPcc7G
EtZeeeGudwP34D4aeRyfwdxnCkI/oOKaTsMReCeUOtZ3reqRQtnTaUD7stwp1Jvf
gwy399NSnSXBODDXwWXM8XAj9fEve6zgqTP1MltaokB23I7k2q61Y9OrEy5NbsFL
2tfGNWk/l84nBVQa1FS6vUveehQNW2FGu7Cia2WNTnwSBgwvThuivqsmjmfnixes
VhVhU0KkZcsvZOg7yuM7gPrbTslp7nNWm0JW5XFdLBl/mmqyvet9L3Od1eKsET7G
B/Yjeugb0SPjWd8pl8hD0S956JpliD0XJGSnW8fvVPg4p3SABtNGMmBcernSo8dV
CDk4ywEpHj8CAYhLeT+NXYRY8xnsdCzg+AZ13vd8/DxsHJrsvS6CqzRdPjpNtDNv
Iy6zxTiiPA52PXR/7hvhxUstZ1FMb312oqA9zHXUhpFAO8tS1aEDXDXxkqOeXH+E
CYkI4arc3IZdI8PBOMI1th3XGMmzu6IOKjs1lJD9fASa9XHehOBij5RKKjGSO8ZB
Bkp/nWAIhFjprrS6LSUBfsP3tnm664Xwc/n39Y3vYQbQoV2+rozm4o2IWzmUCEvK
IYfw8EP6ku/LDtZLRXm+4zeXVum6TKfsBOOycSJB2pUJxSRwQyk86aDE0r/A7cax
D/Yu07MI/D4BiFefWOtU62kfw4qz1yHRYa/jKWq8LieWsFVIcJvedrMltaqf5EeF
A0Tw79X4gx4lDYLBWO9wwf1LMFdER5GKXW2ht3V3Q15jyrS3xHODnYogntxPAUPd
4+hJm/dsgZLoDIhXIq84KyppaDyjZVk03r9iGuaitIFrX3d1NqWv7uKtqwwWmdOq
DazNLw3KQ09Yg5wYnmAC/XKJa44ZOHbt+T5UFaSSHlVYW6Tb/jloFSBk653xKzjP
WJ3JHnoXpNIHNQzuhWcfSMrOJ2XgD26ypzoQ/HV8LR8cGZ+76u6UJcB4Q6XhWs/8
sGH9hafZez7SIQe/dqspPUPZUnJzqwzNVQVvHzlzkDV6Ur+H9xlasLY01uVknJf1
keS6FSe/RsQlXKYg2TYYr4PbKmsaITLAmSXpLZF4wgrJsMEfAd0tr7b/S+4TqDqu
K1oTlbq1SmbixeorUNrvGwvm9fLaNVgeURJNj6RbzPEfN0c1n4nAkirweSK2Zt3Q
OwGhBKXlzVyn19mWig95WJob9tINWAqav4c9BvEztHE/2trGei/KK+uq4Mh6yVTH
4qYHLH93ICqKe+xZLPKhbGWYOXMZ3N6XBKbPSH2cu9jNNT+VXzfXX/AnQVwdPs/7
53rZG67Rz7fHUyCnoojlQgadQFRJ2o6WB7/Q6qLODYk3kBFpSKcLm51Dgu4GVFFr
jd5/dk8/w6ieCS+gmRj4qwdDeY9XLCHDjMYrLnTvldCCMq3MeLv9p/2ZlDd1iMaz
0rjCGEXwaRgIh3Om8PV0aOOQNkJLppNiMvuzlCqVvyyTdofYB5lL2lFGTtwh8lDd
UYpIcrQeYKLRUgRzH83v2DHrrF+U0RMDqfDrqNuCH0ePPGXRg9MlnTsgrZtxN72+
mwNA7tsv8upXNBm90O8cZ69iIZm/lxYWEG01cRaFjWtM+q5/MARwIKYfLc/BNsAl
25N5101XvZRxcN7C8fO68p69qyuYEpXNPIuCm/XHXfdHYKBvqBjuGvYZqs5x0hPe
4GZy1dyCyVyqFZwnziRvOjZIK/I6DuEt8969HpflXjGm792m8jd0yQqyCXfGiyxm
rA0X9stotDeA9iCt+XewWLa4iTqhiHDEOmLWY/iRV200cDefxPu8GQ8rDw9vr4il
cz1KmJLa6a4hAKMVX9lms6e+MGm1HVxTOAadhi0dFCKJL/6Vnk1tK+0As333esoK
v+hlJY8PHj1F7YyrbY+hX9rhGhXQvRXSyiD+MzUJGNsL9oPnJjfkfF26aGW2mv4C
GktxvIIFKDiCPDYpHbQISZUpI7CPJaJsmarxQuDYT8cxn8bVmxz22XtA90Vl39TB
yzFsE2j7qrJxL33RKZSm1oFUIkOZHDspDmn72YIO2SAPOlPLzR4fkPCrVGUQlBS6
o3Uvmvl0+9DL2yEpG1DqmvD+WM7eXBSacDRPOTQJpc6wR4A15Gr6+m89qHSpryPt
Bv96n8u5018qFXA9lFTLpHWUAEAv0Ziq3PxJVvriTBbU63Fx2yK64A9K+40QMmfr
WB9u/esQr+ePzo08blhMCDox6zXu8PTPAw1dLCte2qVFMjhZDzmgYy7g9NzBfJ5l
aMkN6Jt6YHHU5jglcQaD20AB9ug7NZ5JsD/Shz/HoYlPZ3kNX9NmsV1JxllSgO/I
SONvu2khkuOY4XsgqfJArovvtHDUb2aXLjqGbztJlUqOi+4CBN1UDyQf33IK7uAe
TCB6JlBsBJYuv7FpsQjouKoWJCi2bVYGr7xB2ubODZtRYA/dzheNpgKcaKwIH2W7
1jb+3A18B2ly2PwZ9z0GjieT72yM8Ko87CDdGAM/lFYN+V/Jhq74GZERZc87Hadz
pOBTTTFL7aR3lk8JYFXD8BSm2c5+8C+zywrO/ov31BtFjJbW0stBN5qYXdEl1Nfu
427o8FI0Ya/X9y1yoOXORz46Dacq6KNxniHpzHii43Qg+m+cWoIvvLS34tNFotlX
tCFYXavSI7hWxxdvv7+awiTDREIonq22iJld2OLhLYEYa918EHV5efPIvxjXUmee
DCpAcxegZFNE45+u4ibXCGRiQcGe2YqE5vbDT01pqJ3+pI9xteiwG0/1wFCy8kyp
/PLecuFLGAmhS1KVerEYVoTA+61Izy7Yf7lT9N+Qdg7S6JCBbCvg+uieNEoAFtuj
qgDmXpRYGdRsgUu26aoaUPNaIUtufnKJD4yWn0LH66w9V0171wkavxoxKOlqBhIE
Gacv0DnFtludj/UHwmW6el5lbMtmdu8c08OLmISQejZgU4pFoX6imQPzZvMRKEta
/1XiF4n5hdkDxf0zqQyDq477JE+deuXEE68HWZlW/jYLuapQkBtgbIFmbb/nXikT
rhX8NEjY1d/bO2Tw2LBzl4xmwjyd+ayqGk1dMW3c63BGKwwRmYAQNEJRCzmeAoqC
LXw71hHaF/rz9RJKRad7S8xq6L3EGembUHsaLxcLZgwcqSfjAwWTN3KmdmDTIQOC
rskfl/jljz+l5E4TytroVdX47n1UtpBwAuIU+xTqsC8XxiwteR7JoyYAYTu++zFE
k1O+mJKgaodcZkjeBoGyZiCncpaxUTQXWYboRk9TJMhBDlSGQKH2YXbPVjzCvExQ
YzhRBl2n1dnPdYZMK2hngvtXo8810Q9AFiWWRK4uhXuiOc5S5XsKGN7qZHanFe03
HKH9g1pxnhytFziL1ZHUrLNS2ibevRO+q3eTb0rUI9Tm4LZwXiwVSBzgJYaGWHGW
kkhzy0YSQ/HhkHZVUgMznLFse7qiaS4p0Flmp+etd9s1bCyPJtX9VlUzVscn4GX9
q1um0ZTx+d20cY9dDXBZ2l8f9NlditWeQkp37rL3Ku+M4+t2X6q1hLlRVrogqjxE
pufRIPD4p1cxAFRLfj52Y3JIGGBrXkbFeH1uEU/SYc+r+KEmUE2V8FHtUxFwI0Tb
b0OS9mcB0BC2ZueFbj5vCpUwUJi8DNQc4MoGxftNCxUAtlU6PZ5USMeGplNNDuyt
NUUvgRI0+eui/cMCS67PU+QI73YfJCQx267U9dDevW9nzq9midhfY8NMwmHzDZtE
87FEWrwwHCmV0I+zsxrHb8v5ncMNgcdUjrSLqMyS7n2ZNbXHzlrG5VyQWkSNpDK6
JjsQFetY+yqhSZTiBcWi/xP4/rLGLKY2CE6V/GJmwe2neSdz1mvcOEuA00AdgJRH
+FBVntvEvOMKywDELlvKPRVt0WaR65Ib8vYE4GaCZ+bd/xArWv57EnHsp3QX21Mv
Z90bIVQl/j9tXfoedFJmkfq018JgiBDKdLYl9k78zGAvU7tvw8hbCrS7QJZZKpLg
QPlA3LhMCO9H/zX+9rmmAZjLG+RljNQvrXe2UMBNKm0MuE1uILD+CpTbcKduVlaf
ImioYGptIMubkwKDbwy2WmlWtT/d67K8IwobT2I4SOdEl6fQjq0i7uZxRHqqDAnh
o4uFsdB+v7OVGdkAGECk75WLrPQjNRBgISXRAp0eigwJJYVgcGRmjeUx0ZTvH1AS
XVryyaiAeohEkvsSgoyUkHX6bjqtiGxQNWQuV7RYgaLt96RWS9gtbgJIa6jSR20j
y5tp0em2+VDnwkLpU8yw+CWMRh9aVt6fOXAu99y71C8skBBAbD2InmJW7U0A6FPH
+qM8Mfi5iYr3GcbGiOe/0IANnK8rbGSQCC6o1ijiF+FhDXViapms4AZ1S5pi/NG3
09iFnaRZ1FkhgDTzZK1DNIEgFefp8xiaAxNu70cMyrgQ2UUNKGDdSaCR0ROB8TAt
ULiWA5cuszGByISGtQmctxAJdie96BLUsqTN0XKGK+/2KmGSzaFClIWlq1b1rAU2
PXyTpQsRKSx5chpLPEXqzLjV1gEHlwgXKy5dtQcgioj4bAMtFG24krJpTuMhiUpI
7c6zDAyltuuk64NO60rZPcLvnT2Ir9Ct5Qv2rct1uUSM+JJVwpJ8qXHEVTpCJH0c
pBe7sX7xb7b1uWZcUGSf1Zv656AQKRlSeyCDWR7VBC+SUzRLVdRitLEPY9EAhbxQ
NDW0SywitwrrkKGH1YBFjdBD5/9Yj8XSJi6k57Aveh34Hb9Gvy3w1bhqKIAugOZq
Ph7uWjJAw1svJM4UkPN/yD0Gk5nyEIyvas/ky51nUxBjUsqy8BFlTtUiZvslNHIc
VuIzYjqJ4pgVzg+ceJoyJ5ez+PDKyn7pkDVDvGq8PM/vRAurEFhuzVteUGyxb/rC
JBsHST330ABwjnwqYqCpYmqVK2OQO69gzWHZeDENOhVWP3/KMluIMElzJIB5ikZW
5qMVGSxGMB5lMMYAdFR/jF8W80Rz3+SkXhv1K1lgaliXEJwhED+JcvL7bfDBfUv2
Lj+8s/SW/hJTHAbMtw8UFUCyMNaLrApoFnvNVZvl4lgfNvZq2Bgp2TfZqjTua5q+
yrMbGt3f9TE0+8mKFnLOLk8QvZfe3HD32PGIvANQlQ4R/S+9ksZKyYlndq9dF1qJ
a1FGtU+bzkeyhbovb+Vfw0cMO6NFaEy90zGR73Et8aVDE4bzhKNBG31Z1Cb7mWhj
AttJHrr79lRdrSsU3PjQKTXRAnOksvqs77cA1D1EgF/T9ZXXDru/wZUtOjuiURov
iO/Uhc5TUv+gf5ZCAGyY7STHO/cfbxqN/4LGaBxGGX6WZsyO+G2EWho5XSN70tGe
BneHDfFqlZynAc1STWnem9yRn4zmMMKInNa8nOG2a3e4zOTKqwmG7KS647dUzzQR
fXFTi81Hfd2ZV/scN85XFbSZSD3g/FOmO+4R1EkL+Ly/N10b661UNHw40KVeFXHP
X8+UqNvkptzrZuLOKXeQ2sMy3reoDoBUkVchBKKkEDDw5zCkwxx+h/+TzOP3HH+6
CT4UVH9i3YMma9EWO00s3fC10yowOh1j3pFaufxvcZdCAdnUrYcvFdPbySX3KnXc
Ce6LaXumIhr8Nqy23RV++mo9C7uyxu1r+whMda9CKTE6cIDJqTRJeGNFP35xaWI+
Wn3Pb0d6u0nd8GINffIZxalivTLjwCPD/WeHwLNcfyrhMmhvZ4LZDnLCekS6y/+a
sVTdRejlfr++tXk09jSEWL513j+GZxsGSqvec7MJsW0HPhZvwXnZgtzk8dhMymq3
0K/t+HcLHyO6kN10iRytuE7HPywHGOYfKPj/USPbc2JfJfSuxMiISHcJTr7pVNMz
JOute7tKHSMHGd3XA2ZMGtBfD3THQpLqtXvIbDpRsuh5tjBVcPAuzERWClq07Yjw
mQ0YbG9fi7Vv9RmrZj5fV+RWQ65EL6sN19g3KzJ6+ATkUZtBJSkai/d7O1L5rWbY
GPk4V6XgzoCVrAVZAaO9/Qz0GJseb/C1u1rSLHwbKABDeWwwu4QsnAnTAKWKl3pH
9RVA7CpGkGXUtQRpOj5Eu0Q8xkbh9QW1skrMcs0vzYBOO9TtUggURWEdvic7i3p3
rLWhZZrDR4LtlHNpOQdji9WmgSCJi9D8HcZXq6EYxJwt0ht9oawgqhC1rX4uwO9k
dpUZfJ/3D7KHOP2Tavr30VKPU3K1I5ocdvkrOcvg9HMMqEy5DxWdXdfitEY/cxVg
atrSTiYP6xEflYkfyfMf2es+yMtmjoM5sKfBrYGbPhNXCYJ3rr8m1+NjBq1E/HGU
ND45J2QRUPWynNABENxvqCB7x7Aa5seiscJ+iS9VNTzN7/v7mwl0nweE9JJ8znMe
H5PM+YGREQ3DzPK9tzmySoESGcUggm9vK9hDdLkWiPeaNzoaqmPWUI5YMu/TGako
GpX5KrcGTdpKXaaTd6tSNUHGtz+aoRB2nZdTY6XY+qlmta8dXXDhSlO7D7KG4x3y
9Nq7Pyzq/uMZW4gI/QTOtm3LDQH50KhhSMLORyJBcixJB/qMAOyDMnccqga1swil
KXua/sRrX7LqFBtt3tuZ+KC+D3Q0Hr3/t5vWEXJxNjBdTfogry36RSEwJ37duE9a
zSs9jqFMJQtWj507+Uxg3mD8cG4DCH4rP9qiN5ckpzDfc79FzYb2PPuPgyeIAzbv
wsDwfk6NQGY0/YEQCQO9gJdfZ6dLi1SPpgb+QlVeodFYaAbKOgvLpGUi7eI69ucv
2LKnKoJjFAIfy+dlFuzICkrdGv6s0nC+7lwz/XIYOv+7r6z79RuRMdOoXnF/S4VH
Bw1AU7fxSm44msmIkJ13k16gIO0D75gf79IpFIwNO/NfJv8TRA51NPHLAEsY92Le
S32hFzyhZ+FE9PFPSprKjqDi6MADnwk7jCifIfK8Du4BjYCnYh7fcAcCkdwujGx0
oKGAX/M3W61gd+wr9/ubrKLhsf7+PcbK1isTR8wGfrINUVbsowbxr0RIv68H8pZA
mxwFw41nDEANGv3oONH31N7iP46QDAA4R4e345Kuifot1QdntRkV8Zb7tSaxkfhh
ATlkXNe4amA0dPnB6IQX8BTUxAuoZKiLOkanUBCkw2CDlTxyVw/Q3aP2j7Xzciov
TByw6nFUd8iZJjh/k4OaaMXbWWzlKlcZZao0tSx/muL8KlqsVRIe/Chf6rTF6Qtc
h9Rto835yip2GHHaIAhD2pEG+nYezsTGTFFJwgWGXwByFY0wUtdPxve3ju4tpsv/
jB/oTbI3Q4HEEiZxd/pg0yxomphCP1HO0H5z6tPS/2KsoA/7Q0WPjyH2uCqyF0Q4
DPJIntpks6s+gUuXWelHnw7x/N8/4obTaTvWws9oXR0mTWXr9cT1FiaZvZhVRESF
xUrHRU7I12THc/tnl/fEv43ZCb1tmeKWFUUn1pX5bpq2Ngyjwq4ZrZoYQ+NZGqD6
CBvbiEoPlue/w9KbUYu6FNKVgvEi+ZZqRfJDLaYFp59251ZpfUMa55XOmcvojksB
PBa3QeCTJ6p0cSfmQ2i4yjP1Oob8ONUHoK/0iCrZYXOJ04trhlCeBgAtBQjOzAhW
F3Y3yy0r1edkVXKPqp1X+Z4SdFOxbaarSj7TYuQUDqBsZA1RBH16TDDjdY6m3Vw/
poLj9eys3mLwL+LDHSFcusQvHqs8qIzSy9EApQ512t8AAKSfwN6+h/QsQskHuLzx
rJdtKgnVp9Wbru4mqc+dLDqDe5kkueoehdmfEnrDvEonoFQvxUQZup45Pcp8JZO4
s8OqVeBFaiR83Kv4/MEJNyWcCnMjzWsW6Q6MbsKq7qu6jRhymTLytfCrhlTsy6LZ
QpJYEOK4MlffUxpPOgQQnV4Dih6VxJdd9ISk1a7zKJeV8aG8W0kTvy0YS4pkJ/nC
rgmfhZWcoSck4o3VR24Tl/nNG+rns7AnGY9jHAzmCNUqBx8Wtq2aGzI9nZKXrH2U
zv2aBtqua30YPTLiIUyzoE49dYBpEIdidyi3RkICEyThP8KOeLtJkN7/7RndRwaS
SsUbQfUV4MhIQRXUxMNj4NfeNE8JgXvdsr3X/7PyJe/iL+zUZ51eBc6Iqdif+mv6
nt0VUNiImMsnkrXjSET0AAOwUsh5wEuL4MKl2kJJ0dmb9DDcQboIZ/qToC3OMzTh
h2D0fbjw0LrrdfxJJGZe9eFE3gdwaAPADaaqfBtijU3AgHLRZ/h3duj5dhjSi3sw
iSe1xReZZrOVuZrE+x07gWK7Jm3pqg4Mr3o7ftfkc3MPVIx94VHfJJXGuyEy3Eog
fyc7FNKF3zyuEiJ1EqDF5TxpcHKIzZWHP+soErxeRA7VYmTGqTrpMTTFchAuR7nv
CAbvq5JT/7pTcySyK2Y0bPU7UZ2ch/jp9+8sq7rHPJByevsvENhWWHmagG52Odkl
g6N50YPMbkR8NdktFv1XlbBBV6FqNe56yzq6mWZC752nrMmt6I6uLEo/U0bB3Ieo
Ho7od8u162n7UnofkM3p7K97pHGIv0hykr8zMHyMoygTOjIdkhoLFuYyspkb3zcE
39KSqcFsyD1kG16y687BNLe1+/aa7wjIZcualCBseXGhNsQd140i78DscLj5UHqR
EATrTi/laWDGziCCuqJEyjTzZUEjtzBGFHG2oNksOZCKQHad5PRFlWAxQtYvn2/f
KYeABfO1g1k6aCu8IPz64CHIpvDSq9qQZ+MP/p6Gg52hKNSUxmobQJzLz9trZfyS
RAURcJL9ewIdMfE2VcShQRotPmuLMWrSJI7abRnl6VGBSYZvdeilySaPiqNCD+dK
ACHjAltLF6pJn4w71Y0EozGEQf2xHleYpEoZFfuk2FPtLnHqk4fuo+RQT0mom9c+
5fYRfHgGEAJJ7hd/mFvH25fv4rnooP+whtwnGwTJJVUql0zVm9Sbkb9v0XNTVodY
lJ63QlNq7QcjAuogq9rnNxbIdD/CsHmahkgrplxK1wh5iEt4ED73PVrbe7Jodq5j
e2O+gPrinIUvgBiqqYIV3GxlwmKDQKtA5b/YyZfZtQGMoBxJe7YkF9w5y8JcW92W
EQoZLiYypkodjLqk/H0eASyqT9hgjpEKA3rnTKb4Zn1wA/acxGgnmv45Y5y2hHUV
S/8UrVADdfePhUzXQ71mXkONzNky8Ah27ylpQWdZKwp9tIFPBivDmc8Gu8APkivr
iud+uy3pmK8K5K9uy7oy6EVUwtRs5apGEGX0Es8DBe09Xq4tE+8P25dWHRTHAn1R
GaxuSMlseT2qJFtt7+IuOZnOu9E5esspxxbj0lYCxSB0cfxtq4dHBt6AI9L1KVTF
vF8ht/107IGhEahBoKuacpapaF/g8qydZBYvyMMiGIPmZGGcCTEsv6B/lkML+rfg
hM9jeZkd1lL/FlffpkfgtwNn1ob6dftAFfFQKSTv9BhtqcRYSI5jPW1BVdkHArcu
byc1JUXNAOs5+Y37KUjB+oJAQkXuH1ple1hlKENZrVQeoieEtlzVjW+8MNZWGLXv
t9peiF9UTASrFAQri2HkJgVi4WhSf9h5ztvGJTgMsiEK6Nr9Tfw6NxVNg7mgGboR
bFPFWPkVbHg8H+8rcl7JMwqnNIKseMYNDS0zW0M8NV9UG47z9GuUNH60elSC+OsY
Vdb3TbxytF2p2zEf4bN5k97J/Bvpl0Rwt/1hhBE8KdaMzrJ8nyDVLUizJWETSaY+
nUWC8YD8bpTw1jmqxpORS8iI3BhVGZgyGsR2BcwwlsFpUMciz78BZA9tZgGXoDhs
/mCBi2h4pnUi4PnkHdS4k2B0kvi5v0C0gp9M6itQEp2ijPhivXvzo+l9RVt79knu
U5yMH0XMNXOjL0WKPaNPYwxMmEUvbLfn37myU2THqjwEkxi+Jzc6fiwRDKeEoqdL
s8L6AKKX6hWezQO41kKDRw1CS6hCwos519qNRaN3wC8U2Vlg3JtPryOVBMch7VCo
IpMz586Di7d2A3s9zIeuYKt4J96TlGGYXSBTgYgc4fQIiIGVz9agGqu6lqWs9t2x
mAq0YrKVhdBbAJHugeYjSG7caMGfWcK8aLkyLOY8MH3ImEgu6N5N04y/hxmBUez1
cXc5xxcbGVeZHNRQnZbgDahHvahv9x5W25e4DNg01R/kWttAmnRYOXof1dKzUCAu
aUAgo8w66rm0EQetZFDyBbxRwveokYuF4Ka8KbRaLoC8Cy9eNQxcnmZM3kZT5M8K
qwPj2NIzHjhs8QmhSG/WYMfED+SINj9cPGwgsX/Hk14iT4kwKo3NqehVBDfPiWP5
9kQ/Hmd5Coltxcapfzv8HKncM5UQnQXPpn/SOF/kPnx6UgGJs5OLrgdQwyc+xLwQ
neUoHut9Wbx5TRe3s1qgkhvpd0AYYdu85RmPDq+OW700pVeiTLbMh/Z7/5oLe0c+
RnrCQGFPRxj1Wo1RjA3YSP1lj1KTV121SuwkXwQB2uqKNwSg3AmsK7ZnSNApNMQ9
2fXVVI1v0grl4J2F/NwbJw84rFSXjfp1UggsbQQFMJGOkrcBfFaqthJMIx0G0XAp
9YResna93FH1flQwwKIVwfu3td5jvjN23rKjSONdD4zo+eaFFeAmAfP9AnaTZXbt
54OTqnhddy2ir9kBsMesCUkULcWGR2BdaGy4xIUN2BE2RNOBNOtJjJunr5exbLn/
BDlKhMs+mlamAzN2Fdk3LX15nYO6IH93bQ9yyMiLhqJqLa7STp1ht8Qhl+dogrz+
BNP7UiTlRIMDs9RXXGXzvYJrC3pxidwKs3mM6DGxKwQ9sIMDffUsAMXM4nwal27m
6OLQ0q1yDLV2YhEXxo/GSWMRTWp7C54jyId1qWzOV/5pk0R3zk5K6tWVIFLw0NhH
sxDf6JRZ4njcuEwDLIagh4OeWjGAK+tdlioY3D/z+9meALSvGoTxKOX/C/X635sY
MSwrj0Aa4Gcd0iI8BhcUgAchw6PRCtvOZEsBclaoAhHJzT27RfEIXYtW2J/UmRtM
OJLuf6ZPIZqRnk3kuLlUlEYKp39E9Xhk5wpVzxC7jJEwaSd05YFFWzvVKWKUjLoX
rsPDSKO0hrTCkQ8Wczr2+T+IiWKdcVPB36AW77xd9zWkxxynEjzohMBbX8+Ys4vv
ucfrXFOcY1xuz2jFwfH31boZ7F7fGSi1vQ7WqpeE+jOFLSqfHPfNCGte9XQ9QXA+
+bfyW0bjCVVeOvD4VkIqjf7cAxV3iyxSUDHTw7jAIO1vrXZoUrCxQ8d8kssyrMMN
nzTlOrpbq2y+ZxznWU8MTd76BO1WYxVimVgfIzi/h5uuZb48WVBoMm2sUy46lBeL
njRhk/X7N2kSI6IJzDYPJJB69tA7VOL9xVg0Ke8RHGioMsoYaKFEZNKis7S3TxiF
a1eEpC7crHpdfeH6LpPnIoeq80gG+Rk75pxUiyOmbJhDWtyC6cE3wW9GFLRxanTM
LbhyEqY9l1UdWrS8E3NCMeUhiYXMGwpiJx5NYAsEj4+RXrFLF8eM0MX4X/T4c5f8
qXEr+lYgASQkJCNWbGMMzBDGk5QZ2qAlAuvpJgZjCsH7eKUdLFyBPUwvFbk6D240
MPmUxN+JarGj8cYC8E8McDzack/9U/8u2aAelGRqCptIK9IFp5rpBCx5xaJVDSOm
cqdRTNUiF//gMxtd8PlqEY6iRWs6lPfwvI5asxiu/fn9sBAoOtRZOR7FiHVNGk5L
hjhlfsJxP66RCXwS5GerEdD2BUIg7Ga8jWSHnQ9U+ISUUSEtUUFOnulA3rlC7qcp
JoF5zPql2UV6ZiqpYQjfAkGALM586SHuTjW6RmxrnVxceLlR+UaM/4gmpV77+ZCH
QY+pTuq2InyOkENiOQHDNhB1iT4nTBuBo3FDPf9HDLk00X/X95+mqNhd03vQbPs3
KCzWF9TqYgH8Ipd+QdUHbh/i8vF4DwWXIr6VYZw5JUwBIbDMl1WtYTM705GsovGi
Nl22qoQ3JnLyYfUUymyBIzg7eNyX0pjktVhfDs7N44P2j449Q7V3nOBBOmQt6CNw
MJ40eT0B4XdBQ+b29iXDzH7bxfTmMTiqP8fRS4dFpTZpVORHfMe95n7B5kQ2qFf/
HmWKsEHLArRgAYX/1KFS2l6odIqobl09GHQygEaIfcbrNFojEZrL3IqhMsbUNnbG
Vu+yYjBdwq5jKkZTcVMUo4RqFZLDCGSLTPJ1qGf90wMcbWnPFd/KUk6gelIb2C9q
ng24vSAUnkk/fInr+A5mXETSoxvp+L5yOcPugOwbLcCb/rQ2hrXvsxQNltVmUv5d
2e30VMI6Hd32wY8jO1EM74qJWfL1SwcRftj9zi9F3r8BdyFKcCUxTwPVGR7xhY0m
4jGRwgaKOq+XDBOpDNvLuDe5smN7yZSxQog55bs7k1oLZLKCTWdS/Z2VYzm9IMwE
xOk0tQIVkM7Fc7ieHRBerLb89puaAB7fsRS+ghwswR2WfmVLyCAYgLWjDmO1h2Ro
rEGzt5p+cr8ovscxS7zauPz4/VarZqDwypJ6SFRteqr8RNKvETj9cCOw32lHaqwL
nO+0fbCWECsSN4rqgN0a1CiqmmbgTfH2QcXok65WQ9opX0NG/wEKMkux8AdkrQ/a
ObCS5X19j2bnH+lRGCYeFMa/yatxukDJnrZieL+Ots+JZEXvhXsYZH31MdfTCcCf
qwOtKrWEysjgMNGp8pbXydGoFdbASIbjoifbZJ/9rLyK9w4GYPrpRm/XGPYAV4fA
O2juJa92Pb0UufZhwrrvVGZsongfxqMN6NYq4TxEi476IWQu5zgraHQwmgwgO7GP
dCitv9gyBo4/kzIChN4DidEUni+ODfeTUTu/NjKlZcs2/g5BrI6cBuZQYGVDJ8JI
bxPWz6Yim3VsVblwUEpvljbiAJrk32I8W0G71IunLlzyYzYy8LDY4hvIHTl5Ld0P
gxotryOYYxGA657H4k+j4D7CZSCVaplk3x/zpah6UcYNA96gpEZFzLJTA+Oaf8xF
KncY2Jyo2/SlEPAN2TKdBr1ARohiwQIfWckNNlek2oIEtynBXL3vEUVyo3nEkhVp
1HYpPCsv4qSEuzH75DIWWJ1Quj8edx1s4nHh+qxZCahx4sIfm1Sz5B3A9PvRWm/+
HVftOuI39dtp1xnJH9Ey0jPjQfz4xrsuAQROUhSjN5qPUz3N3MJyRKCdmogRvNbY
mcXWRLIJkIKmdsqvsIkN/XqNEF7I5dhSf4ppqKpYsl3tXqHg8Gtfv2cq97hRjJiv
tflfga5HQfKP5/on6YRedRC9wfcV9b5tOcUmDJPrmPwUJNQFQZToAA2L2e2xr1VH
y9iX+CgGeDvVH7uLTDX7yvb42SlTyWB099fw+JWPUEgzl0eYtfnpDRv4ICLOoCY0
4k66kJfp+re16a7T5wO7kfi0wVULMwnLgmX0w3dr/FRDxwfAA8fBrz044btIkYTp
ql+frE6vg32+5hNs3NXYhZ8CgsCGyh524pXCd0/PnJ3/n2oL02jzaoXZ70CnASDz
ufdwHK4n3TVmRxVNrqX0egWuh9EPqYoiOUMqcpBo2o75ImabLg+c/UemKm0rZpQg
J+u3+pgOpBB4K6vEl1qw59FXHWFb3JHCFpmcKfIUj5lNDAlMS/IbazPIJdpmiFu0
TcqTN6FBsotYGeypkKyy/x82XbtKZ2sNP917qSPSaZ1BfkpRm8878ebbrJga4krs
DhlpVnhVERzNFs4T/wsmiaJfm7MRXbPZKBjMYxecCRYcIWR1Liawp42VG4S20loe
nERmmxYFgdUtlBJbDLeaoRsLNPlSwR2XTi6cOKG6Xv7BnAi4cUOhNsPGxg323Z39
J4BscwJq5ijmqT5cuAodpuFKJZIaYmfknPE9m2ii9p0keZ0/hx+JguQugf9Uncog
i19Nq7nwBANLrPGT6212INWjPUvhCaNMxeu2+gNg8T0+IrmvSKhwosObeBOYbpNj
N6nnyAOQy9E8D/K4UpXX4iZ2dqaM6wf6D4JlcoXuuuU1qMRnamgNsfiCKcJbMSpO
jb8XcVjQTHFXcxlX/nqT7dsC2BVl3RerTKptro/yVhMuFG1k0IMzM2T+RlvdtDH4
d4y0tjocu3zPd/4zabEvFaXsQ3k2QnpvD8e1O8yLjsHA7V0NPdSZAN4MeCbcD9fH
7xn6aHdMEy6oA0liLi1hI0Bx5GHZ6EXyWCVYfF8S6MbWedrmSQ82nCsCYkJYjd0Y
BZb1rrapo6iNs3WGekfKGf/j6GXNEQCP5knLOM1cG73qlO2xIcjyAoeom9giCKqy
Xc1UfmMN1lghRx8/3ZQEXknSYSJQGDgEHUBmLzj7Ecm8FhtqL2xR+uRXPsSFXXl8
oGJLcQ7H1ySznaNzwp4fLZv+rSTw7BbNdcjeBbhw9ANmgfRgTRNpva+wiOUkls6g
p42LDc/zFyn16l7qHwFLLTvEVXUidH77j1GQfDsc6ZPaFCwa14q2o+pY+WyNRX6n
mCD4QRrBrJrw4wgrfHqlnWeD/wyG34jgqN7uUg2NDBP0s0psz0OIu6fGX+eou+7H
9MjVjeQsIB0g+zJlIvO5XHj4LlmC8wOETCdILSZIlN359pU9/bjuVSdOj4gTTXxM
jBdWhJLZQou9a6ZDYnCOVFLXDLYPs+z9ehMM27BGkyItDIWWLp51uzdUTp1tGLJY
uRvKvNyfng0GX0uj7CMKExjlNe++xG82+lmeK86em+RRj8GKoijPYQIdWVjR8oGL
z2ifBF6zadR4twg0qMquVlF5NUirkA5LJLsS0T63PslfctSTRsASZ2QEKi6insUT
KTT4V6svfN/B3jfegoxOxhZKDTVfhNMpfUvlnvhdCvWLbxA5vgS6ce4Wz7s6XKH4
Wo/Id4650o1qEyS61suGfmvjzyMy7F/tfkZiTx/KwhkjpJQr9w1e/G/X7MzUOzxW
c37JyW6gcK31d86DDvPaMWRwmuEcREWb/jRMbYhhp6jEeOcbPPb22mvmjeornvw8
uuxh7K286boKazz7nmcyuevCOXFR/bY9qw8Zp5ktGsvWGaAuxUFsj13FWBTE9MqQ
xcgdYzgpuV1CjedKNn+IWGEV619gwEsOqaDt8G5yg6vntwAK+h2truBEYhEqiNfy
5cYiyCwjE8ap8S+gWLmy5vlkGHiXpEmnJEpMf5OrMcNTkHITvfyuaonIpgLj+ory
KNYcvvcmk8iGWpiPF07JHZplS2sUbbiK3BfeythsNHQnHKZfzP2/98Wbg5Xmw+tR
XlX7kJwYd6ZFe2zpCYv8BqvNnAFOn5Uynbyae1ppSV7jyAxBCpX2V3ySF6Gd/ThF
acpVozn8bWdoRP8s9VaVH769QCipOQwtyiqWYO07z42dif9MA4JUszcyeuHlaJOb
1OO1hG4de4TIzmoy4vPZzlBUqNkeA4RigOwBwnx+a2fwD6qxZFoxKQ8YkgtHBJB7
kKMGDG0K9AnYIvVeb6LJVr1p4uYGu/WXr+CddmnHQ+sBzA7Gt9W5j8q8D/+8gpy1
uqZJ9k6Fv4r84GVv2nwXIbVpg3/NQhHl8FNXq0WlG63XEjEr86//bKJ8q/4BPEH1
+6gXF/uQ4lKJ0cWi7b+Fm/1y2pHFUYulx35N856dKA3SvN4VFQbC5HLMfPBm6wOe
N1g+uts+AwiW4iW3XEeKgt0v9sCAstPJ9pfCh+zPo70OCf77v8aqq9CbzViXFcrw
kRFMo9ojc46COXChewh6CzHRjRkgNGOWl8NN9cWnxYndE+FUAUKH99xHqEbKeb6h
3wR5AWOq1VT3mTLqmLyL4C0okCz3JBVRKBkkAZhT0hxExYJ1NVJZ0m4Ho9mP/KeE
NJ1xNqOFXPOI8zX5YXxoRjzjVK92Z3MWEGsrJuWvYaXDMNILTa00jrwRz650e5Gk
DwTiIFip8ek54gCK6PfBfOjJsEdLClsKn0aEUumh3ZRRzwiyG4wwZVd6t+qfP0M+
FYvQlx0e92+zcR1Xgsvl3WJeWAVo/KCFQH7kpedFdzx8vmt5hCU1pDIhJmj4W2eY
e55Dm8KZhNr3Eqpb7HilLE6z5GNCh9rFvLCO+ZEgDJZ7srbCnlaGEnxfiNOriEMX
EoMdiHxocwfLe+HX5mhCpdeXx6s4PiRuczMJTjFavqGGx+yQLOBDUyNKAiVjs39z
8IpXyuC8hr3U2ipDwNNEsX0yEXGDMXRNgn3pnO5cTzGQnIEqt0bs1z+ffmnIOp3Y
F27XCjKzVfqVAfYgYo29x6lEWYfAZd2jt8HR+pXePOehFbiI7pRIw+RZeJaqRKEV
/8Jaf5cUCeS2WyxRDP7JTzaXCimkBtgrkw6kyHuD35LjE9tJrqsRsiPO9i1A2Bl1
KTIJtDcsP319/HFsAGLdiN1hJWdOh17rq9Ob1MkQGa+srBLn9OVGE+0bNNtBHLel
dtQflc2bMWz1XHwsKMWl72XZQCv39N3DNCmEmpLCWgLZLbde36jWDAFdzGNPdbYs
xu0FiCRkOvjeKuqfFP1VvrxX50Iqa1P5zqH83xhbFH7C+LJOE8bU701cnGzRe2u0
13YLMZuvdZBbqa1E2Gv4N1jzZkGXTWBZ7PIMZ+8RJ/qjC6IWdRdsLeYCVCyZZfs1
AKdt4HPuxVbxt6pjw3FgTHMsJMtr+JA8N5C7DQNaEoxxhO7k3cuRhoLJuqr95eOG
ElRgqaKDbo7KuYpBQlasO1XLgi8Yyy1ekOAkvbjKmFcXNQzU6+7PXHnMTRZhZHZt
Z7w7U6kSgxh3ucx/MhHOaeST8vd+eeBY723iNcRpj3hp+bRaEfndqRSALl4FbNLx
a1HgpumBuhSg4bQwk73W9rmYcjB36MnowvFnDJOb5GHOF6mcuX7kJNfmGXQiqwsX
hXEzA9udb5Rpe2eliZCMepAnu5ADGrqhjOGqdKeJy5WxKquwFT1pUB/UiZ6br0ON
Og+P1+auH63FciJm4Kyb/IxAilglvNC/f8uEJseYUqtMm6aqbTtQ9EFs3G4uCNX4
cp1ZqJX6s84EuMkEfE/zb5Qg4bBgml3Q09vhxc14uKV9jyj5P4oRiqfop4K7NXPa
7Pms+Mzs95LZJp2SvYdUNBGqOYxXoLdZAUT1IjU+/VIjGFFixknrIxAGGftSa1Qp
I65nCqtZ5xSEHz/FoUlyrIZe+G3CRvdgjQKmQAh4cBvOA/EcPoi+CbLO8PdXx0kh
0vUq/YE+kTdkz7Nc8Eto/PH/pPNuajaaeLLCT1JLOHQNfhqziDjt62ufjTp+xCpM
7M2AaesMXSRu1ttmsptxKagfdYLX1FRcUMZwElbEtKtV6BphKWogMvlMUFcDtWh7
aM4HhP0tG8T5AC6CJIl88v1smKYIxbFPCRtMdeu9vdEcH9d2qji4sMeQ5WffBv2Q
eS4V0GmG7IRtW/N4uQqX+3KPK1xLjAwnuAM4XnxsTYea1yaQ3p2eBc6X5pliDL6y
KnIniGKF76EIqYUL3UGzyo1rrYUrBHPcoZxBd0LKq1RIWbvZKXFOvlwmySkVELVZ
TsCQaTeCOVgHNa9cgXmrCaVaj8koNC7y4f4peUG/hkcvj4j6pT0UGaRT2lInrGim
rv2TXaj0mEvW/ekVxuenyOBSTBEYGun0hpOWe/GFepH0hWz7YUzC4bGr4z48Pjpt
RYKp7rgFEB9YO68N4q3lGA5akPDflibxtctonBzO0zKm74YnmZkTdwru51bqB+oG
ByN/MHynFvBmMzirC4Cwbxdd9oqwuTTXS3RkDNJi7FC74GIsMD3W8ctiy1/BvyH6
ch0VOM5qnDHYoOFWU3uZa4+SW/uvxB6amkBt9aeSSv2Mn8w5W0R5cPMOiET1BJN3
AeZuImD4eG7Mm1cYiEdedu9g1L6OEKkHR9hEz30PRhjjHoPDEC+quOQiZzvydwm1
u27ruJpE0qhx3iYCuUcvWpCbkp1vJxfxcDulbpoKvuzKsUgnWgpWOnFxXqtdXlsf
bLu/dRYM80W5U2Lesl/fz9+GAKhztHFWpcm3S5YktxtZxXxTu8iSEl9aHuGQPXc/
u7+km77H4nSfockqwhSWmCyZyjLB7CIepleIDTumBDZN4XyjYNz1DJNIGR7EvuZ3
6xih9kui4v2kldKLANEZsK/s6VEtH8VqpTdVCIqbB1KLyNrfEkmS0VtkiXqyAZDm
19iB1pzlL3ACdZgzZJ6JsjmnJ1ugKbyCiyKnK9kwF6yaOGNxrxBrH0g8x+Rp5SBp
GABEPk2NPs/7gCpXnvZzVcN0W6wB/aVmwEN2me5uoRIPA2NM5FZSQd54ezL6djJB
JpjuIcGNDx8qylr9Wac84PgYRh1TEY0DYt3zTzc4/4AimNNvlJRMhXZhKH6lZAgU
VjuL6iWaNn8iVljaSJI6jv/qPABav6lDmwP5fGSmJtaOnL4l1/A0q+S502yTAmgN
u8ro+u1Rx3QxejhM99fO1jDdoKX9uSG5bDOpDUi8VI74FUzrLcI+e/8rJRvuo+zb
Paw1DYaRWPG9Tb+hHLJjTYgYqplJY2TYJDf0DwBhwNAkC5eVnQkq79/ndQz0BFdw
JzoJGG6hUl/j8nR9fELQ/IJBBGB5EabLMd9gzlZAY5hTMKPnCCm/Q/vwMLuL28BK
1ev3WC9bMHGbonsWT5OYwagSbpEeMtw81mlPj3WwR4vGLcHC8f0o9lAOKkOuJ0MR
vRb7V4qUprsV1Ysb49OoG+KyatKvFDwGZ7I8fHuxC7TgZu2wxBaaO0pY5dBS52NM
MQUIQNvHQkZGHWpY4nI9LFCuNgjlzPqv6P/glv/AaUeBk1Q1pwfPC8s/B/TleHJR
0UYjGWxpQXdUhgqqqNNqr0bSCmVUBOxvtMu3CQ5+W3vjZ9EXB+AYYJUcI/NkkK3q
B44qCbycSR4q03+SGmnViuppIJRf2qw/QX0pM/jhyMK64FFcNDo5VSKHuLjJ6v0w
uAS2ReScZ0Z5yAd0F5OFxhQA1nmi56SiUO9MdcxSrLE040xK1hcsAWKR2+622lYI
Lu21/8MQLf08jCycwi/eKScyJUWz7suffJasUazympTCxqeqKVLDNXjfTyuUQtHi
bia07wwWjw8X1RxJx9WU4LAnK1Tmz3TmajZj9OS0FYU4NhaMID04XJwHS7Ra6anx
nKkriU/mvdiDN72YhwGdU7htC48eXbEZ9T48fXIhOioPFmGe0A+LWpty/CAumkcm
YDUaAnWiiJWoLOY0MIm0eQxSYyV5nKM/rSeRNEfh6widXWs9Ll8NThAKhwzwKz/0
Oh6EOD5o5UNRsq+EzKNPEtq4W7+c837ikpCBPCHaDDAa3zdncJIG8nuLHyXAs9Z6
EtgsKVONBhfeJ4CW4SKS2N8wl9qWNPuFV6QMfe8cz0aiHQ6qbN4YQU0mVjNCxaAu
GOyx1wn9aF1AGojva3pMwbQeG0c5JWhMMB9nGkxuv+RUaJsIuMTRxRf8QFERP+fN
OrjxEtFXqzs/OSBJvJ0yltdlMyFaJzzx5idWxeWdMCcNVMy57vNb6WWpzr/TRqyz
TJMADQP/goC1YrRWNNHbfp2wDMtwpS82A/ZslC00gc7E2rmc9ypHPM/JS3fO/4Iz
0Wgcgz5+Zq3DRUglJgeVF937O0bm8ND7KJz+rbDdy492LKeIoxdVAyqxI6XoLJ9D
BELEOB8Yu7O+DF55RVd2mhhVFPqq+Huvt9gwKa3VP2gHeWf5XOkj25RcY6nVLdfw
ujAouVwCEgwvEOw8m7YCYj3xaSWUTQvga2599QHjDtiYppV8oUZ9h37uNR479ehB
l4obTHv8Qfp5b4zBFsFYk6Pdw/zZKD7fZl9PLGIyebrhzvsD/oDgYb65YrBGNYPK
x04FsWw7iJBjeep1w8NnbeDd2Y9oAqRQtGRDD0SLuFu5sT0bmj4d0xH14rsgev7G
tEQYPZdL2TQQMH1p01fSupLLtwgTiCTPVoktQdpjAMmrlTPvDFe4tZpJEPeNg8gY
Tt+WEYUNdVqzqtcPF+vLyUEzzYcTdcw9oKjZVRg6RlNoLf3ovbb5X2MAM8bQjZXj
F/sREBWp0pYKzLFVZyJvwX3/LXe2RxIFqYj+UiCF/gGwQRfqfJo+Q/kpThQCIpXt
KjhqyS1BsrzQ2Facyf5r/kV9NC7tg87pSeDQW+S5piz2xAkZp9plMAn7iEZ2KU7c
W2Hjts3zBqndYveGmw9EyiSkIPK2s57eMHXSXNK4qSzIVlLf1Eq8r1TGX9j3iYei
dd5LThBVJcEdbdo13hh03TmTmIQGZuqFa56WvHmWvODsAUv9A7N2gVtz3ZFW0laY
UiCNj6W7w+LRIxP9C1oBHpoOchgPCSJxQfTAAiXynAvH12GDsQnFyZus0FNvzcdV
gq4R7DPx6wjr55ZnchybUxbeIxydZeyqGb74/I23B07tgGcmta9bl1Pyss8mqaFi
FPqOzk0dL8xaD4YCFizFXl0fUQvVdRGiGqCxhi3Oo0Oth89fyTlQK+uWIPvFli+5
wDFpEN4WGE6wcObsB+PusOt4HflE2n847jb1ewG0sKTj+58SY3719dqAVO7vM8Xt
vYwPYMVQEZ6dp1dEXwh0tduAfxfMdIBRQCLTfMm1jju4Y1CUcS/w2S90gTJ3YIui
KOd9LxckgmUaiuo8BqPqVR+J73CLyvxsOm1VzSi6oRMmt906SiR1TKa30ptcZMPG
p1Of7sZ2MqMo7a14zIYKwszWG+EEUfdPqQ6qRl5IkcUYApXU1wzjvJtNoCw7Dmg8
xrGxbarMa/is/1avYz3GPBFSTbZKzm8bNcZ0A4g2Y0TeS9FVGXy4YJEqhWMeSqW7
MIdlvTKM+6ILHA83/Ud0OoWE8wPHL1ECP68qRnXF5HDpN7SVJbCKeQYDFS79ppdr
sgw51HYd34mtYkU2/BNcFkpA/Err/uknHoxdmSdRiIiQl4tERbCIjntbpPmFjJsY
s6kxKLiZNmSU6mFxFkqMP9OmJFPF5R5bGA9/IyfoyeSelQxKN2EgVnj7ssb5/og/
ywWpP7Z3SsUSH9bg0iJhybJdl+iLrJu4Rrgbyf78zARwNWg8wvmqqupebuoYMRL+
EwN/dpjvu9dU4/0P0+njoTHI+I5jY4xGBJ9Pqqizb+Xvc/v1CftVTwuMPwhAkNXH
tttfa6ph1SFh0ziBtkZAnKmt1wlsnLSmqILrdIIiXqiAoA5kuLc7nR5NEOE7TJXg
EsWgcCCHj6wnGE8ZBNAf+NBn9TmFCRpw20wD7GoTYLc0t+Pmb6zvQGhj3p7oqNpu
pR3bhf3P4qpAu1sYGxDjfw5mJCs7ar/zU0tb0OhT8PCF/+WjMZAs/P3MEeiLqNn0
h8dg0IfnDP9DTdwiWdP2DAU4ZKIlXaMpyn/RKOCuLf3H0NFb46YMkR1K7fcMZ5dZ
zpShZpCO+Q9WkFuHZxiBxq3U8pl9oTJTyr0/35J+2AcjxV48NBtPziX4+NdoAOoi
Kk5k3aFqFKMGdUgQFHU+jjGQkUlBxXjQKzDaxADQ1+KYbpd3OcaVxOvhC86eS5B/
sCPv+y6M6SqPXnKv9lGq2IESQ7eH5jOnRPAcnz2idH2ZoarfyirXpaZXOff3LvA9
kdZuuyqXZ52xCO2WMTXu5pgc0BEmXWHEGE9o2UYMUEhcSJLgBxkZ4tGPCu0YSr6K
sXOnE1OieGjD0XACXP+wIbrFBCWQE3B/CzziAU+H05ZhD4A1UDRAcQzsqj82ARMF
OWCwy8GRwHH6404rNXb2MFhgR9aloTzEv9INLEFEBnuGDCkE6FcInliPhUjymNzc
mi9py+hXS8b5Nr/FpBdGoyUzCXj8aXx8iN9l9BjGKR1xkEp6BxgeDGjGb1bzQi6T
Do86XsOZSwOrOdTCj9lotVmqdB44y3zF4O97GxVBSCL69L4TMDKqogUiSHa3qERF
uQumIzEaEAmMfw3yvKYyow1IUYknkoL5CN92w4rBp3cjgiV34YUwZe9MrrKsLjFW
4H9nhKzsfSgaxaqgLIldZsp4eeq9esqh0X1QeEWWAUgbh0CTx6aGcK58EAiPllmB
dfQVDdsJJGQuuxyliUD7oBK8xpof3FaAoqQKF1vX0lucr/YZlqFtscK096m0tKvz
1SbgaUuGN2KXa8pcnE/8uFqKm2TMEUus5L67K8FzTzDgl4GsVWODQl6B6ps9GOu1
dUtWXjBWDF91ZOeRL0tMlAgT9NCq4QGlSirtNzm/k35y4vmBuD2XNSQ96/Xmk0Z9
O1pzehPp2Z6u1PwB67MbhSoBFw6VyqIGbUrAgbEsr7zIIu2ztmW5TCTdPSjz+BZz
DMYPI0VJpR9Yo590IsgplJ3nqN65dhb2zasMjPpjXy+CR9SRbFZzMMpti/7nV4Um
oOwamLT2zrsoN/MDSZeVohaU82ZPNjZ19rN/QX0KL/542Ql2ls3dOz/Do/mOOkVW
J9B73M1W/apsppZVt4XoeTGM9IGTEfcp3LGp7GTtsVSvTNLhJ1Hk5nRC2b0IIwwD
ezdR/R/klM1FNP95bdIeMQ8vgcqF0uClsGkiEmygPwlrH6W82vvu3pdOkT19xb9w
DOxfJ5ufm2GlYAWAXjaDKWt/X3u1DS6wJ+ywNUKWh1cmC7Y3dgrBUanvsyrllyVr
jNgCJrCnOFiw3rBw8cC36HGfzBK7pv9XZ+6KDsAFZEjQK3En8wqXh9NURPAHQA3G
hdX3yYfAGlZLKhIB/jqt42xPg7d4wVkD5wrj+DJeuCqWJDpta3ZyiWYyIUq4IxJg
nlnJAiLE4R7tOIeGTu36UqgCI+TxHATDKFZOexyOZ8GW/5/stL7H+YRaAHo05DDB
FYDcmQlG5GHC3J+sryR4wloJkn6SKJD7AlaMDIQGXJ23BIOo8NDwJ82En14XdkeJ
I7FQAcC2QoAYaj0ojOsdHN8doD24tYnY1OmtqNHEv9odE8Dt8I1PeWCb0ivTOi/f
yo/Bh9E03hr4kfiZcSxM5LjSfwrUPQBP/CFERoLOFx6WmyUWI0UcCyB/o94m2sZ5
kxt01gxoAVqoo4FHhWKBzIeF0CfTvG7L9QCnKZvRpU6m55BeC3d0BoikqRzSie6/
EmZvXyNvPSP6l8CCcFvECO8etezJClkgYeBT80pf7VOsaaDgfqAgiBHeG0/PmOBT
86jKo6sP0ZojuLChlGFa8+BM6u7lwtV61Ggt+Rksw8po1IeUmZ7YN/5mvrp6qxfZ
56MUG0lDNdrxlLNwTGUUBkFG50L+VLKy5V7rJg8q3MGBonOaSP0GGwKZVrhvAhlK
TDHjJ8abqzB6rHY3TC3O9yBG5Gzah00QAOqdX6nHBeBxkdcCx/0mNJK/FbkBX7Tg
m3+//vrPc8ISyafQar17yDoVUjKPe7Q72nU9Hwu74e0ogEgc3AbPzpawPtjJVRLc
gnLvgBk+JUFAf6gG17TX3MtQsgSF7hewh8TtFKjEty9ZEzZ+WJ0JyBVC8j0ebDcV
L4nEwXFBRgNVlIFXNK7RU3WiRsD62YFyrVbCOWIi3o8vVn+BzVAICl5621uPnSk1
Rc4k4GqL8deUrW6siULE6KbDYuGRzo6gk1iUg0evC9h0dIk3lAeNnReRI9ZQY/VH
H/IjO8U/EXGyeNjL/ResRhStV57qb99MITeRNn72fe4voHHRCxY01a6Z857xWvwE
ucQyHM2Y3CfuW5kBUchmt626qq3p2FCA4k+Iq1SN3ArffcTpyq3sKDETUSFq2zzp
pa3Xp2SspqAhKmgv/LG1C4WYYczGX9CNUxp3l9L/Y5i0Gm6T+4J5NNmAM18xOniV
GUw2C6bmobPyKf2UB9T48kcXA9zlEXtwkoYC8gfgo/NHwrVRPea69pXoGze1VPfQ
LjhVEbu5euWuPGoEJpuQb9/FDVo6w/Nt29C4x652jBY+wkcGT6MWkMZttpDlDTZC
yxuHEXLOsrrihhhGyg2r5qzxwetu8PCe7BHEYUd7nDwMeqqSLhf48GfULW+Sufxv
VRkXkuEG9th5oXvgWfEOrF91zXJ2uUpCvJei70F4kIf2+FlGOQlmbW9shmBJMJF+
a8dbd5RZdU7xYm0SKLGXfBjeUnPnDyP4OC+DAmmvs/9Avz3dEMfSgj3as6rIRPJ0
TF45eTUhzP7t9uieqtcRE+3WxxRXKBQ963lr+xoWvHgB3eLNPkBcaN/6aDB5Y85C
F7zDIe4GuWDQPhc2CUbtKF804IBdmYR1qejICPrp6G20mMy286ipRe8bQeIVusRZ
7ceDuQyaFD4pRkK5TuH3pCLxVasLGPoeUTgZI/lb/NjK9rE8+aJh2Ow/7RGA8+SK
dD0E+AwQp/y2iSIMk7QzW5xApZo8kMvvzPcmsiMq07FxT6WuryC64Vz4KpPqEbx6
/Lesz+ZnDCFBmyrNE1Ck9Ak47XrF+qc5zPfaNqz0nL3LVtY0o/Nj/rHtyKAfd7J/
Y0l9D70GqpGfQjKq9+w4JeV5VAbh78ubkAxhCdKQzeNf5FoKiqUwJOawJY3/ya5G
9tfFifWRqdD81zSBJeU7lC75Tow5RiEsaKHLy5NE+92S3BghDxi/k7dkNHLAxjfI
Gx2ypvwtgBljNCTBC55OunZPCG/LSbpYnYf5ZCsRRwP3vl2kvumo2gDBcpGrqG2R
SytL0DuwmXeRQCXjS8XNakC4Pgkaw/umRHhts6ydVf6iXkeRga+/ThF7pdPK47O8
+gCFXSDgR/ggBpUiDnwji22CLVePtTSzYUpoqFzBbZdyoKIOuEXxlaQ9qVyw6Q5f
WJPQ0y7zS+b8gLFW+jMlv4sFQFJ+LZAP0E4Sy65568f7aN/In5D2nsNMa/w1UfMO
ZscGbNyPqIY78TewncfpAmpVXBdy/0zvTWea7KojhGuP6j+nMdAmQn8xDZXftaBY
/UsweWjYaJKctbt3/WFDW7Z9L4HFTrPi+rTNjATVu2ytlQtLVbAwhPhQ/Z9PZTxO
tdoRr5OZPDL+qaXkeEtGbwmr2fiobOrzD3KmWBUgf2jAkxffORwwtxCXW4Wn8tyR
xlXg0N90pK3fDQ0qMqxIxAAeS1zcJfrkdxlin5524uYpTXdfEL6rmcg3okjvYxJ8
IdIUDe+aNN0WMc40MI3zWojDvOjHrOOwER5wMBk3smG36bBLNeYbQok+o9EZ/kVI
ZwvALeydRNBL0hc1MS+uPXpVI5k1R0HOkvjEPWJP+VX6LgQ91czo9Le2PVrVI+L3
WAD5WfQ+bXTtqXZLoZSPRaS/z6q3Tmm7mfAvOr/3e+r86kegyeVUBvlihO1Qc4Xw
Yc1Uwg+cjOsnD2X7G0/9eP2CGFgmnevx+rJOSl/9QI1z1Tz5/wy3DnQQqCkXnvOk
/w1z0CHp/bY1Kfh5dkh9TGnr1KmF3wdBII2QHt0aaV/SVSb7h0M6wUAAhj1TZRex
xBB80pqAE/ftawBTX8Xu8p1VSVR4+q6IqnVwivYghL/YHYfL/8An0kmQI5YmT/wx
zCkMECIXYl2gz88rN3zoF3oNJzUhSeNCmOiKETjzS1uAEWEbmOnX/YKK17tlIfj1
JefMFKvnLDiFa/XQE96aXTjAXMVNtC3i7sgZNH8euMyzd0cPYp0A5ZmNia4b8N9w
dnc4GajLfTtZbCvXADkbR2pv0yn+9jUpr30BSzCT3ZWjzroVdBGkQjxSPV8bcWkI
bPm9XTpDBBud/VCJdLxKfY3WAnR1+xwWXRVfo7mf5UBNfhC23dJRzTi0pqsW9e7P
V4pBACAkt3TRrxS6WhQHmK0k4qNKS+5EdPFwtTn0DZzdZSOkEJ5ie/wLJacm9l7P
C85U6HPEcp8thPAa032KyPiW4/vqLlXZa4yEjgtgFJA09BuDGAWAb8HFWrYoPXtQ
RXJC/TEswP1RqtO8oFB8TQM/okCzx+o6jOHOeDNNnJpQ1vkNpb1caETd/+m2ukH3
BH0JlRP0NB/ECZhlMHrz5Nz2I4Rur5yrCRLHRwqLkOFIRyhX7Nq32do3KT0+ASU7
31uxF4W4b2pMj6tP1CeefQDqwchUlJz7oSKdRIpdRrNbXt2wVwiIxBkWJArP5Jfr
tEUrjNQTC6IfS70Hg3e6S0ArojevXW7Dl3wrHrAbLnxsGXFdG2VEaGPtEaBj5D2l
CGhzk4RNm3Mett2s+B0LmOW2a7+q0Mf9OoLhX2w1GQdUgeT5TmMeqSFkqYpKEodw
/5CF1WuX57D3DZjFhzLPKl4sXJ7Wdij+/2p6JWTQmAxp8AuA7ZGNi56RRs5HEChP
0qsWxo5s/eNBzTvlwkUue/P78r5JobEuMATc1T8+HW9ytw18+K7YT4wF2BcqZ42I
O5kk5b2dpnDB8xwNszqHXOLkDyDdXQ782wiYEDNcVpI2kaLN3PxGmQ32SrVROccG
7ktxzMRyqVkVBAbE8KiIezkmVsBGd9T58RFUxSVmqfTjW1DasDDE3rPi8pr+u/pJ
LJGDa7PwkwHQfirpP+l6WPyWw4PprSj+Z6hq12jIXXqKOnu6ryM6vpmOe5AWBmre
TbVfpQwb4dyIjYA3w7j3iaQudlgFn6FOo7YPsI8NcdXhlxzzC/DahdGKNYITu8BV
STh2t56Tvc+AykWWR9NIQzVJyyvTxx5mn+kTBNSmSTluKvDlQeY7Gpn+Sy8LG3Fd
CtjCCBRZbvZuNe9v6Mlz4MuPtd9RiYh7LhS1vdKgzzAMxQ5fX/YhkCuUh7ZYVXNd
6EWpqrw7x0v1n6AQ988bu8A003nudWj9TrS4OeOcGmblPOLbh+9q0UdhFNL3i9GS
VkaF2FuxwNy071vy1RG0+NaDbffBhrGgDT2Xx5O0byykmWkoRe/AAxghMSxa+77S
SxX7DHIE1eRLz6jEWSLtnEOAcomBlyy6eTzvNJBHR+UqTSNltsayQv40VM+vxJzv
YkVXHWMAK8F/FE86leVgy/A3pwnWnBYjsFI1cUkAAUxAFhFkr90Yd4oHOuuNF5M9
w/HnsicN7rd0v6+V2IS6DjVtkEfCrZXdMl2ORmzs/h2ydH0MwqH1KTPtHmQOs4Vo
FM13MjfX66Ov7ZVRZWKOm5+gEEA6lg2XepRwSrShBeEWJ0RSD5VIKWErhA9DSUu/
VGNYoSctsbmE+tnGFuwA0bSmeA8D+pqyZ2bed4TTqMC5xnYY+fpWdK0/bSmK+N2X
CNrYDXVZgCdB7jQDZ8ZtwWBgZ1F6zoSmdFOxVeg8A4P606h+G0rMBkxkADxnNVUy
6kiUSkUeRjPTVGX3j3N+DDJM7+HbaPC6JOoLjqjFYD4OQb5VTqNkTB5t4elzi6em
lk8lF52s2VVWnVPldpmIrrNWTpjSDqBma+bInZiiRjhwk4Cwl6hqcnTQRJAHReNk
fDITvZIMj4YEY70mDZ3x++LjxtTtN3eT7YD5uga1wIJkBuvKN+OkIFqd7yftIFSx
vdJhiyOYCrEreZQnpqgD+rqjmrO94AvOLdsXJ6YPWoP8MAIRoGBnje4Af/P5Cuoo
0Fxn/ExAlQPrMZeZjE7uYkO//D9CBx9SzajH8SGAcpp373UAJtUCGsiNohm4PqAZ
u0IWW3+9NmIs34YeRl6/yHl6fc+e80phNwM6v4QoVGbCF/CqlVfXisyThU2QyFQj
ABGkrv69+PYExd6dreklak4dcMYbQOQ6J4FS5KgC10bkCrzRa9ZubaK4BWeoVjRn
duuEElHnUfc8KCFxIRGVXckIF0ZqvrL5c2pSZLDHdxjuOXzvlVAM9TCsGc2u7P1O
nnq5GzQFGfBw35B9OlGHFVND0azk4QLiYmeBu/JYpMqB0dXySSKjYVWd5Z2N+o0O
hm5b+C5aUWGof8q/lBe6MxY0eaqJpr9QUN0LGdKS4Aa/oVSe5ODj9f0F32GjURyZ
e3roPUZy2yf+h4/7g+Xx2Iri/VBRzkyMrbvYFq7d+EcZwNT8cnMCbuoDS5PLWbcC
eeitCcWPQASnQ1ewORI1wvjpZgm1ZtGnW2xZVlRHVp6/Ow9EWq1z5BtYxPf4IYCr
tIKVbOkxC5t3koCkrc+Xxa+LI8pnzr3FJRhhTA434XWird4zvALohR9elklroMMF
Xd/TYLLdxF0dEMIJX1hQ5IaKZSjFfzbEjf5830FSyfkFeMdPmE2K7URM27spZ2XR
1C2DpfUmHQbXOhhhh86upjN4TAHgyFo7cUNfMFm+QBYCqAk4igB2jxXe250A7JIo
8w2Zf2ejVAJu9iOrtm02U4X2VKp52aIn55rsQ6jMt/xz8w+5Cw8vcn3C6m3yWkUB
CZeA9VL0UWbnTfwsjgn4nt9gdKJHzVwTccB1I43/uAyGd3pZy40gxgnLhHcXgj4C
qRNxlv/1xM8ST5UyPLplft+/E2m1TX829uaXjxu1Lm92xGnrsFQkft+mHoOF5WVB
FRqP22TH/zPXiYfyzKJnlYYQkCR8GPzqYmCl4ofcJKtN+3Hv+XGO5TIeCkJcwBNS
HGGpQP/V8wCHz2kR9PwYLgT/U1TGBxmh3V96y+grON+YrtKQwlmrrM8dhshIT58t
c0NpJE4DnNRWWx9KHB4jwQtL5lakoRtwUQvONo1venvkc99vrhWFSVGgkttdsLDH
V+Tdw4+HU1W4uIzYFqeGtBE5wPXmdQP56GKMowjQ7c6UNtuTy8miG19UO0HSkapi
RT2HaIZaP+u6G8u8MUcXnkdR4yXUFfVAlt0ehbfBDPGeXGITAtibCZomfqJlFlt3
5sykMF1uvQ5jxbW7aYECxrY9YKxNC0qQvUQZIYzFvCRghRKzsQ4MP2V12otieqk9
EVZO+GRd/zOOnROgLadPACYp039h7hmh0VM3v2Mb8XABdQGZHWZT6BMYTZNG/E8o
anX+8VxVdNtLxf41iiNS77dXCc83TNu4ciwyyROqvRVW2B4t9YCE579kx3nLWxd5
mLisp/btGRjl/MQ9jyxgPic6vqdPSI68i0sAN/QMBoBTGOiS4jmAJ6fYZjmIYFtF
3IVbjPzHxoIR7tVfUalcqLNgL8Tgi094LKhCbpYrPGwDxScPSRIPiZLbIn4kUVPO
GdCVPlascMKAZfk/8jUOIDBSq/UYM3XT5MQjGamfUHsPogyJ7ubFJwsn7X+PBUzh
0SpbkF7v2AGbeWeLyzJN/k5md+QeCllsZUV984e2S0eFBXuRabQwmAAcDfFEV493
EA/B1p7tU6DRmR4YZxD4DphRXoc8g+N2GDDdTcyHBEGy+GeSm5xKkr3Gmeoh9P65
LYUfUUKnYofukLhMgkh6JmrwIcm2j5vz1ZNgqW3qZmY8pdGMu0H+VJbtpyv9YTTt
YkKuBjewYpov2vJe7BcJG8HaV90u4s4rRbv0ZLkaTC/2ogri0Pzj4rE9G9UopL1F
2uo75EfDh/Dl/aPHWibdG2bfvmtgtynMeRJzH41i9fo79vGw5A1W/05woSVKaxHZ
5dg9501RvL8fFcE8p2wPgkfORq2AHdM+QMBt1PZ0jtE+0Wo/dHS2aajGIIqZnxf0
BQK7yLWoXXXrsVzBTOntopeMCsqHiKGM2CSD1Vp+KsztQ+6T3eBzOg56OQQx53lE
6s3IDAQiefnKjl7mydqzh9yZ6jSccefVtGN9gnhBdzQ9l2rBd/PwyD4T3yCyJ5hG
5u++tAmShOeiKtR5T2xmm4VJEv/LSThfk12YYbroO/tPeTB6WOuz4HnfJYBQqETO
b4bUN9sLt4AXp9JtnMQYM4AeOj/8fkE6rnzAqRz69vywLqGqMgdR4sWltgVPjN/f
IOtk89mNTcjfDUqOSDHukf9HVlAxc7VvAqxWawpF7TpMM0USwA+NCssNQLOLK2cF
uHd6+WDHpNAIED/dp8I8KFt2FtbFStA2BngWVcOjMg/ymnxv8uEU5A1+RGWE3U/Y
sQiqd5HKc3wOR5zq7gjQ3/k0PPOBey5IdcEcBMIrjmJY1TrR/X0uLxN2/8A9PgCG
YNYu2UwL7ga34V91RrL3hIZrVcCvLPnJccpNeq8OHfl1nZ6isSKFTf6ZPZd6Mh57
D6LtSev0/mUxvD4jdsANoQ==
`pragma protect end_protected
