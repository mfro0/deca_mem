// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WlDXxbqnEwNdscZD8QF7F6M8gO67OMJa7pqkdT7KJ8CLvUIvS95gQTaT8OcniXP1
7oDxBUhRU4iIIDCm82+TC3kfEFNYEkw7mdE+r/ziCC5o+yjGe1X+Nwi3D3/paqjo
U9xEx6PDgzr2y8AJrvHmvhJZtY3bs1DUHwESsFvydzo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18512)
e1OG4N3wtXfS3kPJPrpuQCTmiHHBrd1YCiPBI2kFQZLzpuhKYbH7atWHKEQAqgLj
EC+YtPuMvA7a+AX+ELHjoBB8QTjQJBKy58G1ozbhdQo3u09sxZ8u4GT1zYEn1atT
Ni+Pozdy9pnq18xxjW0zv5YOb3ZgjnOapAiEwbNYiFpArpCk/Ao3jC9+gdP2cC6x
HlpKEdvg3xqmPusi8BFf9TapGllb6+2GIE4taIhMW0l+e33Lqdvl4SgRB/vbqhmG
nKCGKDSX/eUTxMW7CGhATkRy5tZHuYFON9Vn1KtWskC7cJZRM0JLPB6T/vHgrWOP
Tna4m+iCZOEUTfP6pbjL8vwZejE4ik/Ews/RJ0t5UnVNgIOBBue8P58ki94AMxcN
/fq0fELkxLmjqRXlJ0Y81Qzah7d5o/1/kJRWky8fiDW8jtxUoKmdCcwFX/+Cv9be
wqDhxpdIL9elHR2gJLbf14qgLXqRaZ/4WYA8IHeNp/Iwz42yPypM3eB+zW9Xitv5
OFwHjV5aNdYKfSD/iP3t5DW8SEMncl7s6l4jxqxX3WjUzZKOWUtBB0pRwSBxnBsf
0MrZCg2Wlfjej5AH403T+zS0cyRK5AgLpTtwWie9MoMmoJ1gGrdzNLF0tUp2NiYh
IR3MkQibi5gCxKwTsylUqkSdLCBgGEIcbGcIuf9daCvkV7XS2mt6K/jW6q3T7j6I
Cu+Url+qk2buDRaxUnpKfG1Y0RO1RVZeehaqqfIkPYtpw+wp/7oSvwAV5M+7DKom
w7qqWWWWUK8cUAqEbnoNiEgYiw3bt7s9e7JjHnaNohjXrnkhafppFvbfQ77j60Xs
RBw67FdnLIOrRmb3csbbKNqF0wJtEDdylAasFE1I5hhldsNVVvu9+8RvImgk1521
JEYXUQs1ReSizUoP6GicCED5yEuvXdt47VG75FxDT4puTwlStROg9URoZTpw3Jh9
sDaqbTh6rjSNwPtgOf+qcwHFe15scuVFmSjiKIFTTIQlz0upDqG0zX7l6AK2Kj8x
GL7rxuMQ/7DKanZm6g6/EloYVujoDv671g5CzLFbGwbQLCRMFsgoL0QHpnWZyWkF
6DEjt+WYT8yz/0Sp4ujYxNV/5cWjjKi3NIXwf1UZes/TcYyzPMocXJBxIcbpUerT
zAxkVPuw2LO8a17x/gxD0z46X2hLNt3wWJFj2LHW7QaKSCXpBR/YfA3x0xNUtCyx
2F+lBoJ2/tsNTccM+PanKUL0s2QfNYOY/o3YdT+jXKoE4HJJP177gqNEwvqyuFxN
eIx4NOaXNln+4oMIy/ypmvlkyiR0sMzatFszVEJz0Xosp2xPw2nJr10a4X13q8vZ
s1ed4DZZ6ygp1Wyjo+BjKciZcOcWIJRxrI4Owp4s+zolkkP0k7Mzhi1DMaxUlhVm
dz7BVV0Z8WSj+ynNu80Lm769SDLzjL7hGDYEAPOpH01FH+s4+ShbCPy4nES5DyhE
DCFGHDLXweg5iF/4IavNo7PU9ZsH6IEyIxJtmpkyqQ8psGId/N9HIItYYMvCvHd9
RcVF/gF8c8koQu6E5LvGbclSvIEdglLyG4foLjDf1CpOgBqpjj4rLFIqcvsfZRnT
+Y3SPTvkOzOPUTkApFQKr1PY78JvXLn7l9AgPOQtjxoS1yG2OvXW9Zc0Wi39VnEa
2Nn0Jy6Mzh+akGLl8KYS7AOcdOPEmo/898uqezPrmircOtqxWAgC8/Tjbq+Vo+kT
7Kz6f0J5K5DvYj/mei1FX+DdRKRjb+3//DFisAx5PvW9KoXoIvVPGBQTJ4qDDZA2
sKgxiIbjEIWz1vbdhId36u7numhZgiW4ojY2MQC9oc2I6LMK5blacckh02vab4ft
FRTgks7X3qwfUU5ky78Gt8yP7D0Nnd0Q+3BvYHur+jkeDg5EFjNmCaDtjq5E8y1R
BFlZ+HX8reRhjMNsWZDKQHxdcWd3TJkz5xdLS5OF4EpQR/b3CwshiFSKfmx/WAr5
k2Htm3FILAohEm/bgDf+Bp4mFQc//3kMI9fcQkPOtKowSs1mzDLTssSEdDj+kKYn
mbBdybarOgltzQsvcVBUWBkJ2hLFMxdsrmcFTiTwW5lJM3ywr08edq5Dl1Ur3DCF
ST4eiTTznBBNCTi2+Pt45A3Bm984mPRnvh7UzEroZyo8fxo40BWIjgPKLHwpiSTJ
in8zC10mU1eSrTAqFrxGH+054D/hh//NxKz9D4YjkszqCi89905TSJtCKwJZFbj4
RsnxJkCnnd05xZb+ybTyBceLgjTb9lTLRXyzE7kHSKf4weTCe4eendkKQVH13Cgm
fe6fhcpgAVZEbh2HxK8OkMT3+YTOX1beSGn5VdkQJg52afCTRvK100qbetdVRwC5
7Qj9hqce6uLKqMCAD2VfPATEvs/KtARxRSWxdNw1qsmhvgviqiQwkGLJbV9u7MgM
HF2AuMUg6FMT+0chey284kg6nb21UyutdzLFPCpLewJ8mWVCCQOmWOxxtgXudnNx
ORQ13X3nX9kXAHyDBBVpIqUgftVAQyAAwRf80/oMfB9ktwmKo4hERbLE7RL3q4f9
Owzj0AgmWsQQYf3EKGza2wB/Ky8ALHWYT8ng+xJHCMFM0k64metNqaKWJxq81hJt
bpkMVACyil4sgYPT4CUkD5RQ1ZTMZoWH0yduNmAZZsV8lNBTQRn8hTfYJ6YXE5Rb
zDapsjUtJeXBJXQ5EGzC87O/XqiPQ0XlYVS189IMQbJfbXczSNClWwmslaenIeq5
aWwtO1jHLO+T4LpjBm2LbyhwAxHkEmrsDBdeWkPBmKlmYKR8N0I06OF7iYhHkf9M
L84H7MWAxBFWOsAtfQYHCLov9/66qpQVcc7xUiktzgZau+kYxkvdyH64NMkeRuGW
mRSmj54z/FbJPnacGCgCqlSMKU0YVaHWgkNKtLLjrtlihsZPXjyRpHpjvSjjIYc6
8ckct8iwnj2wlq7JsiVQAwcjIO0Yjsd6y1fj/MNosx4JniL1D7NqG5W+QUnpQ5Ze
3581t7SmCkATHTEgGAxtfSqmgg2bU5tNJ8XvdcW8IZ61nP/KUfVPBd5uHe1MHlCO
vgKuBG0kyqBueqEnf1LXmZD12obMgUKUtBJ/LysequGH//LATaQ7HQ4r2WvNhfVc
vTMVItUXGgjPERApoBW/dcuLMzUGkhIW6TfR6axlHWPTxtFkot1oODL/jr6opC6t
IIGUXy8cmqELG9BL22lSGPw7o2nCQcGTJ4+uSYi+NYn5eSSGTIEdkzZGRxb7vYMu
T53v3Rt8QghvBguPFQ2gOt+D28n/XKrAyQkSwnuQI8938CyJRsuj3HCB8J4wczM+
kw9jnGTFHn66BFgIuJMZna9kCAuNyFfE2wz6ZfGNjtW1f/xHQkDkqPdTI/Z+J5+w
YIzFVN2jenbk9NqM7WhKCe0xh14IXSagbFnmZKausIST6XRkh3kIhlhHo+Ok+AqT
BF2oMlpjuI8WQeoUxphO32vcGzmu2TDNfkMntBwo9mXX8B/d7jUm+HdLKW1w3xs5
vcRF/5ztIMVtuz9rRaJNTwbMsiTFiv1xDzSoIhBRe/yYDsNEipcrYVpZ9W+1Lrs5
C0bCP+QfkXW7kCEqmMD2LfScxJ3mURWf3S04+MElbEzMIN5dsc6HFFPZ0BW6qxFe
kMfYuJ52peZNeaxj673ku+DqJpAYvLa564JU6CxusT2yiMqdGgkRGybRERDDE/KV
zRGe96zB8JsUtKvmEl/LlC0E9SL5O7Tiql3wrqyWQ6w1Q5x2LyIZuo/cKaZEnFPu
w6Wzogx0E/krAi6tgxHe1+n1paRClh0GpePonResOnIT/J8UqpkCMUkFglgkxZq/
3Mvif+bw1Tzn6w9GdM7kbAMimlVBnmwwkbFp44ObcEn4EwrVTi1bo7186Mu49AHW
4Hl3icLNk/mjMUqGYvKLrxpkWpbVaxFr6D0wF0x4loqH8Lqu3/rCme0ImKpygo+A
fmitioWVyVrpVekzd1ElWLrkxmPBFeUVjnkAka630wt6UgA5AsuMAK9rWS4ly/8R
OiODnBIvPBGQhh2GnlpKhtlyU0vyDwsr3w4YgGb2qNkRv53pXy0kymPMPH3Sr7tM
vycpYDN9Ln2w5cV8Fhh2TAJmXlmEsJud9Jc8OwDTN75PrfyeQ1fAnhHyw1zKauzJ
GTJ9g6Kss6ML2aFP7pdNRBIa2/OXfKgYz7TLwmd1YWcPbL0lyb9hOIVHO6NwUrUU
VizdkwvwtZ3KVyzvaIKaT2LgT/AIFAhufywOv+n756X4HDeDmvsYewyG+GO2A2gn
msjfrNSw8zF//9WmxbgOILQGz7yrCF4rUEjbcX/FrKu5vOfxpbn1tf/c67fpkdKs
aYFJlZmTfhpPKuAF/wsp6ts1RIgqkCi8VwrFoLLVsL8kLp74ptDwmKmDz6KPmueW
Dljvg2bsuH/+5Ep28I8fZvhNi3Jfi49+YVSYPfZAv6z7f2bTUHe/ZpXmHRh8NkKH
pDk+89I/AvLncx/rMgQzoBVJ8b24cD55J9vWMUwtsaI9Rg3aTBS5qyXXT565sTSA
NJrvqcpSO5m8ekB6OqoVK4ZRfQnP4eM62XDENvCUurFWU1gr8/5p9h+F0C0p6Nox
QNShyhwQQAggCDCkoqBlVJqSMOVsUdg3OJ2fq/hopPTJ7mH0sdlMZSTx7OGQGxn8
fUv2LBIA8NbvO5EVzhro8v8JCVcq0MxOGvS8RR0CgiEWWg/ZBfXw9N1wQcl+6KP6
aSsRy8f9p626dlOUoUO6yWIkQrSG5Erk3gZM8YPxzIKFGIR7XPh2rjvJ88MOQBNZ
p2haP6P2CkPWpXLfQvrUGtiwMHRTnuXGHAJCObQPSSEEG+0NrCbO5+F79nCKYZZO
9Jcl38o9aSvxsVOSuN86iuZiVMq9WGywBRdn71hus8NzSopIrFQYtpJPV3wThAMB
RMNFIjJdsvvpbE1gi4b++huIrxRqrZzJeIlDqZI2oAI63dYUWLa5LDqY5TBTUBhU
b9ZDwIlBi0K+ERmZm1LxRIpzixhP6HymEzGDbuBn5+LeCM7qCroAv8i/ajtpb1Yp
hLs1EtrXLDhsi0VtrVnzYBUqzweCnlD1UEDC/dICB4Zw6+hcFNeOIls6W+cYpXDv
79RmZ6WZsGAsUgmGuV8g0Ls5npctgkcQYMctBTSQKXu+Iwe/Rwj/pRuEUPGwkbIh
SG6IQ/wx0/1D7HjXB17d1oddzdMK79ihk3n6/TLbOEeL3+ungRrwts383UlKfKft
7+K01txivR6kbuygR/AzttP8xvINieW/xxpJlIkW9zsxJC9jTDSSSF1Yv+TLiZD7
WV6hi12flxGksKNliUSIlOfI/a9v2f3M2ykmtsgoDZzPzcnpjE3mbNo0rc860kzx
xZVYzREVlZ/yIzwLQKoK8FaDfdpFia7Lqa4hcgpGupml0X2D4XQBsNpl5KL2rC62
3JFD0sHQjEQMiqJMHlgx2CZB63wfTrFPXYcuZ2F4c320RJwOalMQScwMXxCapvYH
uw6qKKcSrhfEOb/GAYrsR6ph7jLMokOqYWisNmyQOYBretYq4XFstRLahNDEJDku
aHVj6X8oxk8h4ttDqGZJc+/NnX7RIa9tEEkddYumx+0+xoI65P85QkJColcKaXo2
OReBBceJdYBRuMDWI+qmu0vFzsdefa2Golb6JhQxGzLvyamhFYCs2K5t+O7HY6Ip
5CSUD3qPk5Pfj9NodghLRfq9lj6MO0xhAfwnmo7FD9LT+VOs/Lqp3QHBORLCWqAh
yQeqdzyTbXb0ug+t32aK6/ur7ErJQ+ZSxfMTKsH9ZohnNCmpBxZZEVbeoXAot3FN
O8xLmtd2y46mQsFz9WjTiq0BO6vxXVZzyYFrj2WrZsTbmElqvX6x9+iGVzY7+kG3
J8H8x8yR11SPlZPRtEsJ8oQoZbtTue7mtkGwWoF4PcryaIOQ20u+KpDm20qfXieT
/sOgJGqYZcGoMVNUHTsxoBrF/g5nONVbe+46D9tq2qnaQ9vJVMW/0DlI5PQwScnt
5GEU93ywmeE0HoptGYrggJrJAoEFjcDPAOzi99PjaddcKOT1A1D0IRtZ4MmerWAX
r1RMFQ4XyqxN+WmIT9QCHIfjkUWwO0qUTeHlgxVEku2prZx9nGp5wCR4Hrd+uvHy
th+yi9ghNQ6Gi516NlPd/K5J3uxE0ehR1ddXZcXw+oL+QDVgAY9YYUsuj35XmjHP
8EcijXrlI8KY3S/oAq+AYdJJ+uPva5N64tQqx4XwHwh/mR8+mjQa9GyXOPsekDJc
v+FMzCn9Nkl2020oBnr2qvvr46pSD6LJCkox94eS/cR+1RnDqkTPJMf2ev3sgw+B
p9+whuygUipyaXnt83Vm9k9Eon5Uq4HAMjtKTZFTUNhaE4Or25aivslWwDHB1wJ3
TRa67gwCh7hE1WcBSfIK3yZi5yqY1pPEt31b0Kf/GZ6i/3DrdYI8WYxbBpOilmE+
wTHYHIzgND2201Hemjo+o+piziyRfozOGQ98GAOlCeXH1e5ZLYmjo+vEqDdDOihR
661zERmr607K0R3mfEF7nbsOaCy6Fwp5B+JJq+QPgn6QoaRzWe34E42PYZKjto/k
2A6j+9IeCb1wXsbgF5ewzl5wkMKubMVkRPznsEx5BPUFEyCEWcVRu2fxkeJD4Gmf
UeAZ8dSr0LwZllfqQZkUe5D65ovvhzwhIFYKfw5iHF3emNmBN8TwHrXGi52m3HX/
2fxDmLp135skPzms62Ro7l93CKnAS4zwL1nTxChoB6eb5TtjsAzm36Mf3jyVGbGi
kwg4y236w8Y8heR3fUO+v31s8HXYsrQshh1tzYjO9jzC9LvEH46S583QTKGxgeBh
2h7qD9oIE95Io7j1nDGklaA2lxnzc50bvMhL9G3lxGmDTW3PP/tv7uOLHkBOVj4f
Po5RXzUkesmpguCG8x4R4yTqhVxr/4rx4G4lhVQ0g6oAYl0XBYMF8jTGljdlakCt
xqUbLJNV4IWNiiIhkqhVv3PpYML4NrdOc795ikxf8qrK2fv3mSYuJ57D5dCslvAc
azkfKY2hhX7T2QGEffTYuhgJvWlMyYNsF80M0uI0byJBk7CO7Z7E9lGpAIaYAl/h
+/EAEW2bPZFsZKNhsXWMd+NOsApEklK5M/sH9XT/yQWrHuOjez+rmB6L9hAhVWPk
8It3LmKYa/EkVDqamzsfYpwUVeYnoJ63j210tIaCPV1sYGXGgU72zYFbHT0YsH6F
/MMj1+72K4kzk3jERIKlMFY3tc0Z1GW0Fp028iibeNa7O0Tn80G9XiIxsJBhEOUD
imd2hShqiR2lSgv3mSF66UF97/6ABmWMFaBGKkSNLXWgdn3v6ydonivIafRBEXir
IUu30zrfBeUdudbgvvqDyOcIrFm9jA46tC4Rf8pD+EdDZBvb7jWLshamg5xhxmhV
iC+m64dzoavnsg1ZrDyTYyN1Io7y8sAASaUbZNyxJhGowyc3Wyn6GTQPaLvL3LYQ
X0RB+0KiPWh4GebYeH2RfDDDWPKLfUGb1VI9it1G//9g2uD2f0KLYclx8CuhUfLr
K4/tQUAuNcG/Q9FBZgDnkevdhueKKf4GgOK4I1BIwFuUJmS7+y6bceVQ2O6EByvS
4i/JXDelqRYeN9aRb8cfeDrzaa3xTSPjuF5KpWyiXoy2ewUVFJpFgh4rGDiaTJW4
icqQDzUw3o2HSbOg9CxW8Yve9/UNZ08seNGUMEAubgPqweOneuelw/GMojD8xk3Z
0x0Igaru3enDafImSTtQjPve9sWeEL0bQ2hBS/kiKNmsnaBz3NWgiJEQonriSeRg
thsw9Y0hnkC15R2kPB7Sg7Zd1fpopNDy0STB8Ij68OHczfFPUhN9vr4qUwN5P/iz
/1Njr1dVGVgthn7XdlEzRuA8Yba4EU5gbj1vBLiJf4SJIK+kKpbHTfGIZFtOKoHb
hylzsNS32t4fZvrwp4StsffKUJfJRL0gVcTUmIvFhQAX71wSyMWoOlTz0W6WbQve
f+BaQTMQa9CJQ/evzzcm67pKIyretM8bFZqJ83qPd1/kEqjyb1/7CbPJcyFGcqJP
ClCizOoOW1IGbGWRPCLvup8aUEnYBYdu6g0G0jCPPDVxya7mmxdj1fiSf/v5qKVw
lXtl2IJDXDntlGkH4lDjVMj/jZVzOdhkWhkykZlQxXoVBsW5FhBkXSYt89ZCbQHT
CNT/f5YEeo/3Uhx8dA9GodYqErQILK7Cpvw79mvl0GOAD0XcMC4VmtX5TRmyxLRy
nZ5x0FM7iF/87NubY5FadTOngquc0muuAXl4lj82UmsHyS5tKRUyqCdOJE+n8qar
CNFM9wwzMXrfqKmVsRpQghwpsdjY4BqesZ7YPgHV7QEzfsSZ0QqLCVdtT0rPF/Tj
ZaCeGRXgzjtFYrEK5UfSAVX9ZlWzELWqibJEeiyJK5fNLbcTJJZ0LCI/zasncf8K
IUZ8rcVVSf4Il8aOowjyJMDmFLzyqenwYJ+fq70r6no8TknE2RarJHuTSFGsW9lq
Vdo5VvnZqvPmGraK2DwUgFxYt6Ajaeh0p3el+DngO1h959kKpXb5P0sy5HSMhKHv
6RH2RS377MwP2rnJ5dyAPB05WSSZqzmWnjdw0G5Lm+K/JAppyrgPl6fTm6qjQboT
VPGyQz2YdhB2vJpsjJ7zmUeVSsZYrMdDkMjqxqGz7x0cB/389H4LWu9DoX0j4Nla
ka+rnByyL+1l8dzuigaDjQAFjsfOCqSqYBSLQiieV95Czq24bOoTwyzQ4SbombaD
19izc9SAiadcnRhKR7Un1TCKQHjHMnH5m0dGQf0sAK64LTaGECh433ePTj8bVHUP
vMlWc7VJ/+hpDg9/GBENAFfYmQvDo2N6uoRjXcyc1wWYiNgBOmvgsYt2cgDrFaCz
QrDrPLM0WV7aF+mVdxiy2RE8Fn4fok8hKKVTEU3IyqnrGTp3HjVSbwVVBtO4OZbv
Xyvn5nyvGF/jlp6RAyQloyYikEerGQdGd40aDWLpN9W64u+eqvH54lTfXP1hvN7P
NGtcasS1qVJR7D8y6L1T17sfRJpK3fIJCOmdhuqsPp7jxMFROyEFUxQEeWHmDVd4
c8J7kRA5+F+Co/GrDyC2HDL+HJDX1se5Giazao2D4GvLhOqIp1axx1oiJc9EIrZM
2LHCQlMmGe4cHwlpbX7aW+jMONFPA9CuLS1pu6PzPRunp0qOQ3iC8hhYN7z8QMx/
MY5WBb/y8EGnArChsuopc6GxCUDHpMXyfc8d9oYOBNTyGwYz3utm7DHA1vJ/IBOz
mJdC8WAK3pDfu7St4OJo1On35FvAqG6wKVO6fLEU/leNdn51DC3Skz/tdYj/B8VG
fbzXl4QUClnGJGsfwLqMZpDh8AXJ0paIeO3hqhG+YnMQspErMovoupjVx6f9g+nU
jg3panJp2iLfzNr399mO1mI9eUlIDAr8weMm6cEbKjEp7129671c8efhoAHytEPk
QHbi6ik78YitPUSDxLGHzgeMMmN1iBkFaQeoHLjahxt5EKbr3rkHFLMA8fQFDMKy
ILVHfQOUDG8i2WralrjWDBBUk+UGLiD9/0AWKiKONu+21yXo2FM3+6Cr+JpcbfVL
1e3Dzl7ZpdHEIFXlULortgNAZ/rolO65w3424CJwoCxrSG10Dl53mkqiUHKqt+jG
55vZ31O6r7SlIAJy52GOts7T6AzyLgZwKHxbFc5yMMluScEecxu9ZmDwfU/9draq
tfQcPd+Lqa6/Ojp0Z25SNVRDvUJ6lZXF5IeaA0gXLsSX88PYrYWUBjhuUNhATHzN
cjOna68oDXWnCpln00hUD9InkkUjIQNj+rAUHymmgwimdxHqMb5KTDBbmkmzPTim
4nlUKmLeyzHLFMNkI/HlHY3C/vUDxP0XVYvlr/O7zBv6T9cbrU1Y2R4GWmnCa49D
e0KPqD21HKnHiYJEVpoFCJbK1uZKrcLxaGaI9v65OSAZuy4zuajzvcds9JH7YCV+
isfnKrFyuFuNVVb6m+so8Zgzvg23C3GV5mbl+a0rSZ7mVvffpSVCWl2sOOnYE1qS
9TB6b5cMFSlWZV16y3tWtvWcAhZvxajzc2KRvvUdgxXN/wJsshDfmZsBTAUFO6yx
Le3iH0wog7W6PT9bkCOHNLmk3/JQY10d4UGVzRiAUvH0eNMoDWGI9yad2NBaqnHA
g5+0XR2r7P0f7YfPewEzmtjnLZwAqToHIIr++IH2sYNyQO8Lxo+TOUaw4iHYDS+n
2y6cGYzwhk6r7zcp3hhA+cRJ6feby+PFVlF1QSpR+mH/ofv3vQrh8vAEQQlp/gna
KHZzAuLkLFEYp8WSigYZPnUsTFP09ebur5h9l06eqbxZ1npbCGn9FCZecEhOYaYB
WJHLikwhfqi/mENLzEEILXC8JEbqJipxB2WoXvtXcki1Leom4jIw5QJ8DW1OqdAB
h9y7VBOOYTiWPr3gtgtf4w76OT9eQOdwW/j6uqGUPb6AV1C4paGZ8GGTI5rfXb7c
JSkh08DueM/U2MpEXWF+piZkZLXDVjfKuMksEfVp+yhuBlnnWMEsl6D3EjU7R5Cd
ZPL9A1IBCh8d53AEhMiCy1SqOF3PRbX0fuvpDoN2F4XjMiXXBBKG18YV6Tp0YK5p
N2A0VHY7ZrsRjQQjBRyQ5VUgBYcPaQ5go67S/Adw+s6rdF0erb4Am4Cdr3p0bkV7
ujmFG//CaipdIe3FdWwdIEBXHReRBekJVst7F/AR1iVCEA4o/dFxYA34LIK5RIi8
L8LN6OdmpefjTu7in5mu/OOcfa41PXEvO/vAIzkKXGGcZVXClAxNN7XxWIHZVzdX
fdhLejau+JuAvYrk1EBiUsgj3Ag9LPG4qBnuEeNcbBAxARbOezss4xQgw9e3WUhP
nd3GtQvkD6Oth/YnJXD3VcnGUsEdMYxLw4yldvZaBhlaHrtn0HA2V5+db0+skMrl
DbSj1LjmUmz/HT+wKrMTapip4sF46LQ04ITr2O/gSxEDmVHrvrfujE+tJhxmWH1g
qTOpIjS7BqJEdcVTGR+bcz3Xv7JRa70mYsK/RYgD9h8EfDAEiEHQZgshKI1suAK8
WQlqsysGXwgV/tV3I1xs98RqRbPWst94KD8H7wgUgeo3nZ3L7/0Nxmo1r+a862kL
xoCE6qW2zCUD6rUEs4QFJEwglX2UQUZx3tLmZGYqoVG65/7LYfXZtPbkW47h08wU
B8FMmiQhoyb+PUmbUA2Q7rkseseCr7ZPjOfHCEtVra6Fo2bsasyP//KOpADZcE/Q
xMgcH6P0jLDBk2CX1ghCKuMOIHnoitSyNdXgOkjFNpNnIg4aXLThIpt0Yim7scv1
Ii2qEhdOgRqK2GZCmYIoAksy6AAoKCuwT3ATMfooxC/kz5y3gTzTF48986Vd5Q6t
n9hxFT8FD77P0GMAkb0P3aG7DQMGDD1VyrLEUQNTubhchuWOziy1oUAgr2+ddbJc
eIB/bb+zlyjf97i16HK22ysZ+/F6nT8hbO1Gc3WtqfaVbvgDxAZADtgj43aiYgFb
KmHM74obTUvDJL4ZcOJBw4Wnwq0JpJWbXOMW9z2+lvvInXOjZcsQc65pbF3R86Vg
yUDDTamX+HsCoecGBD0DxuYUJsNan9VFxAKc8ujeLm9aKLeUpjKl1qsrGysXP2ml
L9ZPBya0xnD4G+d0p7lKyGPQ8xFi/KmvhF59Pg1HsRuUbMZldo446j5VuHoYfELy
FoTmUtLCurH8AcWES5WpKc5FrxT053GnrWHoVJn+Ka57w7X51kT6+VFIW2Zyuxom
OmJbIVjanpls4kzZwMCuUH2exUcchyrBhkjtrNR1+50w3eALCLYVF4GnJD69iX7b
YRK2BMwtwRPXkHa55osDYtMpTK6sg82FFt+sBoxQAjH2dMHl+P3b0B4PbXkEJSxA
AiNlFVe7P9rEuMGmlx7L/tXcWLjsWxRlL1XqdkeVNbBufBJ52r7MPbevF5LDLOzS
FreKiPXz29tlb/D9o3i1ty0t6Glbu6xZcUElIIvtOV951XwugAiCzQsVoqNbqUZG
siYf03qlARicoBamWySrqwnMUU4BzNI7FjTXOgVWWxC2ekpa0Z5acg8z5WhhtLlM
W2g7e0Y5gNDOQAWMPyG5xhGoHdzJjSQOECpR2OJ2YHuR36GeuAVWXw80JtOWENEq
dozYRGe0Zl/PrpHf8tHus1rYqJxmVMcbEVM0M4OuwA8UF4i+2TmJ6RN8aaeaGRpd
pl+ht2X0ySAF1Vqm3hICrLIxLn8UqUg9fDxy1tQaV+t97vrgrYM+XNuSeqlLEWut
OvMewd9YRjt8GdrT7Vmyc4CzYseLKpEHBz2hqLiYiBENXAj/XpvnyzW1MO0UmCL/
I8rZbJT4zurASVXOBlJL6jx16S7AXPcoqgOky9BB+YEjlp3eIE4foqqPbq/73B8P
wl2DsLTrMVWlJe/MLXw4iW/eUJTtiXaftZwAjFE8nls7ogpcMY6kFqKH5szHBsUR
gYGlf8b4vuR3l0ZCssFMJm6e9LaT5nPGuMyd9MJkeahVJprGDmvGOFMbA5W3AdTf
rN9DBHlWktbXAQLGoIjUflCrdcX20hchiO8FRZ8+kv/BFB83WMj+nOQvlCpGAjOa
lRoLlmPes7aWTh8ZwmhNEz9EqmMIFWoGqYtPPn2ATzrR7d93hbtpEJRVC0X2SFoX
3Xt0rvQwAl9OBf5/s3TcQE8tXMWKY5sJ/vEMm/HuIl7ITL5rYpgD08blDXE04xD/
7ch2xA7jrI6rjZHlvL6Rwkqp9Tf5z0AYF2NpzQaNAeRt3QIYy+joWkezp6g/N8iE
kWWtQmoWnc+NJL9XbKV+9cuCJXbhxYwuli7PJEiNtUAqXYQU82Q5sytVQkxT5UiY
p8VkNv18golfcKkKPP9z0VQbAhqPGUvL2S9GT6J0syBIfsW2yD/HNA2lSxP6hGCx
IOJSWGIQTtLaJ5kH59OfGCj/4g6/YsfSiInPkfqVDJnPVUI3IVYXaCvhTwHocYBS
2Dh9IOzXNmCCWJNllkgQhHCqtkYKpZwy602a9CST0O1PQCmsslY/QvVBgerQnufL
JsOk//7rIaS8dkdmU78URzrgndLKzY2Ck1zcRpR4pZD7Z/h9NWHTU2k56hixhbKW
ezlH+fA9BgXvWp3ItbSXsluzluZGdPFClc8YLZx9tyh1rkNq3DRi3YvgG7tY8oB+
Ry9HyVCgprfXLcN68xA8JE+PKahF9Y8SgSVa1+/g8k49xoiBpCpIf5JbnD9Sb+z3
oCFEbYNQb4j++g09LHgXRXkx1XqfaALxu09ThMny1EqZBBxaAcb4vY8vzGdx9t2S
MAltRg1zzUvU+B8pLm+hrTUxpJvQcOhT9cR+GmHMrzA5yMYGNV/2IIiPj9x/bvro
+Qo12y47700oYBW1NdBobWiU8mdwylXwZ9ZSM2OPKSpZq4UmRZbh7iIBbTollNAO
dgQAIre7o+gHxt5Tj+KYHYkycZAYHweGQbcjei1ko1yah3H9nrlHmE3baJhQhtN2
51D1dKkWginkO2WLp1THMqvRC6W4QHRIGwVgeauW3aNASIWkhFjNOPXEAa9GgXy2
ybWih4n9HZxkTOi7WVIeeH2DZNxe/BlEvhWO0OEuuRoIjG48fzOSumdszY4FFbaw
SiQp9Lqw0HUEx4fhjOzcQR2g+b0vh0M3yKFmZmArJYyfSeOLVlXT4Rx0QbYwzd8T
8JaOEkPzeQ5tku4xNux+fWyqk8b8Ab6jGQGiaS2MKYgiAFJTZwtO3cGCsnrRZcgU
Kk4N9K10Ig3zhUMUXAIeuWFCV66Anz8zJyajHDzKqF2zc6vT5Ba9wI7wm5CaHy49
bHvaxfez3Ls4QuCtOqF4IqMW5WB6uWLRFur46pZN6mjuO+b4wryTfC8fA5v0QHsI
ChNopQ2oQhNFr3JhW5haHhVxnk3xMWJg7xb7GKbQ74BilDZr9g0Fq8i/RfTv0kxS
MTub53GvZMHx+rTDBKOhgtnOF80uynBBUXyPzw7K6NKi9X/74sD/7zBqUPqXj+jn
dsuEyrN78f9zIonvvU0uONFuszXp6vL5qEwHOQcPcjnOVgBMk/c/LUs0hU04VLR9
ZPRBMytSVpUdqxQI1eza6bevZ6N1K69lKbnlOc+ylaBz8gzRjqmt+d12farie8zH
Y7xgHRbE8wzaumF3k3Cap5lTDAT1KY22rjLN2YfWsrE/lH3pth4HU0YTdoX+Kc3o
3CD0uOjrzqKEFw6u324H9qB5ZpGmoLkQmVroc2EbgAuNPkeYK79YGSSuFhnisNCy
0g0gZCgD6nJUMgv/8dPby0Y32Bou2/STMKJlf+rxVWjP3DDXxoF/XL81xKNG7p+v
7DTe3y6PrBmkCgZrdzzj2AYomUGPErNYNAsqjrbPPMBA04EXN+7UNWYoFl1edf4d
V0ouaZu3BJFx3Y9gF59/JlIXcZEv/BViWCP7f5+IsXYmOlxeV/BcCRRfA/oh6KJO
2IUCE1RsQ4LjOoLV8ocXP8Rgt5Cc6KKj7rUhX1jE3Q0sgFsYMdYXSgp/QLrS8rhz
oEcu+ewSGAowFPQXWyMmq42AthYK+8squdKf3tSJPbUKd7R1EozsyiyYwua4Wib1
TsIxWO0mHpERDauoz45bK48zAo0HMvUnZNln6mwcL4FLWbpW6GhrJDerc+eQgLoM
ZRLvQViMJiYTpXyHWXxKWpUNICplQAGZvH/f06v/eLId2luTqDL9fA5682HhEipT
Oc47fxpYwnnNkTtUc27xJgl7Cvzqfv3r0PnqDytxzXjZha8PZuhbx8dtQhK+BCZ/
QGPsHNWp5GW7quF36FlwqaZEtYusY3TTiTQp7qzzRkWEiEYlrmw4o2hg8O9Kso6a
gIeNNkFu/dwZcCJmVZCTCTMEgkp65FwcGky2f5d7k3FG+zQhc490djYG1cEd+pmy
tCpbezBbi9Na4lmXob+2d/BGGWBwiedsGBVwvXDVAxapJtRikHcziHucZcPlY/Lr
XkP4lTJrhewSzNQnzK2lB5pgJ8RPtle/i3gRhaplu0sNfHU7hUE3H/q2vu1W1Nq5
plF6WbZEz0PCjRwhy8/VYDa5iIjVLVOpmvD5sRiOhjFHkj0V2/pCwVuk3VHFco6j
EVzEb1mo5UOiW4Rm0ANx0IditNPDPoRPt9gGMf1Df5soxWk2Yxr49Fx+m9mJ+t8w
EJAtF1jeUXvurJrc93CHPMCHPWNk7sAWCAOP3DMr65503SnvwzKQmy+q2hKzo3yV
2MqhgyOrx1Sau+dJPvgcfqGNiuuayWZX2fQanCkTulLchETg3bsiIXCFMTmETzPp
DMaT7aZB1+8fViKJzQV9raIpodYfQ5GTdU0QTrpQgwo/HDZXjtJlfxHJgRNdjni4
X0mY3kxm47i3Qe0pJCLXlRScWvhSHOMg096l+raFo2ynXl1XndmcnEp8KWo631il
48KWLM7D04kfkl8m+E+YPtlyzMltLvpQtuiB53S+aSYRFG9u5Am2fEblpQ2GOFxv
LmGHSq9r/J1zSkH6uuW4ZQE7nqBgs+ulo4S3p7FBfPoT4BuL+MHoOyl3XlV/yU8P
pwT0j0WiGrZWI3ZWchzvIcTbDSF+/riSfHJjCLEQ6HVeAjJoMIJ0qnGfIUFHuqKd
iEvPiNyBk2SS9AXEHiXjI/U4+ZGTsj2NwXeLWNa02SMgbNgTRS2+X2AUBhh/IvZV
etJtV/RNk4Km/jPNkV0YlVyl7pwao0+YYg4wSWdhY+YcmbhAwUDbrIrGnJGTElHH
7h4ARIGcg0Ln0MX7QYYKyN7pwfEpBbz9kwAJ5mlDoVLutGYwhCpNy/k+yl/lK8Rb
/fdMRIS4k5ir2F8JRwDj3fpZ8zRZ9Cj/b1vTyhDSz3Z0vhFL+3qpTf/4Qr5A8RhN
qgEJvwF7ypCML9lZWuf158hJI0ui2ILwEAdG5ohnZwOvWvyAsoF0U5yl46N7G7Hq
I6DbcrbwaG5seXfEmRbkPfxbetAWRGyrMlpzKBDnA147FVJ8CLrj8uVXCh4mzHMw
8Qtcm0sXK/u93sxd2CU9wUjdadFiAby4HsYYXFyzESnel5itF+tgYwsp39t+JcG1
xCQXrd9L1MpFrj+RA07E6WC8lB6eZKDabdcRLbgXjTG2tDJYw912F1zeSn7ArUvP
xcDembR9/l6JRmkGPv6J/NVHQSlvnbh09VJt8yt2YKHdmVqWKlL6btuX+0gZRIad
xYoKzEQP9qJ7uiX2yrK79ZYWhmNSAa8PGKnKX/BE+Kap1tASEqty7HGxX317AU2l
GodzbspgggqdlbKIEUm5dyuKaEx5YZRuTGrlYZqFLDFvORgBHaKGiJK2wO/iQrNh
qMiXJpZIkDeyRLlNx1twCIIF2GhfB8DJoB3HrAxX6Esk4fdhfHQnjCJZRKA9Ux0/
h3lg5Hep2x8fqxtnG2uu/oPoJn81AFS7wtb7UsitF20CfflKuTt+1qlRVuixgTeq
c9QH0fGW8NKYVW1WMDSVRBRtupDOnTirkeNM1m5WH8lutVIdApFfsq+F8p39Lz3e
yXK3N0X/fscMApigfy7wrbyrD1H6VR+19SCa60yOij8E8D3/VdAusUzF79l/RoBZ
LOROfHF9toUxn9WamujedsGwj3BpPhcZZ2BAlV8BHnq9MAmFlDYPHJj+o09s+qSj
lTCYFFGoEB+/a9PqDZGbZ6KIkcrnR8m9LZH28ZiKZA3BK4ivp7kjdpQZmA5mREsl
h8bCmPVffscq1D1X7GNbZ+X5wJxA1vsUulN0f39brqgFcv/6uRPfP650xH8g6kWV
29steqjsEsgNP3fEEymMG7QqNPJdqsRYGJ9ae3jvUmljzdDGQmam6QnUS55vNY3g
8yjfW5Nan8rqLQ0Z574SP9mKC7ZEGeiNIzkL+FZsI4iqDrml5eL6+Ti/U7hRFmhc
QC+DpU0Uibt7jPUVjpIrS7BFx28oL5c5Zf47cSfZqtf3xs3ZaRbcsCGIKjoGMQle
MnfFVUC8OQmaiTg+Dztf4HZqaF7qttdZ3/Wza8hZNwwsuuQ35dfkKOJCcKfecRXO
wOw9nxo7+LMAQuSh2Jb3oe648lZKMHOyzIuMg85+HpEzTYuLBKby2Gnqs3sbluV3
1PNFyeTTupgcpc65loNTYAOIUtuZuXnmQEylakJ1PAkccVdh1/zfHr7vHCO/VNjK
H5mIeo15p+gl/6/hCEW8x2G3TU6ljZ2zzCxP8vWIr0X/dOT/a+T11lZSIn6OPsFr
SNmkE9ZZyQqzi8tshKMYDu3O7GBCGThnB/gouW4Eqx0K9kXQRz0H2sqKd21MhRRe
+hTuhyokaX/hYacdOpagLZIb4vNg0izGXl0HhRkNPm4tH5IBKjLDODMBhZYn7/7y
31KLzbhUn2lK/jXPmsyL5p6hm3RH5eTJ9s425/fubXXa0ndGEqTYC5k3wzK1pNMT
hJ2s3uD6jx47i+RJDfEAYJd+rDYpXIHZKfVOVpkOvUjDnZu7qABWWnW2xXTbvmqM
wGbnXKnr42gbqB2aZ8hAHQoQEBN5BCsGp2VTucYWRO5yPEOZ4u1O6s7ij8prbf8l
P4yXjr9zF3FLsm8KZ9kjR9tkrFlxBM9n/eLaQ/WbOrdZl6laWajhjBTuLmAD+y4i
AMSohJxacv6nFnbnpGxeheP+UmIS5/c5rFE6HaIFO7GkVBsqKCCvFEEwP/aGVqma
OHXmdgLi64AxwkNdQFoiNqjCP88b5prHdZIM30dJulwfCcdNnwg+h5HH+6In5lbd
w6Poz8Z9Dpys2vF7zEOdxs+YkxeLFusDmllfpfnL62P0VfqIPneRSO13zfOKdRKb
2tPW6av2syjphwsAgoLKvsAAcYmrddDtJFHHVU1zTHZpeLXMVFHwt/L0zkdi5BdL
NqCPYduTwZdxqHzyXF2DWVPhJwp80rea1wpskA2oivggXDrj9XHaNIDbq13gyBCH
QVZzJkCCsM75CnVK5IGYDH/S7NLN5Lq+g/NqWpv0UvuiUMUciTCdzQHZWMSsOyd3
XLNpaDqIg9kVnJJiBvHWLIQzBb0vgQ7n3jFy8AKHwZVQLiPAg+wJuDspcnzyt5Kv
+YeB5v+rwsInLx8LlVcqJZ6snWLUBnxpVyfQPNgqiN8raYl7x3RnompV/FrY1B5M
MIpQps/FmyuCeie3QRmkt3TazzOul4CrEHdYgCAfJcTd8diO7Jap2VxmiUj+8tXL
kc+bP+6LYd+CwZZjn6iYlIdeBEzRFHZ0RSqJ/XsDuL0z70lShiRBZ0LE9vEtzhc8
q4w7X5yLEKOs2DzI/JQmg75MO+Iupyl4j17sUyQ+cu0MtR8CYDWf/0uzTJQGqjCF
y1EQs8bVe5d1saGNvWsJ96ZDCU5PjcrncYekNH6otRR+0RJ3gpkEhhXGtrqRG6yV
9QB/Oq3tu2XFk+JPPMdeux2reRPC/pYGeG6Ls76yDZlGmyn0i4Fws93NqRkKRs+m
saMQfau2VDo7Y+gC4zTK7IW7iFqQKPjMMLXJXh2L5qu2v8dEwmXPgoB7v3HTDt8O
B+PJrpKF67Uq3Cqsw/LsfpgJ0hw1ynrwMQvgb4ExtgwBopS7/9ypnIFoSA3YX+rs
vYJN7gkzxd+gZ04SohcU0yFuOWxtquQoeldEmZmZlmE4ylQoYqA3GdC4XluY7uZa
UlgiS1hrO5Y9tTCI/vlOnPn6XFmE52TYy+T1zIcKpnRc6DVAS6wahOXhxYSkOLjY
a3OTpjuvELJlZDOqdF2eD+Ja7CNDXiUi3+9YEP335U28zoHTmpI5r45gUVoTZ3wU
4zDT3o/XX6BFphMAWykXX8inNMKmuN9N0y9BsUwrDFxHxcv7AlXmsA+LLhPrqsre
5/ef2tFbgykfnPIqVN8qi0FgRMHn4KMlxfh9Ex34cx2cxXvwepPVkEKukE9R3fd4
8CjptL84rRKattqd68fUdxCwAGFDhxKHi40iflj418tKJeU2Crb2KTwVS5RTi2xP
S3rtmSDobVGemkPjPLNkhBPu1E0njNjKaXOU0plYheuqaiXWF4Igur7KS1eD3/Vv
7LRV+CGyXKAbh4RSz1OV5t3wk/Ell77CLndEyguUwjTeWFxjJ9AhixHJaX6XvOY9
XvO4RTqKgGhRPlHrLzk4DC4Lepsnw9gdA63Ibxb+amtY/pseKfUMDidk3AxcYxnX
qpDJT380pTG/VwuvRJXsQDjp9UdnCE+o+1daj5qiZypQ4SC2n62E2TSe0SeRfUgV
mT8OFkMsUamRc/nD4zPiEcRFc74XtPzW2OIJmQwRXZqPD1PLcimzzm7qZsihOAnV
8GGRzzX3vuvAzyWKKc7QaryKmxs6NLmXt3PEJfPZ0rPsiWaq7exyfk93Ygl0sy95
ptqGJxcZhe5Tq7yEogb3VDgbcKwYJcz2zd323UY0fxHj9GOqsDQb0HhVfjE9/Paq
/s+aytG1UsWbvKXr4/JsO6o38X28hLXRjAccwqCvmivHLqKs3a8XBnjqzabqjQUd
9t2z62vEs4ONq+m0g1DDveoN1hbvLxZD2/nE89Us5yrkNN4wiYtFhLX+tHQXu1vU
MxMKcPdUO1S0K154sm4hnOWsBPE36ZFKYbgDeQlIMqy+2zwkTTUjxnNT8XQE50S0
YgvAjTVzsPWKVakpoEMwPQBQTkiN/WijERqv1Sil0GCKb9HQZ8LXU9iv2WX2XRzv
+2+046LmzrgJeKJaW7ZaVzwmJ6ALPYSA/45DWAGnODRpM+Gqcgl5zvIWsMx1QzFT
H5V/J2YLAMVdUIrIbwTZCDYSvjvsXxpvxruj3p+fn+8hIzayIAk8MPxa1OWOpvSO
YWbiyYbrDmuxW8FsYyDcRnGk7gZVCG8NzTILY5QF0X1QlY5JeCBbg06g5ANJfWSX
PcS672z3eJzqEg8grtjPwNRMDBFcq5UdhbI1ibypJ02ClDp6EUkfrHt2p2b786he
/BTl+nkeJ4dfgNtsSqbifwo8nRm1t8m1gW7uT3QzvuGF22QalcYrUDm7PG4JYbfC
auPlYTjRMYUyWPcoLsO6QmjkgvnOID0QhmJXsGjyJbEvK2tZZc3XW5SYMInZ0lOa
OClvohAtA0W4PYdvU4qS8xfcfGIW+DhEPLjYhmR8HG1YcoVNtJVdYrJalVfbSC31
DBcO++bdNiDIELE+cObMQmNhyMpXi9fx0O1i4dw+pX7qHTh+HUa9uAWOz0BHinq6
l0mEjjB73x3u4F62V21vWeqEBZyEMciCsQk8tQrW7vfWBHEDLFLsCm8vHNAcRx35
FZ3rUQF+YTOch7GUbTyJV026gf0d6lR7K1rajLGAY6u2WXWvldAT2PcQ0R94V1d+
wqw6h9CVLSELr837YYFbuTJlZiU3UBazOirowT7ZAf+Xtcej7D3JaAVsqu1gSWBv
oVvVNI+OaaeCSFGVV0lHGRmnM5V/Nga4HW1mEC/an5vZMYPScxW5Ez+2LQsVa95r
JHcuCDpOLYYKxH31z3X9aWiZZiLS63D4UH2bIb9dzwcBX0xaT7b4bYkvx7Cb6O3P
844PipTrhDKNGQjZGfdGTR+pjTBZoEbmmq/kGJzxh1/MVRDwNo/6IFigbvKup7sp
iqW6ImMHrjJOZAgNCfQYRrHloSxkDGQmq2U5DHm/HYM9nPjhefOoD7c/IxbbrQEl
TJN5ichYTHZo4QVQ+4LoMxfBcmk2fL/bH+YbE/ycIt/Cat0+k+Kxd9fK0N39akWT
3qa+Dd1kl9IrK+cuNPIiXtIRauWBYSyNG0eFkb4VTHUsATqpy1UwKAr9SaulM1ZX
xd2tU9X9MnjB6oQAsNYbF9E+w3unjhdqhEw3pldF+5n6mbNMB+RIDnqrXBycug8+
T7io4GbdK0D4irqF6mCzMMW2zfsoFOkLwo14yZ8XlHxCDNufZub8YA0R3KuU8+0F
60krfnP6sjAuNxmNc1G99/vdbwGj69zDtxwrhu3SeE902kHZXUamY2WmgK4aywpC
YiNleb5txFH7wap+EisAzfwtc6D3r+vcq4FOsKe900BPpYLpJyeSlU3hudAx8WsE
VKJbBeHVPUVoh0f1I73tAm7iWaaLhMtwhjmmQdOlSUQfUGv2PuU4agFvoF1bkWDZ
oeXNmqWFvu6mMKrGN/BmhfUTaTMLnzk7Yj7hRHMDvJk7VehwiwmmRrkY8dtpfCVK
vpvVsJPTzDKCsWvdmbsBqBFyD3kvPJoIB74KmhyPXVFHzvDXhv41bmGK8Jmsfy9G
DAdnlge7A2MeKj1ho3Ca4gSEyQzNgdL9JU65MCswywh+WUHDe2wDpEzlFhopfVKS
vCFf/HJayYtnL9x1Bl4NKkBgXCAPKMJgtyqQwBwa2gfDTRD1k2aERCnUE5ZTML6Z
d7t8MG5pd65RfvLet8nZbKSkW8KwsGm2jeLiHhStCt4NwSmWGyuY3m/x3eqE+zgo
yd4vh3eZB0g3mMO4ERvhXbo1L5lcECW885DcLlwPwpOiSdxgDn++fh4g3HpBJyKR
0Y2FW+Ryuy8ghp60Ggpbn97NMXx7kyZQ4G2KKtvX76cRfruSmWdt5xKy2ME6+EAQ
YIwpc//g1ctjnQ4abBtbdB3PRB7CPVWXklk6OrkN2H2ITqkb0B4LmiRgFDjbz5YV
hbRdEnNQajoYsM1yuP98KUziZuZeCjwj3Nl4R0CSLljAPbjobrr51sL68bKGJlDf
3Vgz132mcsW/P77OsIzCv6iXNq5CZgGkXtkOkTK789ym/o0OQdctwqAyO7A/9tSb
w4w5zJK0FVXH4LlmpTZ4q8QEmq+FqDbMcq3f8G4bq7SUuHhlzmxtz1dELDbyowkX
omorbV6F0X9JsiX/SKD8L7dKXKKeHJ4g39+IiPc10IBk2+y7CHIbwLw18JJ7C3kL
gm/3lKQyK2D2xnjI6O6O1MOB/vMC/9HQooH3ihdSPqqQ6ZtICzDqGYl6X9iKkzFQ
yncQZb6XnHEnmHWx8644DPud/rAG92+OssCVw5MixsPuO32Nf8pnySB52Zetqc3D
a7qbOgPd/kU5I5+aoaZNuZVtwC23TMy7wpaSEqEh/qFTLXgredKyLxyintwGmJGf
019D+qyFaH2bzPqkRDvwh5uGepPznWYMz04jVg+ltCpzqxQ/wXrBci1TSknWDzUo
fmy2hOHgEsMmdJprDgLEIk8BCWiNqye3uNbrSxavcLAN7G0l9cG9EXw0zeBQx82s
o4s+YNTGATTpUbSMzhBkCGG8qqa4+7wyfFS3JDImfHutfTQm2fhCoqHwgiiBO/Sq
tzNbXFVejh7JsM8FXaAoIH0QKXQZ0kutNK/iYellvFkgrjXKpUM8ukwJS/oxKhWe
av9AU49gUF4PwSgwUlwyWMC7y91xgf5pnzpHxcXKmoKeWm6fFwl0iaqPxumj5tlp
eIBj31mttN+S7MPAqZzzrJksd2XeOE41asVbJ+oGjj2O5DcV4/rw+OZRt0O9RxzX
50W6OMQ0h3KdLXFCPk02rXF4S6UxZiZUdYlL5K1JnqVnv8mdQxPSN2QwKK2tg5Hm
PZCz0hfCLFSc/lJZOSjl/qtxQIkReG3ofgRdN4MXmE+IQEOl0XKmTCSip0AsP3v9
HT11g6TGtQZIL0TmQIENpsMkAzK10LBYWyyrwS2zIV0S7b+9nPq1qgJAbLwq7S0v
LEVLRDVKzrhKoi39wFO28NOZBYO4SNfEx9pbY1nH24UOOCR2UzEEiO+H3noIo0lZ
XMuBV81PbEheRuhO3P9vvWeOwDtzALI0mFWRCsQd8POv3OWRgxqhPXFjgtKiwohq
ZDsdH3TboQyC0ZqX+NXmi9njwaPgbXCr03cuQgCyP5dZTq37/AfZScm+fEO+nnRg
Kb3CVZjrpyxNWojT0rBNoADEK2JtX+FuclFY/DGf8yn4hK4vLXnUxqdAR6mETnOc
1ht3RwTSpj6bIqGDUlt0lx+/938gftV500/HIGHXfraQCpKYsbLPnI0tyfujl0lM
5EPh47ekcz04oy4KQ+k+oXKchK/jn+v2mLTRhmX8KbLIQZyD4cVleegVvZFrlunc
r2+BVJL6J1rYAq8sXx+uYT3KmoaKmcEptfRs3SeHP3xmwDDUhWhCiRVIjPDOtot6
qajmcrHzVAKt3CLzSjyse8KScfomtN+DMFPC3CeFQ3A/UskAuNOdwgHqMaIfNl1k
3ZHxMm/ztuWeAaOGceEuH283PSHF7EUH6AZC15UEiBoezAoPUNtuy1pIn8Yutfyh
1n9YVsnEBTNr4kD2Wb5/iBbLL9bFreu3qLJ6SIPz6RnodljjUpz6Z3X1DoyFC9g5
jH59+4GetR7SvG7Ei4qn7/T8UKSAF/TBBkDbhZROgCClgq6ptCo+5IodhCsvLD4W
3bs7x78BhpyBH9XEPE99VAh8CdiaVzRQ8MdeMEuSwoZIJIvaQr7k75FDV8j+K5ug
BBE0mgkrJlCCoquyMZUQFOTr9d/Uxs7Ufyp+hs3Az4XyLaCv1vH6iSqID31srqqB
urCdSEE0mCi++KER9ONyuh/JBY0og47cOCzalU5DmUtgGua2VM7uK3G3gQUWCYDQ
oZNGbAichpKX916Patc9AkFrH3I/5nEGx9leDaDzOQeVeqNCOpyS6a+XPWG2+86G
iDMJ0AKpTCF2ipgDCQsUJLjr+ewd0uJelVH7DoKal/3lTrrHI/ssW7RTiGmiGVJL
5QXLinQtcGCIb30mLHuMH2XFvFMO78/mQXZgbJzQ0jeHbT78aS6MZ5B+5rafxhRD
42sZGI/v8ybVE3fumNHxq6gGWDkXalc49m4kTtQ55tggx/3+vT4nHpAG4j03tLlb
odS4ITFHwKFtm0sTLmi1UYmgRx58WvlHecfvo5QoZ73UYU9NyktkiDzmv4jFlDBf
ifExIrgciyRXuZblDrSFN4ktvPDEYpNti5DPXDJgYtpzgOuVzDGAY7poe02rrq1i
MaaZXqijkVa9jH31313qpYpd7iuLlw4OAX7sJI9KJFfyo/lwpp/MZx7+GrYyTGMs
O3w62PVdNEQcXr4FTLR0/cctlCQ0LuASnMP6Cy10y+sHzH0T6cPU6p93D+l1vjbQ
UO2r9CfQJye8VlUcC8mNvy5s+xWs5tmqSj5jntyRnajqZjQqEHQYlgJs80Cjf8+Q
QRGZ+zCvbTRmfo4iWSyB71XS0w1MzgypYtXPOyHiXeokBkrgUKDBPFivEL9dYlxA
OKiu8UtMmKZmNlcElhQFqf8msiFsppiXwokwxa49qGw95XEaBOzFNV5584lE/ZN+
K5V+wiXWlrpFqmekOcMOufSy3yoEdocSuBW2AaFI5i5ShZ2SrnfVudUqvAeh7Htr
DRdO9Okz7Ho4lqzdg889gS9Qp6g4+nEFsWV/gStcL6TxHpUWWh1ayomGbEllIj3h
FZqIlQaZn+jktlSxnYetBX/eI5+42US7jZpS9e0Yqlc6/rt+f064enuKYmF75bTS
h+tAh4QfJEUaYv13wAWjNmo9mmB/wSXpSQ9b7hFNxCVgbghq8hOAbWK6k4BFc1CA
N5CZS8FVHBpQ54cePpWNgfNUsbn1FATDfyyZRM5O4bXe68dOkhVcQVZ8NCE/jO1x
lnXw3xxQVUO/0ak0FbcNrNVQpijeulAKoSlEw+hbbsk15as1AtJoN+za8DWTKwjL
6TSoomJ+tFGo2iWOpN5B0GfkQq7M/uRkowHz8T6UIq/tf+D9w9+Qk4lMsKhilovl
OLOm7iVfjaEaoSN3JhraRZZBnD6fikTkc9Tnwj69R9c=
`pragma protect end_protected
