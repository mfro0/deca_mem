// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GLzTEAB+RE5bCIVK8p+Gc0MWeedNRI3bM6WdUUGHSBbBAtDxhM8RY5co3XziHq1i
HASMypoiXV0Ja7fEkyC2SmsOoyz3sp3KMMk5tUXwkZ/zaHcPdihYLldrKguS6dqb
4BLQVT1pe43VqH2VOQbvPOQtbN2Ri6nx4hCC3OvQVK7aRApJ7JUvgA==
//pragma protect end_key_block
//pragma protect digest_block
onfnYZkFAEKh95/UsLX4KhP/iUg=
//pragma protect end_digest_block
//pragma protect data_block
wUX+YOxt/13NWpQKLH/DBtypCBaxvmOAuxgrab/tFGALqitJqehjKT2kQZCuljWa
qepXA3eJnu/sAaRnDv9DZuemFwWUm3ARaFsijSPs3hr+ACYpJ27rUFfxmKnZi5qS
Q8QuV+eT65Ix4n+K0yHuY6JqicrH25tCcIPR1G8QcgVQeDmphqxsJYbN5wm28zwf
8Zr2TmPWRAPolBDEdnt+ACly9Di2XLCv3M9zhKIQqWWjMiuKNuAAqHei277xhCW7
o9c7tovBAlGZBy/8v/T6L14ZBqQ3cIHYTQQbaakPbqz+zH8zIXQEYHrebjKEZtzT
6KE/l1YQ7a8IRAD2nJORfW2pJtdP9mn+GGeT8DMLTR5NQF/2jQmxsKgjP/tuU7gX
rxrR6a6wjwo0JmT01Y0aq2mErx4x+4xxxeMR24pigEErsA0ytQpiKs73JyGFSPc4
mBNKg6XBUjMm6jUqXI0rxY8xoxGfa3679TVTIGOAf/vSBI+Yxqd35TPDksWLLRpR
xdtGBZgvB1iHvnH+VtiNNqbJ5jeOn9dQVDc1NNlwABZc+ZDRs1IuHlDaGFF7UZuA
BpzJYDrosbAa4jqLP0nnwykFLHPZH8JbrLTWJhMD3opHaG/mGVEH/31wResE0IXb
LRA05mMNIUBl6ZMdF5oWET/OXHYRgObdJmmf8bwruzvwHfTaUOG3qNi0m0+amr8i
TaDy77i9a9VUFWcUtUlVfwLRwv1UDrsjELXa5zDO+nRIFj3SEM4M8DAj4z7MZ2ov
IezYBQ0jsqn9KwZHcse69/TsSk0kqnKfw1SD59BetSOhRUJ6z/omXPWCI5ZMeVsh
m46lAuUgwe9E617S5GTrPvGzNT2CCE+/xLjDIQqcCdPwCDUI+FOuGvN4zyOpIonq
IG+G4jx4KjsEN3HU6OT2PJYiSvCDCAbtSEcjGvouVlzJLStpi6CHp0PZGMoFYrH1
yO9C67B6Fhk+8S04h1/fKp6Z6HxQuQMhGn+jcbhFeaDcvVh082z+iJQ2eQkpRIUy
10UAc7LhuNdMRk7FaeQt0zCtxDcFD64FTMPipX+xv8NaPZV7gh5Ik4SEU+hn611a
9apf3V9DiBJlnT5GlfEAzIJKX79dG7qjlj0vgnNgAldUdFahQLY7+107iS3OwSHf
PY2VdOzS/Za7FYsAX4jNRXsNf5gH3UsrVdSGJIr9+Fr4t3jqy4XoLJMcSh4P7Lux
zsAgTSX32moqrfw4WUj7tUIHzqlVnuuJ3k8hrWYDUBn+WWJv9AOe4S9/HkGgBcMJ
2sdmh2ivtRqiYBYsvLwovfvG+rBNxHFjnHtBQ4ywzR1x3n/md/5rf5AjvOcohl7K
2OLgjqO9knzYb9OvjGXdKq9S72TyQaWh5Ip8z7gSlkMh0VP5pFciYJQmMsOI3Oof
FNIYjiPSvQwupmN17PaF94wjwA4ya0o10UNF4LgQd+AHY0me1MA4cM1D+mGaSl+k
bpmZtxv/S+mXO/ZYTS3p5Wla5LHT0DaRL2U+ByY361bacW2XiZdCeeKVfp6jCSa+
5QCXXxa2EKQUKEiSBCvmG1MfF46iV1boQAAu495NVuUwyozXptj+GvScC50+t4tt
DuvZ9niM43XAQpWxwolOCykGqOgvK8h+sJFLbixxe9KiHhfn55qDM6rCI/M+/H3B
fGYO5H6FoxqXWfTmN0pBrEPqi9RR4QbNkzW27yK4GePuBsWiw8k1I15OVac3/s4M
C9kbcWH/7ruGqr/F/lEg3Tks6CRQEmd6RruPAWzn/iHZfH0blr6nMmjyDBbDHoKN
cbOHr/3j9jzBGHpSk3XvrgLPdM4EVuDREdv+rIos0+a4VYcXnbzXNW8ixK9sITW6
bJNNQc56i5z2ZV4Zghb30ga2EE5X8SqJACYY46lDxYW6oIESDxiQLV12C87L6KGF
VqjZtGc08wy4h3Wzs4sv9mXC2GpzZLvZvBUIjPf97hnRNvCGGeMEMXsDnOas9RrZ
ICuxoFEQFoLThsP3GZAQPD+KAYVeHMB1iw16OCi/8t1/ACtQ941qWlCl6z6Ydly1
weuc0hsUb4p4F4LzAtoBSzu3/FybMHdxtKa916YoDncMj4U2YMSAQgQ+AqUFuNdy
VeXlhQwzl/k53kmFSixAp9xD1GuiRiQvlh8MJsJm6Y4720c6UmPKNURdDqu6Wmzv
RSXY3za0yzp47W5AJb9xcBcj5q15UzInuqC8ytnJ7lQ61Z8e7MOVXjEDlw9aMep9
+m1HeZls4CgAH4jtEpE1PKqyDaM0wAqRVosnC4wMPkarnr410jN0ZWksRjXJQkRJ
bxrHQStv7cXZbVfEFckxw3RptQ6BqqWMGxTeHGWeqExCZuZ2+DR74MBpwt/CxFEH
oTT180TvvWtfMYxev/gDaR9Zm2W/gh4WTMFDIB1tPcX5UmPOXgelh/H4Wzma7T3D
nDtNSdcOz9eYOxlRhWLa07fdPvdRIFI+lKEfmswV/fB5GwSU079JGL4vxgbOYqhr
vLPX5WCMnzF400rLxKQewhblaqkyqRGWajhFd0Ht+W8nLKoE02ZcsHPdKX97gXxF
WD5a+4hYWlcd6K7+B8f4TU6Ng/uEo9tZ4Eo9BYtkqnGZLbOHeUK5T14v3i2k9fF+
lcbY/3v3EFdK+0B5QXJRDspRh2uft/6G43Lz8IhLRZsinbyhLIdHUGL8+hv8ZLq2
VI3ct8DvOypVehP372TVE2h/Bxi9kjhCuC9mhLBwd13dYDx3Mv1nvOInQPUkU/pF
nNBS/FwlloIa04a0D9M/pxTvTV6r+BIP7qIs4TIXC9Jg/lVIq6RYf/zTMPZ3tZDb
f2XjGa47uAn5mZHQ6kf0St0ljbvrU05JybG3U9TjDvTbBaZVVg3ZWhrnndMoZqkc
d1VaNMeCRNRXY4jQkE9P6S+41fI4undCSYAO1GO+H4GRiI/Z1fdsyBBOK4l4a+wI
OOM52o+4lXsuqEtbOVye4FRLdhYY9AHlenYyASdIexhyfp5R0qXdBIh6Q3dXrLA2
1T71hnTAmu1TO290+DbCIiUTP5k3PDNW1zu54hfBnOqQjAmG0M4Fn0UH+vOQtPwx
8sqf0YTvWWsNtIRGmGG0q5Hbj0gQK7IXi9Ajig8CSqJHXcS9aMbKOrA5kiKAy5zq
BaFeSE1DwpisnColZph1OwDv9oH+sL+s154wt1Mm3A7GnAhmqwryTR8DNj9TNaqd
VT0dQaIg0+yRmJYwPaYqTqRRwa0HoBZlXvbzARf5kJURx0mdsVrm+QcXJPrsWnXS
6mwJzgu4E0JTx/2STLlCo/Tk2eYrvW0WhWFMzNL2iUaGcCZMoSrSfh6UP9HhGBeZ
iJmiXnpeOr+dvC/7bYJeRJEsAVv1bXVtyLNa7UMkM8uRVykBh3baYHobAi0aWVb6
9JODMTGManhBNsz4YxHp7J9KZxVrNb9Re+96lWgV8MJ8hA43FTD2M10+4bCAs2og
JucVnd6cuq400X45WZC7rfGBv4sF/T4REv9OzRvMMtTxphamW81RFQ2DyngSSqs1
tMbyKQbdaIPT131O64a2Do0RHjDws5H1A7iFwad3v90n8t241G0d0yqXGO/kaFTM
Z2C24x6nBGZE4BzQVBfM0TqP8BlhlymzFKrdFn92SkyuUX6f4KoZRcSxHLVMDRnE
EBtke/Dccs05habNhHPiCTWyMEu9fVEoK3f7njFfOtmIkmBvFc0AWiu1lGXhNGax
F6Lf+5zaxlTg/BgTutdlhaTIOUmPx//ekg/d03kmyu84ukW0NZr0ODHdblggs6Bs
q7boWHSFa88a05GZ4RIkIVfES13rwwTQsX52NV4FLIHEH0PkKD0DV/YQ9d9nZ27I
w7rwJTX0sM/+SpO8JYE4Qzzhz8RYS7w7/wmOiB7qdnZfbze87+3YWvivPJ7bccn8
qlLv5L8H4HC54wxpVNvYejgYc8rabpmJAbuOuZHBs6Z1CKekZz//83fsGqXPhqre
yksjRobm9VfrgGuSVR6LFb4nyH+4C8cq1IOPpvdKSXnTS6nQjmH1t4D9VShx+tWj
v/G2k06FKR240j7VOL5G2zHmfIYIsNT82+ctCOxYN7CL3aY9XxGVw5t8roxVU6rQ
svFpXaKmq/8pa/0Tdnw4rVlc5RjM+pqZ2O6Z6Ryb+SheL9hosqzZ3Mos3OnGfc/9
RVgyEfwGPRh+0FX+wQqHMd9aojZ4d45DmzUMDIn3EZ0ETX2Av4TtxKaIXahMy8X6
INJy4KfiMkxXYpjGuq9DD7YTECKWM0Yn7sK2V9DWh8ZwlYQXZB00a4CQ3pPFgBuu
SdJ4TI2frTiRNG7s0wjHXow5QFaDQJ8KcQDcW9PcmzGq7GIFFBmDIo7/LWYFoDuo
nFSaDPxxH78hfwgamRvx+FlnjxTGfiFNWKX2g/Dr3FscXZngtQUmgRIEC2B4VDIp
LVr6zzMEvcdv9ZF8/+2e3KRnuxt7W2Pudj8j+2l3dDCAHkYh68mEUYUegjYVEb9w
BhUYsHB9INPOm198CB1rp9NtG8poYaMjH1bS+e0pg7RDb0y/uc4cflDTP03Q4fQ9
zdc4Sij8tSgRXmSqW6ZV6fxljE0Cj5uDMYSVJHVw+jpcEEeZmv+BKBX5kouShZAD
RK8PPVKN89TzUkFQ5of3GiDydNwe0hTQIQfScDB3AOWE2aoyC5Xxnh7q7CIMin+p
g1lTe1POOTzIGzUnGea4ChYDwM3M8H3G0HhFuAbMQx9s777cwhM9hYrjrISpNrdS
QrRUjpjxT+mNehTENImqVdbK5RG6lMUK4ra9xUMnWZiPTVk7rPGEofK4u/XziXEX
P0kW3Ra0lI5QT10kRxEauqs/5kesvg7bz145utHmH1ITI39Na+6umcT3Vq4zX5nr
IRZwWeTST/iTu89u561lOt+508qtRKTmZEVLqBseCuhSiwkqRCkcenESFPeuwXSN
fpretdcmuBIhscJ9/QxEgi6Fo2Rv643cQA9T+3XceKZxMoIh0pNdbQ60ZzR/6Wd3
jeYaiIb9dvHRQ64ETpCp4H+1Ms39jLDgRWQ7qkM66jf8gdUio3eqwglPdcuGXHqC
2phyMurIcyvLCvWSYXiqkut/PygCcPumK3cCHH0fERoo6mLk2NNnkFWnixNmOdG0
rlWa/Q6urR9Ht6tjv0nSlWs6UzXekd4mPDxCFs8D7x8Vcu7OUU00WYvl627rCP3c
askgvW6qeYslooyJ0K0TWBgarUpwFUziF91nJoD0ixsIBKzgYbaHB5kJEoJS0ITG
GG5u2Ls8mfPYkbWZH9r9lEfU0WYSFuW4SnwEKqjchXFA+6zFswOF7JM8MCvCZ44d
3xVHrkQ0b/DQ7SVrVRbyUEuTViAoMI7D96Cwx63dFD2zBpMmCjaFDxe6pG/iDXBR
Xe8hqeK4NxNwkmZnRKr4zPJcuJmF7iWSb+yvCwuVeyk9gp5r2FIwBhzISPoiLhre
Bvu9avUlbB6zN1e/QDJPeTv2/inZuKZ6bch+Af2c460FdxkKakHpDYbi7aNycWx7
rfMrrEfwjtZU3MKNnsk8hTsvABg+QIEm3vSxzFTM9SYxbO3VzYliV302jyBg/nxK
9vUrU8LBALSh+BrzZ44MR9KQgLeZuU1LkosyTHQV8ll1z338g5evyR5cfw4+2nwz
S+JNJinOuh4uEsOOfEYh/DBEijC42yXN4TuSFA5SsdCgxzygIdc+9l+mn1glnTWP
Aw4TDl/cM6Pp/aSPkREL7kvRjLBnfpyMgSMMhWsRjiIGg1pooZatVUvSZ9ka+4Kc
fJwSMV63K1J3nF8oGgNp+Q/n2OmlXU70dd3qxOyuMTpT/VFGMnz0GRwnJqWyQm5u
VNttJ1aVVUqYkCCi+20dL8FDLNtn7tZRIefrbaaTCAHhZWGtyTx1oA1vC70a6b4l
w33TLtQcajQGNyUYtubPJtMxS6f4k6772gd8m/lsoeEf0trSDdBNNuahQDow68FQ
ugcZsDttG84Vh7Iyo9k6O868YFDdlC1hjA18goSGcMGw96VoKviuQ7j3W/Uop9kN
UTa2ICjL76nTsMBZukNgXYCbZOzNFXFLdcRHHABdy98XrYSwbIGnrRxAwUtwVQjK
W8v/ql884OciJHrgIi4DrIfh/FRvgPE8LaHc7/rKDN2+L9sE4gk6xNpDzSkMKM2j
IEIOt3CiFMvbKK9gWy7py1ii0Atu8WMUVEXFsobGS4BIotuWdgvh9icBeyUmBnFF
qHCGua1xUHHBrvm5ES6wtYBF6MqWVuKurWcS8cv26dbgH86eHN26AWhihx0ka4uj
UCQpDwej2PZ3DBtp0HwgPFVBsL2cbk4EdgQDhpSsjl0rAbQyUz+hEPZCx3sZEmOi
vINasXDYuzp06DyoDJERrMNWyM3htw3j1nN4e6e4xr9tU7zPWJaQlFgkyTSDw4b7
EsfZBB7+d8Qsz9+2LWNS/F3XnABPGt7alTTon5y4fASggOvVgmT6n0KMvNXIilin
6Zao6V+jkOy9SKNxB1yAHgLxOy8/oHXOZYvdlaRnxMMMHuwyXo5frSBUbjbdZYir
nsS2KiwTg2gMexQQF+JiW/ryl++ytYbP1gt/+6dnnxsOfruBHSMTEQQnf6I1aPAG
uQjxHE+Usvj5sB8E8PYHZ96xp2dhL4QsaF+zXLaVJl9dSDEbpVwGGLVixU0zR00U
BkKZ8GBXwW5/sYjf7+XM/iNiGdmCJ5aCgHPTsN0CYFHmBIYgihNX1F8363xrE36A
NLS3lGtsm52dlb0ITKSl/Zh7mzrdRtYoYCBR5nCGw9bw6luUKWj9uR6cEItjBdo+
MJXkFwB4TDSmvQNEpmz/dFuInoJ9kuDBPCo1umHl43yeU5Sjg8J4K18SVuxhpor9
0sLryIcpEn1Vw3eCLrw/8xaPhrRJqVrsIcuIY3ZOf/32LFgpjRgUVw9go8s8UZ8K
VsI1qlV7gB+LQrrq3LacrVpfBUVOKIWUOVCjZSecW+33AtzOSs+vDLpX1zdRR3qh
FpHp+uzSphbLPe34tCo+2N1gzlCgpJpgxWwnsScnQjO+DMDhhEk06bZKy8qQsc9e
rBKj9ChF8eMg4ShfCxS2Vf5YVC9gNlvHUZyKqXx1I7o52nlltRgHjhOn8wQZwCIz
gpGpJPOs/g6SqEoiK1X2WGs3UlNhGAD0GCJ2/n4dLMYmiq331aTAwpQcY3zD1XgJ
zssyL46H7WEmM2V+2RAMitLDuXh5gKMX/XvQGgXkNihmt3aWd40o3MJkkIeSWJYw
BCWrxe9kHus2Xjy7Yl4pJnxiH5Dnmyw5FxusHlRBsLsl+qzBgaeJrQ7hwpyaxOpO
7E4olfxj5+WQme6/eKWgob67cdiu4zNFNWYFXgBRjsx25dT1ZMZfeuFGh6Ifms0n
DpjykAIFlZxdognrvgbGAnYNqoIup8+yBaN5xxFZepivdX2l0KNpNAdoo9bRTbJ0
AB65PyfwKuKGdxYmZkZWsAkU9fGCNeocCGls2htMPLFuysYNmJP+9FW+2I1jRFBP
NBfzg41aNFmsmf4zqmm38uwKBekR0ztcpThg9HJUxHLp92XoabJMPdyLml6Q7dWF
gtp4mt9QhKa7n+nAHcVYWuo1nYI8M21aEQy+1sS7Gx9BDsqAvj9vObl/CvoU5ZzZ
UNcoUOvPqFocROtX9XjJKyDEfKuWhLfkn28luhZVIfyb7z2TS9UHPp5IHa9UeI+s
dsGHvJtnFyX5B74t5qAESNcIFT98a/Ee3lURJu7mdxHowRYZtdvAT3NtHfVuX9Mb
dnD231yn3qHXF7SGPUckjZChiXE6s3VcCgG+9Sy+EbC9endWAX5S/9U4QbomVITw
p+8WYnlav7X8FAkLnl2XIG7qabDQtVv8GL2ixCvozu6JV4v0jQkgko96BhsUpEa1
o88Pbe1Y+PX75Hnj+XdbhW0tdOyIzcy4BiLqiJcLMpaSFhqMZAqe+YNygZIOE35J
TWsdy2O7LcXYLbRdmkPcxQtQEduB2rZWkHOCyreQsR8a3f7n5IoVucQ/EDBdWyx1
6OEbPXpjuy16ojTXwmFbbLq3mj7RgjlhxSyOsh4gTKsNdXgIiRlHSUP8hDR8KUX4
X9Zabn1XLyOL4DJhfv+H1ZH0SLARjXJB0iHnjzvBI8Pq2tlFeviia3gfydmgsbAs
5ljdcg5e8d02RIkQLY/j4X+TWhSt5itWr1HWb2sFwoEgXIwUXxhKjYctE9gViNBJ
C8Z1X48iZakMYAW9JI1DbRoiHOoh/0BHhV5XmhJucQGhU0ItxKONxSwxqikjrAYM
U2QMtXsZy4UCEgwJgkTUhLpKUEzvCrb3I9pGdHFTJycdDs0vVcRT0MDCRRwMqrjD
jaqzMSwLhHsd9wlVjP2pO29DiPGKmnKSfvZTmPdguVUDdFyJwxRuIZnYor8k83hR
8ruWU4rRFj6JP4/kaSyPvxqREw+bcxOjV7nK9/s69mEdM4v4nPNlBU+eac5N1G5y
aZQQD64Y6SW6Vw8pNVcvlpGBCCCBy7WWBkpoCdBNRKqa+GG7Sh2lOuDWubWOiU+R
r0/NTk7zWBybcQnToN/6mdit6uhhPRCAVVxIhVlPEQ7FCscO0usktJhhb56CUKZy
xQbqtSYUvw2FRanzMMWVQMEU8cEfNyEV6UFMiAfU+xQG10VFl/H4pRE3hgWwFOXI
LUPtXjoHnE86knFP+oN3fAITls0Sb6vY1lYO65I/mjh64GoI8qXGtOpGsZR/+FDP
LhiRtgo/MWXg9FKY70MxeYsjgvH8VLO75ST/bMYtJJoq4Osvy6r71/qO2MirNxzd
yLg8AAt83jvzbQxlKht/3x2V06P6lfESMosz7BFTqnX/DT75iZ62onzqB6HWqP1b
gYgAucmEhqqC48qR+CKyEcFPfqb3Hw1b1j8DOTjI+0HEpmztIEpaAqMUdzxYo7E/
7JDOkZ7yfAeAQToPBNGg4fIcUI5i1ljpWPt4uy2JqRHSVar9MC4jlpVfFht+1npd
+jUBHBHDwqHBU62l6UOvtyWLUnHo9TtoKc2yTMaoM1V3pEvzEveEOf0XnxewNJln
lOAszZxxN7Dri7jrutdWgDIDBrquvEQAbYbYIwXxVule36v0m9/AuiMQ9UzLTg5y
e4Bh/Bx+AiWA7RYqVrOmM29WwXe4uEWx/EabDN8gYKGiDx9S4tgYDd+nqjP6ioJd
G6wsQ5iO6pnEz20nh4RDhdupTmN9M4P0yPpLTzElsv+6XRG7hRAeCAKq0ViZYf+E
LNIRgKD/nfiVVlpY9D4lvw4CeLDRSvSOqIQZrO0ua8mmJdMzV5SUTHNWCrRS/hKv
mIqh7rNNu2OsSSPOnft3hRddXycp2tcAu2OTNf9p2kQf3gkVk9oF8Q5K3RZUH3UR
9JBnJiE8rBUTQCZve7SwyPbQ7/1OwpOv5uvw6uPYEkdr8N4lW5sCanNtFTA/aBjJ
F4dEiixXFqM3WSgRb4flLjiGysAPq+CxSLV8b11cGOQIuJw0Cgvv1vG8fJaVyGIt
Ivc670TyK4XBsIKSKp2lr2TBc+Z11iT3JmBKuB2aLPOSiz3Rvibtv6qYAyZid6/T
kgknnBdKl5In9jQFCYm7U+NmlXWf6Anvah6HG8eyQtwbWTQSa8fsiymiAXyXUCYl
aFaeMPI3F7DilcgGTTm+P38eSnjoF4s/ikK8vpF8OsSVt/pCq6QTQTdulYiFu1lA
rbDolVSIbhPKKhCKzR4m/rlxwg2bxlFEe9NuDhfENFkiN56IXYDOB3d+GL/r8RS7
i/DKktDOxO7CeW7vpIVrqgc6miNG9AvDsYOn480GrQrLwoqZ1nnpd/OaJeznonqC
2mbR9oYPjEYlOJXaXb4u93ACR7f+utmutoyks/ZxblZ3uI5wz5165wuCOFG94rfD
oISP1i3i4PrmuaaqCGGpizfs8gKWZ5MIL8SXz12z5dWsAhtVFFzXW+GxQbp385vf
KEYOY2a0hJXlxhZfSIdrppY1CgZ9yUcK8F1Y/jALLPUOir7iT//dVgohXXrFZgoL
bjazaIdcl31B45Z3QWOkAv+zGmDeRRnEgl8Gc8zv6eHNvv3EaSTnRBdUvaUTl8JG
yjn4my0ndYhDIdmFYKY+3q4H47dvPlEQrUX/uXFyL76qiK6cZSqDFGPpg5776iFv
jVVfc8AROKrO9bfhybv8B9rg3djam+hZ8sZXwHi7Dn0e15lsEgniI9+m/th8QcCf
WG326bqvSogubp0XLOvgP42KRwcet+Ck7L76+VpJxhA3Su1Vr9J17SrMZIGRJ++S
Zl6LXdqIEhxfibD6iRojBYSDS5L9qNoPHOpdCKj/ToU2au9LDAKjsQemCUB5YY7t
5N2lbUFy2j42t9o1vGXQzGJ83QkBBx18N4LkDKv2YGT+jjl8ixw5t2ecjwjFb0sZ
0YgLTX/x15lqgy2T526DI9ebuURDsySVRovYlawgu26bi31jU3Yp783Z6PUMKC6e
8V3C2cR4s1aQukGpBH4zzPqih2fj3clpsZXRie64wMjrZNDn3HqdyaDzfmL7jIAu
8r+4jbDEk+nKIZk+rFw4TXH+o+BGNIFtPJRnNWXW68ThP94cDVRfndX5/EjaBg83
tKRyz2IqtFKJz3aPc+erwPURsjBrUt/Yh7W8CX/w9BYzwANN749NclVXSktj5Dyh
O+9quheHRFLYZpqLXbNWvuS8mEKLZgTXLEFU1cnTjetcSw0jsie4qy3m1J9bmxj/
BWfpDoEByljy9DgOi83YFg6TUmVidEBA/OiOb+Su59DFxz4unv2252soiQvSa/oj
9eJRo7NKZXdXM+eZVrOyUqjiB/k3aiRLVpqcsX0zGv9b+T4HNWfrU2zdFjxQLrwu
LjDO9HVwW0euhgj/mH37fUuoBx2FI2/rirMY3N0abqGWPWyItl0C1NLDewESfLHE
JuJ9CU0HntyDwcbHFNi501KSLJtkJB6JYCZRHpTWfA78sul/eiw5ZGYayODHNpIZ
8tqH5nNh3yLwrpIgQmaTxG8xtLfoMRlCPqvrv20Rmt2yo0gBkm4wEB7ejhHHgpwb
sca8zPw+93bmy8FY1EHyqdihb/uAk5O+y7Px+kgtmervpOZFJnZxBLG0GViYXxjL
pB0b04paqkapN8HEVnZm7nyXw9N32/UDePvH/19A795m3qH/N/zUSDkJn4gEF16X
HLB7///adbdU2L+sh29ecARj25RF0p2tfDW3ZLzso8uO0oWIl/nq3mqbUxDNTg33
gnB5OaTku5u0eaQXFc15kotU6ywbSQjWenIIUQA7EtW77egp6w1NhUqXR2TEOhXw
CC5SciFns+4QMPIFPDrcEBb5wKAmnEUYTtmaMriNxHJnxGR5IsOz02cK1yn10PfJ
qEI0Z3LX3tawGx2DfCkCvWPOxO/HUMxjXV5+4fnyL9MJJRdYmAMVq3FvplZ+Flgm
499gwARDRGnVKC18isPpglxC6tAaVyqoN7rNZp12TAtAwZSPyJP5VMQIrFWKTBCj
jt+7PymGrHySXwBeRjyzDIU687YlJVspItrYmyUI6KXQXOJWO1+BOBrvk6vHoJY+
1PR5HXZLb6n1bQDNcKahnimOwp7mI4tTTMQCxJFklvN1autlIqewuC17LGMhA9hM
INXutbXvP3zXT2a5bGNuM/J1CLcldziRDr5lPDY0Uk6A3Pze/JBeKrRZIiF1rkc/
4YcDY16i7sr9R5atD9ryARrQBsHld8C9s+/M3azXJXPIGyQ3H+bnlmDzJ2EmYdKZ
vta8Gtxj9eDkTlgc0IahLvEAxZRWXIgx4uqPkIDfO5RU+aB180L36HK/NegM0HWK
SlMlihECmtPv89xPe0aHtC98o82faSjQlAw6d0r9eU3LS34l7gPWTQfdaGOPuuib
SiSWyMu0FUJNxGT+oDufXoVXZ272mG3hxlwkP5APdED4mKzOvqj3VhkEArVD8JmR
Y0KvOM+kd/4P6lfffPfO9GMFqdSCqHXVJIA4XAW1A99q59sdJMfA/O4RovCZDk5r
O4IpL96QOUyYZo7m5QL1SGY6lSAMWonb6OjJK0Dr1XAE8KijuPPiJyskNL2yngyI
hDq6MeTefYUvg2SbNKif4w/JyfP0aBjzSlBjuRg23uFXUuhGFTmHAuNG7Goq/9nO
21owHdM1DGGSK46G0rsMSHr2eEqCH5jHR97DOfdUb3k4P9cyOOKL2dwK4+USGvP5
hxTtTo4sqUlx056trPv0VKIhRWYlu+fEBwlYXOTFmMthw1m/gxbPASUfXBmIdptZ
JWpoTQ1cjBYaUivvZBLVeDBpnACrjU4j7dNsF0tIrFeH7HgTHElUTQwt+aa+YNwO
Fit4pZr56wZBub+ybPxIi6m+6HQCd/AUvdEsHttwA84Q+GkJFSMoWljSAgkvZIed
Ks5I7hh7T0GMM8La4/TP3mZRYb1ijv9DcVnmfZYcYEGeiQkUHajNt1/FwePo4iXI
V13OSzX5ug1FIGRRd4bkWhR9jHqAmr2cRuD738IEQ27YfxmHG7ztMeQx7NOnBBzf
wxQEYn7djeIRSipORIr+vi6961nnqC6huxUPtWY2t+fdzYC0vj/FGjJ5DR1P2R2N
1CvwgXM5JiM9qfNC3MGYdOFEs6Z6kDC6KlL+pKGBEdWxB0tm6sqWpKxhqLelExZs
XtH65dpjzmYfIKsNHqDsaBa289Is/FO0OIymDHEaR9JEWqMqPY7gsZJv902P4nMk
6xR0l8yyGJ9KpMZOXI6/17a3bNta7p7StSwoM8PujcpmzJ5k65tcYhGprHDR38gP
+Ptvnr89plBJCNUaND4FEfNpgLrm7MFuQR5fWgO2EUgU4xDZAGoWGQqFiEF9qUnc
fEewLlsFDBmMwsJ5HqLhjdtmktOqOfOEZss2q4aLrf6NzlX+JPadTjLY5dNgG9vY
F1F+nBXzADFu8bBYjJcbmNTiIn3+kmHtIPEpjk7eRwBLqPB/lRE2HtSYBYvz8UEy
FzRGQYXjtZdI5+spvEg+BnDXyTLjxRiZq49EGVGuUV/0nxyJ0ORhi4sIoOH9+h2X
MDLD/8oj306VSQNu7NmtiZnBdbigqyNahDzniCTH6Ds6c+FXkiis/yjWCBOgPz9u
z0rOhWRGGGUHfPEWgJw+6druDtdmWwPpWIGZjGsxxJ2YvN7ajCL+BkPwLxLCWxb+
burRkD4UN+IUAsjP6pfEpElmd5edajD+9zOUusBPxcgRtvma/oa1eK9+wNfyDdho
g14RhgOxj1yguKDyGhORe9/dOF0L9O3AyQRnXc2FTMSItdAhJXgCH3SkwwaVou/1
IxIQEtUS+AoJQpWx9XS999gwNRL6qo+H+PUciYykPfuzcEmX9+V1EphjYrjkLuOl
aK5C0WVmmg52PxwclvaGwvNJih5SdqP3TNK3Nt0DhNpOCDFpWxFtnrmLWAwPTKsK
7j3WmiQK0os1OgXhc34fACoLr/9weMHr7RjGVVJu/EHvo6XiNwDEkYbdL/3F/6Bg
J9bxdrlvawmV+HFHLHM/CgYv04BjwxJFiZEdSbp4gNJ646rxTg7IrUKW+0cgobqc
U8NO1kZc+m6rFE2DZqj3F3+3/aSYJXR2FcEMjXpERxljhfQLdGE041DIWkE4p7CK
sltRqwpl7myKXiNHpeyYO0Jxjh4E0d8I1O7VPX181Tw5wO2WcMmCZhCHtTPzGsWm
UCfXpuLJIcBHrvzUlKIbs0+822wyUbLWwiW/Vh0ocrmTvePH2QZffp86PHaDsEaG
NcEyIYP3eNS4vpDlgvQSBfeUM2cZolJNasukTLjKuyylEQjEPhK7GCPcAdB02d5k
jljWN8R52Zz3FoAJQ9ypG5npJYKisgH8Opz78x/wbt2zbyRgXICie3sjggLYuApe
KgowKZkejpqo1N0ochwf35AfcRfKR0kjDpPqSS7x6dzqDIxGa3M1MOawvvjduRBd
kBQU/J+97dIiJKe6arg8CIqmATWRtFrWTpwR0WmPSEsOnxOjDukMRbIGqzuWXgAl
Uz9Y+DxDgsKecLhDRTGfP85Tad1wG6kiiFt+1ffdxzTFmIxY115hd7ZhoNSF5y2T
fI/w/AnU+ujvPYLxbUPgIyl0DO23AlKOD1C3T2UnnPaUO4iO28Ub0XC1ZIAJmDs3
4bbQGioQb1ii2tkPoTRKu7UpnWMJZmlO//iBQ/pKX+9Nu9yM/Q4mwuBatVxCot95
S1kY/Kaq/eyiUF1Zdg0grbTEqAZXSffTPGyocRO5FQQyWdhN6ONFoXmYgsd4mAzS
G8q7IiD0ynbx21x4YzyV9Lz+XPdkGyHxGoaYa6R3Od7AsORgssKBoQ08WnQCLL3I
983SWKU+5Hx+JbBgrl5aIa/3HI/IchKd3JamGjNDQLCaM8c1k7rbEcbAFU4DUzRQ
jfJ/DdB4pFVURhkBSgA/aQt50Pv1vz3Kx1x1Og9Sw+r1yvThbVqGMEuLgoVNQwvD
6aKsl1kRzUd3jj91K7olVnx+5B9t8jS6c1Z4uHnNJx6g48xNifD/SoTzyI10bx5A
WTaKYRTgN5C9Uq5WFubA55TmitVgvTg72ZTwpizVq+IPALC8h3AOHa1FVKUwSoVX
5QxKY4bKndCGlk/oPcD8UWtEdtT8m/Rq6rW7L3noseTftl4CO8rB2+yhP2ONd+n3
XZTv0Ay3hpJmKxiIBimXaJp5umzi70LO/2qOWbeUaRQZfbO9ldDunC9im8nZDP4G
uN0DjJyaW0/pDrca3c+JUarz0+9sRepHSdHTe1A8UNqfIel6rF63jYAlkzEnALMg
MBaFrSpeja0wtaSTySb8DzAmUg9csUe+Ejjx3u7aglmRVUACxxPInLG3zjQtELTP
+sp8DUSX2YzsVXZENNab9n+dQbTR7NsZN0xd0ZxtM1LovYNDF2cqTDW1mGi6IjHB
9UlYkd6BPfDoRUhnJzPuFBfWlnu8XzMv9evGOnx95Bxv/SGrfnj16072UuQ658Yn
6lxmKTM0CHWaxaBJboy1fKzzS557I7Bq9El/mXWMbzVt6q7Six8iUq6zU6MXfCZ1
cAsPANMGb3tTimMU9dhMfE57i7hEtK56lgCmLf5oeuTnwLolY835fsRdGhXD98H+
Mz67+kkYD33L5e200zXHPRZob87PY3BuVMyjMnbpMELFw301By4nwt17Qur/JMfZ
MCodljvIhTObER+kgjKv0uWFOV8CgdzPnnCXsugbtE4XbscV+PSAbGnEXw6G9qRH
dIFwwhiaWyv4mnbpLFybwx7pLRnXVhcIdlMO1DKCknrpltyjzcJJaI5J0tGYrkBd
q1aBDdEzuGR9LT4NnoB7CJ60C/6IpC2DooTxNZfEmzdvoOuP9xn07FXujMyKd6PG
W0xWl2LvbzutA8sv+MNrfALKRkd+j832jTeMAtdTgH4iUAi0d9dH9X0DSfHQKX4r
rhaA+3py9UyL5Nmn/vG6Yl0R3RH8CRteDln3RSoWmK5ODLVHVQ4z47Edc7omiT/k
DNHbpghoSeHKi1nk3HTtexzH8Z0HqQiSo+YkKAde2Gp0CifkiI9Tb+U0mDGCcxFc
LN1JecYZb49bKrmhUUkdKUqIkdYMUIUElqkeUeQNML0/7sv3SP1igMLSgzK6p0Ge
+Zk95Y6ct9eRfq29YMPP8VDqS9dUbAhd9ufEzEYRJOL9gSr7Bqcmt6Txqtzh3lz1
oqBgKwZyXCtHE5Vh5imxW5ENdnc/IjTxIP6LRemRtRcMJyoErNwWAqnufM7dGbLk
2+hj8NBWv7qeaYbqQZdT4sxOKBszV9/iuBDsgJODOH1sf86VZpRi3sz0NuiJRJc4
j6hicycjH4nyX42cMDi/Gi7tHVUomP12+yMr9A+snG4BKs4WaT7E5qreL5ypBpEu
rCSOBAWG+MAPcoSJx6ork56sWWfnD6jTdmFCmig2jG5GkuuvMqAuq4FekPPjxF7l
bKEJQOqtCb+fzikW7P7z1EZnVKiMltW/1ENWX7u0tsfnSQT3xGOB6N/MZOYpYgqq
UzIan/h3FfTR6+Ei6dSaTFU135jYaxjU1nRI3qbJTy/6Q1STgVj6z+NA693YNt5j
vduS869xepOWpM4adJv/gfz5zhk0QR7pPlZXxBSjcZ3EMJqYblZQfu2treYavtHP
vN0XfVTQjIrvPoORa2LNgL04jeZHAZ/2LMn1MG2xHjHginbM/m8HI2T3cYgVm+D0
PknoB9Y94F3noOJY2ov5gmCZ1wDzBwuu37uLPUA2wflzu3ucn3uuadQ/XrOcJZOf
cSB8hSVhT2ESjqSFbwYIxuk6OxeNn/7fmIFpxj7xlhAgCy4Bb3vG3SRJCEzlGzdp
8tN54p6ObJHo3sspgTl4m+lLhLqyAcXPUjW/GbpjDdDtpGqxSBx6HhdFJasBOWo9
uGk8rZsceien5MfsxbvJIG7jaQPQ1HFE55FcW15LbbwAS4uKgHjk1rlKZOWcD+wk
47tPlkDafU+cEocDjSGkdCAvabcNwlyAFp4W83vbC97aHBic3Zx77hJQnR5yLd+E
CDGaNllEMzXA5/ks/hbgazJtTm+cowYu9H+u9y4cQpScoL5j4CLCXRhVdVHiWaAT
uftBm48DUppRd+XeAJUpZJYb5qQNkK7UVwmjIz8+/6QFVPDU9jWNHemHw1Q260P4
D2ljavMBXZ1X/gaLfOjssf8khGzveE9P3m1bBC6XWDBkEDbchNUi2KIyRshOPxC4
SMipKtdJjnULh0f8FqwgXGgkc3c79RljEmVC26Ktl4u9hhSKfYpHIX01yuMolmOz
yp4k0XwsM00B1xfqNWUAYokAs6v7eqv4cF7ubix7VdTWrEzZWEY0q61XPYmpEpiT
EDMZN3wWmyRaSkJ0USwrAO8eZnLryg1JbzobyLGvfszUHKCVPBp74MlQZUIbhVlU
F1vdV3O9/Zn24nlH3EJm7xkwW1P+4SHX5NUPDBbagq3zW75wpnv9zvKRbKKC7ngS
BdoW8K7Lw5v1D0LtesxAjKD4LdwRa1HRBzleplJ1ro5+56arzRxn1vgbE848VQ3d
kHZyFseAe9IOBSA5TkDBoOeIAiEqirQHBif/wpyQV+PLAlNWCTPyMz2r/OAWOmpN
2sXil6TidU8UKqL+SwMimfkdyl0QaS/4jLWUU0USDvZmFLybLzLv5pSLVkyc3Y14
cjjG/p7L2H+n4ucd29L+CbotR+SKAL9ndO617dKEix/umZno4ZCW9IUGk+ZwEcRy
EUmrPWnzrVKPSULop96jPAZcOlopCOOLX6zTS1oLnERVnLX2vTcXUsvPP1TgPc0j
wp20TghIFFh/hmaV6f0mqz7VmeGMm8XsDTi2IX5/H7LDxLPlg9Y258URXTx4PpSN
YPOYT5R3JGsTYbW4qKRd3TCRRQGmrH3lBCLofcx+qrxB/xGFnYw2MByspZ5qQJ96
p+g90qKKuWNdCv+eVPXtd2hyLNDYc3OAm0K9mSXIZcA+K1j/khJXISlknrE3eMTu
PH50IjU1uy+wWLMXBYbhT6bZmG8JoFDK+QsEtpA8GZ8qMwGGQ150SE4gHuB+1K5g
Het4NM5+DA1mZr/IEowK2+UVd7s6S5YyG3PcwgG0CbbDq3E98R6zAA6OmQxla8VL
QyqjczDtzEbN0s078LBOf9qEMJRTAIRT5VFlLMUwzJBsJWv3yM9wpoz1FyG3Z3Ia
V1wLemNLT4ij2Av+o50ikoC4BkSPCGjXfuR29eje1l/W6V/t5gknNUb7K2EA9FCn
3UndW+pc/JQ9TLUKGER4e3S0PGJCGhjMpa0qrY0sYeeCVJlCzbxkF/xYwwDN1ksP
FVu6HePSZgjFt884pApoe4WPlV3Ju+tKZXE60wF/3GNtJG4cyPFpJP4PJX77ftzu
wdWWEWgmNP1612iBj40sad6VTGXaZ50f34zIaYsSCXANwTcWZ7ymc8UFgi0Hn3cK
1QN1V0YYQPgGuxtqponVs3SS7qPXC3dhdyum8hCzBj/7oyxFsiddTSnijCsBay+k
IGrWzTnjKpQjq0+UFmjcx+FtnbzntViL/u0PQszV2AWlpFZdVD1I4MR6/Wi2bT/N
VajH1CBGWewqsqN/OYyh0ltAV0krfXGnv9+iyY9pbn5Lgj+2XiVv2jNa1xdm9+Zr
O+H2Ky3oxlpnBrrEYhwvqARtNlAAA8KoiEp8+lnC0BG0K2c/G5VGit99UOlExXrs
foRVVquxzHiOTEBjCNkC9KFKtSnjYzjeZUsLW76ZDNm3jakm6lTnKhgZXfffzeeG
VIZhv5WOoFjpHkkcKAAX0s49T1kyskMM3ot8/B00O5uOJryBuQ6gWYoresZqMX5L

//pragma protect end_data_block
//pragma protect digest_block
hvdbAdhz7lg96ayzGHSaZwYW0gU=
//pragma protect end_digest_block
//pragma protect end_protected
