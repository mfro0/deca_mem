// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cFyTE2stXy79mwQyabcVWtkXG7cuPaLIueIhiGddiRjG6ZNoMimurOboqbniZHEs
TTtNDO1cFq3Hn9aXoAKEIMNLPU6TIwdjqIsLoJ1wQMo3yYJGgjrEGDYdMBgetrso
W0XDEuz8xnheU6N9m9Il0Z7RuZu1CZ0Mhl5SDks1DUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16976)
cqu18CBT7irOvQ+YjAL94ZsmY4f2MPPA5OXRyEQjy08FlTEMz4eEllhTFjB+GXF2
rh5ZzOJHWdRrAbWJN1xfH6Vm/MeTSbcA0/mkfXJxPuJdeaSE0yzDghPPN2oFV2rs
XP8j+Si5c+HQGvFdVhUKEpj3hhieUuvyHoaffRFF+GDg3NuJT4Jd5l0cUblJrH7s
zYw1EOnbgihABGb0SFuwExIjkTMYsx96LxaqpQrdXWhmTQzIho8K+V6gq1DA4eNG
OEaXU+IjUYArKiec/ctPodCU7j9owJ7m88DHYCAtFWRXn6GTiJZFL2qbVR7gBJO3
nJdI7hk8ciDngkqpxRJwxW55v/Wd2mhaLyXYKj7w6gZ8H/cRXG1LTVUp/qcbh2WN
mpaGedGkox7LadaZuTvTvcuHB4pvcPTpRdKYKN00LJoXZTxlkEhKy4cQajQccIKZ
0Zw9ISBwi2xpHenkLQaCXov+8j9daIn0NWjzTf9Hob9H6225OYGCPif8pG59qMws
3XG9DpP/AkhBJ+n8pPdlvetqrwNbXYMluhDVSCx+gnp41N+o0kE30ZrEQJw+Pmfc
2LACSRNeDIGbcQergx7jM+rGvccvAQi0Q8e16IJpt/Co0pTs65nqZ1Tz1lF2L3TF
rwTXA66GZdTDBANhfziMZd6f8FwmiFKXFjPeBACNuRUIdV9WnD+7sLTWJkOch+zq
OX7uvjWtJIXKrzbsi40r/HW55A2IH0Inx2tJNmDfcZZIrpDTXe55qIVXxTPKi9Yk
V3bjy4TtjfPPW1aTTY2kfLRhye5QnDPxX2vFeocmvpEK7WQyt2I0T8VP8CV8aD+w
Xh6M7/K82KNMLsyN6YrIevzjRJl4l9KyW9JgtlZwxwZHW8ElnRnU5mO646JI5hLP
blCDuGNzc5x7gwyQrsV9lmtiwTcxuSa+7ffXNJPi1fnUmKuYiXGMi7jOCWfTfGlx
zzuqKHZrz5vCpJTTXkdhM3Gh/D9fPZ24Qpi8Pc7rxLLTlAcOmHjlg6ezHbGYvJRo
d732b7yye1AxNEoyw/nIIbD8QNaKigjBQkJLqmNThlVc9Q74bS5HeEmklZMDgBhS
YSmdc+hX+I/4J2QI+oSV9t+g3mWYrqis1tzK+rcJmCMFxKeU8LjYUoFo/FCeF2Ri
rcDZmZ0SnCGXL0FE/x4WcTyMQ5DqmDEURYf53ufp1wonnhoW8VJjUYklN9BRQtwF
zgoc9Hk4wrHSZGZrzUFIzb31+2ApMItfPPEvyDtqpMR3ZA7Ucz4y3FlFHQCWbF0q
Rq0tOewhcH/4xtQgOiXXO95bJQH5bmvGZHlVUl6OUOEAvaqj3X7/8/wsoetjvV03
NUZEjDePFG8ATI7DUDgZZPlkVbjErftVqbUmTvIou+WW4Gpd7AFpc3gT6wWLEurv
ukRJvhcSISAXLtmkmcOq/ukJVbG9cRbggase0Y6tKgvqKWf4fDqNhEWBe3+T/pq+
cao9iUlvc/222ZOS0yX69soUNFONUIdAy7YH0nR5/SqGQfvgyycUPJt8NXa/CazQ
eTB8sh3qVco4/6Y3wJOefqQtMOqLsr28SoQ5GAxxLjYN4zrxmJma47k2Fl/EupQ1
/mkQVJx0AJtHiAfyqi68NF9rvshSe2VNB683P2m+u/E496u/uOJTHtIuyQ4wAVHN
bHQfU+8/I4FxjGyhISNEuR7XsC74M8wLVpa8lB7IkJse/vQUM/PpH+hzrV4pjxdU
7XQc25WDpFv4lVnhxrZAvR2AJi5+iatHM0PpQgaLDmJ2lDuzSWMwev95d6VhGZnV
efeINiYSgu+swRLidGd6MB7o6N+hKKyHaBWbL9A+mVwm8EYE379vVttbYTaTh6Ju
QbRzVsYNS7RvmE8Y2FoGr+kK59GP5hLpe2VCFLigLsoG08X6di9cv684Z3DA5EkB
hT91IK0jm6/9Km/c5n+sO31a0Cp9O5ch3xmi3SIvYzAD0sFHbGknCGLOcnW+hcwP
jYd0V0O7WUkpsmXP+H5qwQ0HnkVNcmcKqIBULmYgKt4EFNRnOy6/FHfAe5upGmHk
t92nB5TtzGVlw4eKtv3YbbMU0RmkP3PLcGdotwQ3G4ZO5/M8pYm3zSEg/O5OlBD8
LYkxKkzHPeF/JBLd009r4QuNRGuV7EGlHUHW5OmFfaHR7fNvCYGBk2WNK5J2g+eQ
2kB2bFV7LZE0ZRvcEXmtNrMnPer/DNjkFQyHiw4FaSfnCGyoKhgsYKiaHvbFXOJ3
LtB2edHYJEGbF6rbt4twBOs+d4lPOdMCN6HqHUH+THOn2yEA7WEGA9xoY2YIHl/o
RkUCxc2n87HU1uicCdL1yVQclY269xRONDlCQe0k/TtHXHX01ZrLr/WnXyvBEkHb
06zRmCjY3Sgvo3MPd2FyYe3JuLiMITkv4cGWOhu5AYJhAnSJ7s1kq798JPxc0QdB
TWG9C77eVqzBK4+z3YtvHbaag4TURhuHxbkbMq+tbr8Ptb93hbsPqJaQwT6Rrv7k
FqvkhGOlPzTTtFl1kWp9RNtOlO9sMxHPa2SqpqeMvl4lxxRNjZqapsPzJ7g8LAzC
VqGdYUKKzKfB2e3T/60NmKBFbPluowQ+UipnArBG72kQGetSK3Zgv1PR5C+LCJ0G
09Yzt5zg5svqbmk29d/OjRIsFp84DqEeNsJ65jcftyn25j0czMIoag2L4Nogi7Tt
T6yT/WxrS4pC+KQwOLyLQc1Bt/J2Ze0VI4ryJnDA7DIHXvLgx59+EC77vMmRnDgX
+TWH7XhaUVOlRV/6cPh2aYP35FZqW9qE4eotCOWiCcPewxfIAQrW2M7foK1Aq6vb
3G6g43lVTiEj1/iypVtg3LhV7H1hllz2sutNh/HYNtSyClVUmWXemtF+k3KRlmHT
dtlxBmJr/n317qh22DkI4t6RtRnCrTViATMA9q9+tUjJKzZoGPTMdaDBXWFX6Tth
r4mq84sYSAok7AEK8prcmktkaEUuyMOnMuqe9rjYSbv44gPirrwouU/0mV5Sn9KO
Nj+7zjKL0ifhIT4AJHGhKEoKpxKEGa2TZjtv6+TUzATdtY8dx88FLQVOM6E1fUnV
1Xbs7EnBFPHvwWwZO8NhIx5CL35jBpFY74oz1n1RkKVGTn9ghQ9YscsBFXHwkZkq
Qc1AXFFjJPWYJ6Lwd6IWnIhzpxnFVO9kfM4W8efR0f5FdVYlEllK7lgYuC8uIQxV
CzJq3WwsV6BbdlyQ8ubJF70anzQWSFFQIAwTnNXy6YXLn8pHZi+cMY5QVBOYadeD
0vIUBXQqXnvoeA03PkKFGxq0wXlFOI1CCEcu8oM8yauz5rqsgeCzQYZ8c4RHUR97
v/HVqISKjqSbxVq8FrQkW4PYEB6KlfVkHi6zb5XqMMWo8OTVIWixXuFNKFu4lt9I
SCJE6E6kGkRwN3Xh+EAwVeT43gdGE/I0cT575DjbX5lAfzoiABg4xgbzR5IGlsAo
SyNC55WCl6AIwBi/ATZzjovZTYC/KUBP/So2APeKPd9FQTmv2mqCOxp8AZIvEKLs
Hbbt3uNMJiWOHln7gKa2ElFUHaK02o8a5ToD+6gYkrWYI7nodLo9XuXJoR4jRTvV
4TwewNpIJsd7bXDGp53SYTxG+HIz7NPMJyCYD9L0mXzzC4FsPhVmdLwrkS3XUW8W
LiYvMZrqUfpxGI6uAU9o5Z+Gf9DTT/ho1z+bGeTnhRz2S4/vjDF4+u+b71F5HpLq
pPFw0A5NbN1ZU5wR6AO1gRUsyTp3vmOnE++5T5dCdDctmi32yFgDrkDkSFZWLDTR
T+Z/sgld24ID9a7fzVTH+BPVu1vtj+kWtHJqR65XI1TOal6xUTd3aNWU4G39oSWk
RIgH5Wu487D/MNEBPatCCZzNQtF0CyPuFZLNjdFRn8XAL9hYJBb8yNoyB36rDL4u
AJ+HOVDYjFRpPODfYLFKvuM/eJYrZk507a1LZHnXQ7/9VbfdMMx/cwNgcLxG7cXk
2C2dHzGzX2eXRONRG2QZC5cF4ofc4dsk5v2gbWFXEmz96yToLBrb7J+ixkOBaZ2C
lXWOb0Y40CAzBiTY25T4SiKPZn93w6pHx420bgmWKQcqg+jOvVvic4NvDoPPzELr
o0Ny7S/R0PqXqCTmsT3y+fA6El1/fN7iQiZE1I+UNAdChvDVHnziy5P8emkGsDMa
Gxc70yHH63x5ubM5AglznGDdrt15xy/KCUBJnO5omc7/+aat62VbS/uP+ZNM4kX8
fk6tqJlcONsaqX0ezmwootDKG7BhA0mwddC7ZzofuGd9+EJ96/YIo3w076n6+X6c
N75LFmB4LcYE46O5xbM7BV/Y5PjU413WzbZ7smwv2qKFA+qDHyIlsNkdr4w0MKsw
VB3V8FM2q+G9RdtfXymH/P2aJDwU5ZQpcL7qlw9cb3cffBkQNBWTcOGSHIfGPaIF
3n9UDan7kMhVTb5Pm9nOnC8FXiAJQv2gtrTt+kggpYD5NVQ0BWMf+nllXqZoXm2I
P8wJeuDhR4vAp7su9CQt4+zveYN0zgZQ+BaT9od4UDSF/4+0GJOJrHYmfGmYCYAx
nP/TkCW0etX7QzQ5jiCpivHlbVHbKteLn9Ac0ypIw56gfLqapzgLspLX6CqdTVW2
d+hvyZf1OdMtY4k8NH3wgfY1mywiczCdJtaST+VxbC92sFBqENnDUuQwJbEFUnr4
RMHR5TxTfE/KHrk8m83JueY1Qy3Ly1WCUUCzaxWCoXE+H2wbCNQqi39QManeMN5U
29B4qdLw3rN3VBbqwotH0cuULlJF+jtYnGZQoAwAOhANsVaeq/JDUbOgyPMgknWI
c2Obhrhn6+LO8ubwjpMY0UzadYkX+0RUDjYJvI6Aa3Hw86pj8/DVdLkxqu5iia7q
ODF0Y3wePW+ynoA/FzuaT3X1SwDg0oMQOJOUEsdMGMgjGIJwE9sSsCd6GKWpvjIf
1erEqNtblqQ4AXgc654U9V1AOwGzl9jEID9YPnsGLPAPNS/LRRNDpGJlUdSZ+oFT
rJFtAUhy1hN80WldFLaFgfaBqEdDcAcuvxu2nTxxDGXMGopFBUqJhLOOfETaaJ9K
aGCmusfJ55O3jOlw5LOSnHONIUt79/tpRs7l7Uf0uxa3iRw+VRHg/m2sYNIUit2E
FWxsSdbQGTUTrU1xtclZc/CeYHP+xadThoDyoCoftpv/Kgfm38F4Gm5eDYk02Jao
mkihPp5iGFjYBybGE6zDRNZzxkxHyK9KIOvposOfsM3p04w9cs99zcT4mtqeDcpT
fskZOby0BDXaMu5qrwFYp7BYi+gYDgl73AbxhZ2CoE2zAUz0XKTzyWtob45fETSH
9COGfcCtnMW4947sLm1HK4A7ShunWivVJHmFFY91No9PTYYDZRa/yiYKPd8Ng5Cf
neCgptiScAAATkZE3fWQ8yaFZKlJuWa8YPZAWgGJvrHfSWqHf+w/9E314FFPRKEu
F/YIqRaSm5m68uz3v3BgGZqchVM0vIbdvyvhaQF3c5tftuBx+19H/k+5bEG5D+0X
tmIRwpEkIIYqPW40dqq3n86KUJbhp86wWdRLfEZAoLReT27ZjHu/U4Np2K/0bscp
P+M5E0oY1eC9ZVeCHg3rLB6MpubbYtETjovDFiZk8veoy0KzvNATkDHAeIE6eZJ5
+d+4Y4dDwX/g0v9Xv6v6s3rtrqp/iuSO3tZVE/qXjR11ywzAM85aB51bUhu+gCgA
jtjC+6BlePtc4e/HkLWgc/Lg4GbYzknaD66sXl+7WRY/EsJssHeNGyA4nr7s2Dhg
++L/gd4G+7u9qegPdGkwXsOkzy2VJ1yiNnxLC0ZEogsyRuG4Ube5Zzf9NeTZ/CXU
3qscX/ZEoqQgesBv2NFUDD7GfRebteSmsVuCIBjgJvPUCwWyXDO2YpQRZQ2ea6rC
nFafqz1JIqAGoRuOpXLkuzW+CYBGH8wjHWfYPyfOiaw0FIytryepUriEY3c7Xx6Y
1QgWHCZOJle9cZ1SI0Rp858Tt7JR6WWMyWRKkawFfsTps+UcThATsp2iQN/EWmkC
RYXhFTWEMX3hWT838WroUNDr78AQhn1RqkQvJyLKrEb1tDuNV8cfAqC1ykEGnA3C
Lh3qoowtfMuLfOpbg5TmdXPQkbQAyvgdrLcWdFhq8lAmuvoNI1RHj0twh0gSJ5Q2
XHLDubF5qzg2kMvmBNvJZF7+dj8VZF8bk5w7Tpf8OAmuUn4eFrNHlUzMOWpL7E3n
O0H+zM6btZWqOoPjf5O8cUjmN7NPw7rbLZh6q5t/m3oTnbcGz+Lg7auzmhpayQKO
achH/PgsZ23lzNIb1D+DO0oD7cV6EdMfen2CZTPx7wsjymNNZ+9Zgbfq0/DjsA6u
NNYSRwdU6Vi3k5/Z+0Exh5CWHB18zX2mwC7dcGOzGAsip5UoFTJLJ31TGTrs0TVJ
KocjixMNSvs/TTB7UItMJUsWr0GtbW6NjXncQ4DuUvsB9Sw4QpBRdI9ZFTu1JzSA
v96dFWkkSqms2JR0vBqTTXt/9CxalqdSj+encgLwihNY3pTSNgCxjZwPTNRtdn5u
sxxueFrhIHBv4OiquBrzKyjnmjMo0bxP+0WVCaaY+gcweiAN7gPzq7DrX5fO/kB8
GZ2SddwWioL/8rejfwOedIEV8RFwGDn1HaiSrMm2kzkdgRaF5Cx14TL7w0TkXfwW
1R5d0PBQU4QjfL3WsgGfhHfK8VsNpl55dlthUjh3CdRVgIafTK1AhzNCdCPQZC9m
fJlRaPFl5+0wh1Xbrl4J0je8AM1FGcF9hSw3RphgwzKRXJWnS/xHh93dq2sCCHgD
nYeZ+iz/LY3yazHxlCXsVPaeFUMbbhGLhqes6qqQZwqs/fVbpC+cwODJ8JdHlVoi
6fAequc80d6FLhWnhMPsDgZkOCTjPR8zLi0ZbXmZSXk3gPgZBT/eAOU6V7yk05sF
ndGohSLMHZwwDXWzh+rsGDCO4tasz8ejczo+tiizWNs861LCKXsxr/+sLEH7rxuy
nZXm6yDx/vz0ShSOC7TwU90nmJCY9dtwyaxc50Vja5NjxQdXk0mq0Vg/K3n9CcFn
FRv8WXoc5NJY44M1AMnUZJ7hMY2EC4gR6OAWql7s5OkE9/2sAkD9Tue+QFjypShq
na0mkr0wpKBDb+OMfxKTJU7iAGCIIE7A7oTxDycD8PmYrCE43R2DzZ0Zz29eZps6
9Gs3iFzIB5wNcA5E8oyV23SgkpVwISP5vgX4TCg1MgUd83ZRS3eF3Ng/C3KJsVbw
PgSEC2riqGLPFQzJLQmoE5VzipceDJNjSkBdG74LmMMMC/yPVJ8VJM9eBGNOSMY/
WNYK/fwhNWIf8oI7XmiwzEHi9vGy35X5ecCkZStL7N3EYYEHUqQBoZP/Mqt7fKFp
w5I0pgVhxCn4qevbO+70ctB9PFvqVnR0UiN1uISKEkssjz4UYVugiNE65ZEHlfaf
yl+sg04+Vvbchh0wRD2TUxpM0TboAoUHN8P8He226jRl5NkpKI0eEWAtcVl0Jyg1
I+VSVo/YuoZaykKF9sQNleQSD/8kewNaN4xNTUZa/9nQapbQy7KCcjscBdj3jWHi
YhbJhAI0hosNY1/2V+YG07zJ4OgUgHEEgY3vIa94IGaOvp+mZkal0Gd7vRMRNHmz
BkDrxk2McSVAMUwhaorAIggq44sNE6NNtpmlcydLg1JeKLZ/6vUOtqPr77wgPMBT
zdbliWOGkxn1XtKymbgdTlUtEZ2Eh50OPaDrpww4f2YQP9px4NcOuQpIA/wBUmm6
6sY7CGwfQh2UtFQ0kbKF8Q72hYiAcXdAxD8pOR/DBWKXZwYpokXw89A6RWZ8jT+G
gQfYpbi2wPMbCaRMwsuhkNnBMhBlSTEySygfIDLdkZwbR1Nt6ByC98XqCBaq6GFH
o6+wv3bt2EPfS0RGt+neiEZWXbkmBxopSeUHDKNuXdidwYhgbg5xPITN83sSFG3B
VmM84BnM8SFMXVc9Zohq4JY1vNbLykIKQ8o/nJ+FmfhPTNrx1n1HpCrVZmfeaZkp
B3cxawvk64J8o2rkitJwNBuqLn3WQDcLLhFM2NP5G3f8tISlO4gNINuI83EgV7sR
kgM4e4mx4IOEGltUmKdPeL1aLGXegPte9JL025EtSBldfdD1lyO3quWnSUuARTux
ZQdfqw6J5upCUtqmOIqepqTCeve5YTFEj0uh7XNEJeil2tt2hd05t5bHxlptGek6
lwe3tBDueRUF4KWEuTVRTRQmXcuHTh50/8rfzb51ASWTvO9iouMdlaxFrw4viEd7
RPRmpXTKSxRz+jtwHlBf4eZCnPSNCaocL03ST2q5GYIPwJSQBMR3V4w5Ag4pZApY
fdtJ2y5QnEVquJznI3OybPBA70apwMVWUxA5JITaRL5rcUQ+xFvDwl925ahwyeLi
27iU1yuwm5SJH8cz8uucLMOhYjE6mNHbh8Cq5CpAnURImair26JIhu4rrjDTblOJ
Y1r9Gaz/df5d63t0LVX/Dqaz0/NzEDHmgTN4gVk5zOg5gSpvoCgZhaUNMo606ah4
e69XDFURz7kvesVAnZ1Fmy0jEpMlCqdhpG6w0P7Si6NaVi6wd5PxlnPicVBixMsK
i451RnShQ5GAMSSr7baSdkXyjyEJfO/+9RYQf/RKty6XbM/Pz7ZnywsHvFHvk+wY
pv3VmM1Qf+SMa3Sln+MMYOrMvafURB/kPSD0wbXDdC9y0zpNN5KS8imuIl5eu0Z/
1iRXyNOXp8384crfqZY1QZuyoOAmNAm3A06MyCGy2PgdWw2FNnM23GbqhRqdgskl
KeFpPrLnvzL/Ri5DB0a1KpbD38/ScbMGV5smJZTMw//uejM9StAIgygr2uwE/Uxx
KUb018uSaz1kDGID9f4FGOuB2yq/++4OnhzoiyG/h2BXvOR7AH2OwIOrKGigfwOr
2+3222WHE+kUL8Dg9tPejKAGB2csEysLq31xuMu6336XGLvvZkZu9C8B37Pk5L0L
S0k5BvFf9KA9a5Sg8wVIrS/hLFCralWIsY3884iLWym8lUh5lVtAzaEtf7Y34OqY
LkgVmd9ny+PwMleRoI8CK8IuHE7IgkphndCe+e/OGvDQGr9q8lf6rG+7YINGuJkw
idcXB64ZLqzxC2b1uIF7GbGvAV4JZl3xUdJE+VLKw/JMZUsrq4pTBKZdqQ1WldQt
G7SVmN5r6cIUYSWbztn6dA1f4dtmiTbT1Ai1lFQGUX75kqveJpKClJj/xZtPo4eU
RyP8npd5WwkAubu+BWwJxp49500bRoYB6rQBX0moBpZH09KxKfKVVtgflareiqMx
IeX8UUMK2bpXxcUAbxHEx0Z1U5ZOOE1d+aZpFPbqS8gzww6daYoqisoCzpQayg6+
fNKpmNvOMgvZ8C6bIpgbZmBXAEVaO2bpjp61TfMwm66zlF6FDj6Vm9U3Hq0FvKUr
qYSJbcBqtH+ZEQBVySwWEzcuDUE0fe6OY0/fizxZRRQkKRCU4fjLLbsV17Wbkb7g
SrrVNz/tDa1680+1L2bNUYRVGPHOVRmDr9UvGUv7wvtd+LVQQeqyI4OpbpLocB1W
TbBh2NI8oQs89+zhOeCSGpCwJN/KpKshE7gB5Spd88Ow+76whn9VuM5zZKMYP/Sl
0ofW53M5ijhQruVCNdiZ9Dr5bLtldyKcUiOA76Ps0hpN5wiadK6dqZ+oE3KbYimH
GaF6MWiROshGS11cRjRFCcVjvT8TIaDALGanLbKx3G0VWWT+sV6DvM5H3ETJ7Ljj
UKzIymkxINjGlV4lIwWNT6ZcQn/oayB3s8g9GcCbQ0zV6Da1bwoL6unY9LEJNWKi
Q8H4CwxjeTpy5SOC/6otC+N4cJ3qf/PG5sdGmYgruVkk1iBI7aybyRGaFZ1jXHZf
vv9wnrrUKsMdtQk8NrZQNNgB9U5I2+vQN7xama7+FsgMPe5pnbm2Or1ZeAIqc+8m
IZUu+krGS/xPYWBas6fRjr20k4+1xQNQVk4RmYxzOVgCmmer/aIqqOxVn/ZPdtSX
zT6UKM5SMSXdHauM5UvU2XnroHIOjWnjPsoD71GzDwQNK4hj5HhrADQGeJacxQtt
t/GB7uzsurrsWXww4Li4ITOjVNF5JIt0Vp4GZDKtvIkIntJrg/RRbzpcL4aUfVry
bcVuZX97/+iz24lzeAhlE4JKZ3P9keBZhaY1WSf4bLsJr2P7FbrspVjuzTK8Cz/Q
ETR44vJxAtCxW6QOy3WKFkHeT5wDFFPHM3ABFT90i9jG1wa91YbD0hnAEpiDTx3i
py7xoRevIuGxfGxqqU3hlNDN1ZuGQbrikwChYOXrGo9HLkx2GdfOenF0a44CYVOO
pbEe7yCxKhpyz2x8ijyJp+/ky4GjLHkV3UbqRpTSaPb3vqOBXhBDSnnXQjbx49WF
Q+VieIQa2xO8x0pZofeoEoBol9vPyG9/1rNNZjqbK3ge2EyoetJJruahVlHYLtR8
LSQMIse2kgFFFEeaTjGvUPnKTF0YWNxh/UGcLhghePucGrK4JICDgDxxyYV9a92T
q+GVFgcl4dh4YvJxvByRLBTmdO9UasWa3GpKvqQhvPhCXwmsIYE+fZLXDP3VF+Ob
5JGqOm62oBr5IKraB8mgXew+LAtsqxeRMf6JcIenHW+ObvDB92C6POdR4l9lC925
QQf1Ft6Mr+5jiHekHbPCiJ7ml9T0dQj7p2XQ16gAL4KSV4cA/VGBlp521hTsv15t
SHuM2l+udg8Ho73YN3cKOnRqNRFrkQY5PcrYjvoMmBdzaN/HopPYwjW3xR+rNjN9
H6silhpfuwa2F9Pn+S/QjZIdGJVWgQj8dm+KqlRzqpBZgkzNu1obnUwpb6rSbBHn
u6OAyYPtwuRYgBJLAcCX16ziWXtB3/JJNLi+7XL9wDSqsQ/AM0q9D+wS1KWC7aDM
ELj5yVVBhJEVfO6avezjFSb5r5xSaUkJYZKP7ZShhze2B2brIwIRZAZ3ktfRvV5u
8F5F+6a+sOqYX73pWr2zdNBl0rJj5Yzz6RaCQ2yisUf4fh8wF6KNuUZSs0kVEwVK
h4eKa5o7r+eGggOaj2dhc0A+5prawjWYHKIXBnW9I+ATSmZBHGIVBm1/W28XWlZU
vKhrCuGV2BOKx22Gyfuhj6OmkmbDgoPyU2GMhss0ub8kKiupzSTBxW2cgSK+orHW
zBASS5D7oCVYx38AF8wEqfjkF4JBdZcyjnUplnS22GceinsnF2OhbSEk18rrr5oA
2tsq2Q5Y94pEG9iHwC6yxPx9PqfP8ec3/qscYe8biWneMstWX7zJrBneTq3VIvO8
nAUtFVC2nopvBA6G6vDv9ItBfn7Z7J5CFULX7qI+F91H1BD01y+RMXeky5rWD2aC
inUI/G1VyTTBv9UGqtcqiksHNWwJKNYdqJhEgdRK8dISwKIvIIc87Q/QltA5SWNM
H/x63B3E7tY9U6+gq9wrVSNaFiGKGmkDriYACyJeVv03GLv6guIt3miGfG84CKXX
JC2vNawcyIkTA7sd+6t9IGYtdtYNBF64hODiukEg2SgPoHBp0EI9o2eu9THDOnUC
VDSzMF4PIR7hiXTXOINjUez8RWHFN9hhlHnKHuA1OnX51k5fQeSphyPN0596mXdP
kSMWL274MqB/VzNGNFds4FEO5vMxfrVTn/9nD7K6XW8WYOv7S+xHxv5BeA7RDqV5
yLIdB9O3/BlNKfADMJsE87aT/bxnN/YJ7YRD7xLG/109Y+cSkSH+Wgcwdmi8tIzG
onor63Kdbc1UrfoWXdDfaeU0V+ahAV2q/ScokOCZB1/mWtrcngTBXvkOSWssTGnS
0hac9Dq4VTd+qu3YWLIl+ay8Wy7853H9w+eOnTrdC7ymlk+U2ELjZusYLSTPayKF
PCaad38b2xvOhj0RkCAf7Iob+XlfGeFigWHU11d7doH0gVI+q/KalSDZdrnxHB1j
NwbCbf3GeYfPAQCd2vQMWXsAf1kdWAbqS1p2WmlLqvz3YEhrK7pt7DYSCgY6b4dO
kELEOOO2HXquTZ3pqciBKaS6IOO+/wP3S+knqFVWRlXy9u4Chl2YcvhgMuN9cOfp
ayo2YjPjYgh4FuhBMjk0CiUtZ7DUl8DpZv0bu5QFKdykQ3rhYlgD0rzcaDHvBtgf
8R4NNbGJk8WUea0Par7sbiHw35uxc3xsmLA635xSBj0Fa36+wYd6df8HYVz4y4LS
EAnbu9AkfJfdfvtX3tPNsd4+NE9UWWt8360dyml4ENS2Hn56Gr00YgaG9ZXsfUxL
WHvN3Pnb9zklQUXvN5yBzMJrVXXHYJzF9Y+rPn3lP3hHkAlURKb7vzt1HeKaLLhh
C16RAbY9T0Duyn0iuE3AQh6CKx3AI6DsBiGLx+MVtCYLBjczauSo9yiM2HFYcVPg
4ZNRj7V2TZYOw7VZkebyzjbmObQSy/ip5/bPeDJjKEDs/iTOph3z/rkzofbQAZgg
1t5xww3fgBY13pTlteowqShQRAT4MNq8is5FOUtwyKZwrXD6NG8MO6G6D8JXnrl7
AWT+43PF+FHB3Lx1WhO8EOKiSvk8qcBXAOzpPKdCX8MvPlmXBJKCyV9JFd20pmre
rFtr1z3HU+Jzvq9uSTVOkJ5NcbhOIa+EzWpfOhvec3/JhM7pS6qWKup8Kjy3emWM
Av/O8rSFSyzZvvTDBXgx9qNOk3qYZSPz45Kk+QlfcEL8f+mMvPtXBj+AgC8zggnt
n5hqRTMHAcCBHecnUzPUZQ95twKD6i31FzCQ76VfAGXy8bqVQUoyyXe6SfTWAUjt
yuHSJg6ILfpMr0knmmxVOj6fC7cRf7VPiLaafgvucOrqcHeaI/1xInQRDJc7Xxit
r1C/il3MdMQ7SaGnZ+TZUiH2AuqpJjzAIBY+lDXkMnPOvWqlWek1M9aTRR/9nilo
xl8koFCO4JLZpNuq43zvRmM0d2S9xh8kaay1B9nbDWKnnCaR5YVKR1kTbiwPmeEA
uiRlfDVhRsbq+flsw8FseZbDLLIz1RK3HFAKs+xhMFdIIoLSNrF9TC7Yz+yE5XXn
o5pOGPmntXo2onLjcbulLxhjMbjd0DrprQ5xc5fy+X289D94kzlK5MhIKEJtjggB
hdskExfFsGtpAn91N7A1QIuLwXn8AVTY5FusuB/b7vBq6JHGorqDxgJdGyfjZgSj
PiqysQ4lDR0/PeEQpMbovUlgBqb8Lv6/aOinKmFyeAWt0Tb9QjH/BBUc63mRC5RV
+LePSdiwe5tqQ0KJPbI+CH+hiMKhpcjqDpaN0e6LWtNjuT99QjoRDsYQanBtyvxB
JS9Q2vpZbbm4d9JG/EXOvBxJIpbZJYz5GpB5HPFcRX9oLky1SZaznGfLesc1Y1AB
QcwZ34J7dqgvzaoZMyXMACNRAVf0ON8aIskrLBuD19UrGBBnT8Zv6f6MlA6AP7dU
/onY1WP8B6NrRXXnfihh4iEgvu21l5wEsYmraR1Ao6w8/zDu7BHUcX6OGNK0PN1/
bdCTll9idWjASGKDR0i9rBfEwjulZMQDCoyjHIJFTGyN1FafMETHV/WERHtu7uXx
zE/xqIP0aZmDlq2TEMhtTJam7eP/iQsdd1e3LPCq3N+XnFj6V7KOZKNC2lC1/Cjq
SIBjYbXKY+wXtxiZQN0Inyqi54NLkcXLidVPD4UmdoptcPmq01zDApl6cz9lHJPp
Llmq0T1bcQD6Cy8fMuINNL3qhMSilsctM4LnGqDyih9Pbd63CgDtI60nhQcVQp0f
+Rkvco8Xad9FV5N9dTyL5tPqMUxp1zUxEzs83AMSWB3GStIxpQYTufnnf7BklZiV
1n4g+HqtOoYjkGCgtdhPC4BiuMAzcTk0hmqE4ROtxaoc+/+3aOIV6g+hhrC5bZz8
R6YJnQ71uxT/NEQmaseD9OVTyPLXD1XvRiHr2PIOA/XbhzQ5CR+0htxTe3AJCF2G
Fp0gukQolKKo1mSjEU7MS27wGuM2u3wJQsssXIewaTKD7R5t3xC1Gfum/M9GjF8T
ibzmCFtWVOXlZF4c52u4yBmsJjA+DLjmOmcghGIiA8fLLLWXb74LPWg13LYHIK/n
Sn4gG66j9ygwoVXoAEAeMPdVKfOqTZQz3ipBRf2bS23jhFoYmUesGq35I2IRvAm3
jCeFpqv6Y/4y/K+bOldKLWmMby5jHHTZblWp8SkSqRcfqvKp/4luM/WH/TvqlYpg
cXjkLXKtSn3BC3clUnflRVN0MCOogGViBbhKJdjxqsflNnbGrF09YduaDuFYJ+fw
9PxUPq6Ol20Kj5xihzDAFIfWMhRvxW1/1m+va2YcavKlL+EFC3SJagYybaPIA2Tg
pQopcYJSNCSAi7HD0aAkvgNNMA2Hx9/jImgLhbk1h14+ES2agMUMFfyoCvnXmMvf
rj8NriIwIMAn6BHm2S5b+cBIIkGjhrCbaWAHsCugJxjUU46Oj+kuVVjENmSqUoes
Sl9SVDIVkaoHS0OkdWR9wwDxWjSeqkHTy5HUM4AyU4pvix7Y+ea026HAFBwK/t8y
BuxXM1pHqGHcdyQVe17SABqnbHDlrjZNtuhsLtkTp3FR0K+/+4832CSOrFxVRd8p
FsYWFmnrd2Fg13WUnEqT8+vHDNyXr8MwgpsonCceGy9Y1nP7IeUfFS6P/dzVYmJr
avitPtYD3KHilH+joJci4MTPZBqa8rRR/5UyTWZTTC5VgdQIWHHD1FLLRr091uRZ
QGodBprvDQ4SmpfLQzX0S/eAiskD5ZNVS9dNhcXp5VufS3h1IBlgULbFGhaufYG3
eMtGQFNYi+IB5hilrz0WnPKCmRrVW7Lk0t9CfjIELDPuqsJILqX4N/h4BV71mRM9
atGbfqRlyepVR30tT46/R4TES2bcPgMB957vLQoaOpvJUSnrc+XgW+QtLNQxagpR
u3RspmwR/84+lK8f+EsXTMY099l5q9iLy5yoyPfb5wgotKGG62HDpWvB3tapaOa/
lV1khtTeGKNvHwlFTr5pmAxNIJGpyegAylNWI/LlBi6QCN9l5cDMveaUpTGagDiA
6SkqpJm7E9PJR8WKZUPqj6yeZl228s+jGGxgdgGCBjboOWqCir04AdBPUjZfeqHT
/rpaQjcSyhBLuNufC7ReSQKGWSnH109dZIcZinMUcNKxY7jRvnI4vyM4feG5H4mr
akcZbwvZK/lDo8OhLmKHwGsAvtqRA/QsxcOChJazCWEmV5MUobQ+SS3eOJxY9ZRU
kcjaeg0o7V7OvX8VuiSac5icGtBvAouOvQy7xva/SRJGE/3/vF9cunC5A3zwLksO
eELTqbEplC1/APJjpQJAIBFKihjO64Pe1LbiCL3j2+xEI0DmlisLBZEGTerYP2X0
3Tkal02C6olXEvKCu/5rp0DugzhS6Y5TohpAQkaXs9btif/Sls2VOtQqygyPoIjB
J5zjxXgTLmh9/83E1zhvSniMUEL6FzMj3lM+H1w3yo838eUjC+ZmchXK8viaCJhQ
hljgfcKnpSiGPQ96s21IQLa60eiyIjGnY+fMC6CPs9QIa6weWt48cElfYQg4UX7Z
RuQI6fl4iU+8YJEAzXd8BamSbJ7IUrjLZBY0r22gkHY/rtBpHEztZX73/9OERNhx
imS0jfZuCKyoVvv7VMie4xASl0Sx0P/60S2kHPkabT6WFpQEvSVpKnJR+GmZSY8S
r4kjTWURHNqnROKI0fAot+Paf1zZ822a8T04TdE3+IZ0xczlXwv/7PJbehUV3yCA
veIewYiSiTYJmBapSqvP9+3P6yCjMrTc9cO4L4IF5dz+suUQsa9xX2lM2mbKI5dz
/pJgQ9lwjPmfgu3t4szWBwAnhMK9bZfHVCy11HQy2mbaIuJvCBeJCRTXmiRfbQO7
1r9aakET+r8HAHv1JA/DGKjavi7f6IE3MWd9shaPr1Q4Jg14KirBjiaeFj0Zdibs
eYeHM5pZUmC2Qwb1vHWS8LVSnntc5la0yDt3bc0IoHiuYT6TjgAiBStnKEsOD/TM
Upt0Ebtq/fPKvERzhcai9GPlN7dpZbcxvI3nHYTYQweSgqH1DIyXNkDOKpNMOAyD
fgMTKgMnHFjFP+ay0Ow76X9tQvm1MRMlDJg1vQK4uXXOPnN7fq7VdTfNDVk+otXO
rtaw5afgLqOdaVuDyfXCGxzhf55gV/a3ZWhOfNi+ZGYYan0RuqvxxCM8uMic5hp9
7KadcWl5RDVR5hdsRY61KmFSur0VzmwJXobkIT+mc+VSCdLHkSeNF5VgTAtOKd4E
AFLS6hXAHlZ45H98QeUfh6pUMegDfJVKoorvd6kY2rySVoMqPqttoXw0TsoWGDuU
4BdeWVxqOZFvMf6+SNX146RBKNHDskS27k0fzsWDjo2KRLo87bKkHzvP5pWGqZe9
UCaIaFhoedIrYEjhrZks2VKzropUu3t6utLT3/4U1QqFOPM0nBZj9xagH9HzTt1f
oeEWBroK+BDtrlMlaSNyE1cDcFO92eCNpPbObhOM33oGC8+UGCQaEixYt6bmjizk
RsMFGSNMMSJ/WJkwAGtOHj/Xgi9vvV+msDSWbT2LhRh4kTLSCNoedMwpJVLR9orS
hZleKLsk7bWQX7dvgVZfJ9I7ntCn2y7AWYMyIKC9oUfu4wX1yuhr/LJEXhEyXkPc
QQXCeJlhDX6VtMVN702A3TK2Ftwu5SvXba2UcWpfwbvQtab81mLXA4Zx2zNhsXN5
Wgn/FvGv+VMoIcEyOV+ApMsMODk7itmMUEyAoP12iLkQWChT2bU5kDRXbjAErb2z
3AfBOHAHT4AxJf5R0T65DmtNUdnU9wywFMEFIDGXBZeBLNWS0wrmaFnbRwLnCBfE
5EItQsiyzyK4j7ZV7lJVX/2NSE8giR+i3avqA9FxlJZkoztITiwXlSR58XEsKvGb
TRuTyJcRLEu/6a9joxanARBbb+bZfdNfbhVumm40yW+B3gFp3TEd2Ly+EyIeH+pv
DH1qx9TkAf/9TAdphtAC01lL4E4h0OkSDNuNEeiyInX31jn/BrHbf/cyXfMFmIfY
64bLYT8+Fz69SttjjT9c1uAPpDemITk7O2tOktMCOW9QftLJi0/+eVEduElc1M2g
5OFVAjzeuHhFGgPO5IUxj6J/jKllz5JL0vnUelVgMYbGliMFe7tOhIuVzR6z5Zdg
KwozB2sG5lAAo2zcCnD9yVq5AAjGnKDNdV0NxwZLY72rFhTnm7GZ5Khs7wgbCgDt
IAKHz0s6c2EdYCN5Z+ONq+Qbc54V4BYZK9Mm/GVc/cWWNPIBwbJ54ujSOmYS5XpF
7w/UWIdzSJ7aO037cnvRFwzRfOIPiDJOpG6MMVnZuabCzLrTu6x22AQkJ5nmLeOo
dLufRyF7bIubFCtQFpklChWD3OubhTCu9iG9LHVLSs++F/5/ZTK9k7SR5TZF2Jm3
PoW7xF0+4y0MtOSad+j4CdapjIu2IA655ABw93wBT+gM2L7SNhlioWMzs83n5WAH
yuI/4+7nTxRZTahir5Q6FGHz++LYYx5DoU6o9QZqWaMW3iNL5PGextSqWS4ycKmb
QK9c8mCBq8bU9Ewu3HCLbNcV3C1etgBxywaHpBGlHXSKr9hTosIU7xxYRPT+ndfl
bNxy3EiWPrDVGRWildWVUbWA0jqbTRzwQWYOiyC0F/b1cCXs8CU7yv0yMDpBkUP+
kEmB5LPwmGG8PASgH/XK3AcGh9jULTh5Q7xU2o5NrUgF21o5pWiUHdhdUP4ivJQ3
o5kxxb3LgzGxMYSP03TUPx8SZhGcUDEW5+kM/yyukobRE7Kq4YDnXjU6NFMDY47z
/UhKsVXhllxYbXi+VWsNt5M3s4Y2I4ySu6zo6p8waDwNRk3q0guPwmldaAxcugd6
aBQ+QRe2XZuuUOiuCKsYS98HgUTmMik/DLH3yBQI3MKB/yw7wdhd0BJmWOblhVHH
0i+t/ThkkOaKQ/8Z+Bk0Qhq1PwRKYCA0JX9fz70aej6rWmMbvqSEKdOXqZkfkKrF
xqimn4Q72ybJSUZWMTeqPrLVlX/DQeVR3srrllVtYf2Uiqsts5xH3RMhm8oN6ao8
D68sceVsM+RfZ48UbUWVCpV+FgC+i/VhCGT0jCxDpKH2d7YV07U5qqmA4DEknEi2
0tZwUYirkumNS1TC/00ldxHWf3cqkwZ5O6Z8dRRmRDbsbZ2vDCcPpkwFTdpVcFWx
vLKrDYiLEMHTRzp5kz6iaLR/h3pPAlrMcYFHEot0P80gr2Jggal5KU6ErsQHWLPX
kkmHrsPJaZT0S3k80AsX4sxTE+yDUSGrkmmYnrjeUA4dlJ+iJE7zaf8s2SC0aloc
5yy6BMH9lZAtncZc47yvUxr7DJNPtBO97PY1wn7U58WIk8aC5dHxeKuFG/GcKuY2
NI9BHXnNtVVRw3vG0m0kmZje+m7waiK3vvVSNuHh7I8heuPTqSY7Ql4A6pSKJWcX
QXNclRodXQcVNy6Xe7ezalUe9kwl9z9U5KjjacoRnFlSQYIbJPdfJz5kaDJmA7V9
Wa09hTLwZL6P33pDC/Ucr4lsBOH3ZIJHtTQpdJZ+j1KuHMxh9+1t/ABv353lcTVl
fgAvgOtTZA9QXHQkGudY75+VbMzPBso5+hyOZvh5putWx798M46iw+H4jx7j4IGq
/ZWfnRpk/Xut1Cfuu6SAED9eBeIB3zJ1c2Kq5E/SK3IAl71LtXsxMt/93drX3KLn
/y4bgv3SWXL+KErIXqA7ySp8nZbRRIXp0IPA7LmbztB/7awu9RIv5mgqFTlBtlAo
G6ZkbdLJ3xJZP5FTctIFzbRxnMTjI149KX/68Zm5pjMSM2QBOpFttOCQyofvZgVd
HzTdKYVLg5abgwDnD+c6UQ/15/EqtS51nNUeWiWxdm8gmqDd9DHDUHtoiBbbwQtq
uIUF68k2XCMfaI0RaCdrbRwAvJyL894rtjArb0dZLEJnk0jX9wzSe8diPg1GVmg1
GTBy5OM+aajwtc7jOOsX8D6yfCmvOEnRInTrOc3LM/UGADqntmlN2HIrUJrN5S/H
0Lq14mZPlUOF5HOINqPcj67pQQyj+UchL5SmxIyGXWE+Gucf77ogEgyZvmt69fi5
S2VmKcIBWL5HVoDb47mHcdyk8vsA5W2LUnjrDt3ahxAIsn8ZNQYU208C/kpcb91B
MFNIisu/OwyS+NgNjLhktW3tNpNXdDz9NSAIvDeXAByqFik/ZAGx8Dv91VhwxJap
kuwFTUmtKo94kSGs+P0zWUs+lYjoOQhqDg9/Kf0qVTkZlhjAsVF3rJQHo9Z8WqVl
DLipO/PQkdHnKmALkNtYGjrh99ElszuMhfVNFM6eWIKq9vsD9mBOBObW7sEmw6sm
qax2frx0F3vTmbifyFVhys5gEh3MO3e/C0P9y4ewr1SBNijVFDYywIMSRzRwmFVx
fpa3q39+UuN/MdDMaEUS25pWa1BWzvEDGn1StY/qNFtkIVUWJ8cSWGFNAmTqd59+
CoVr8+x0lcaU4ACWeMk5v5psEZwTdrIh4GpvXKOctMg3vyO65litD0PsY9XAOYw6
u9YZi7xNMq+PqAz+OU+gzd9wbFLaiuR0M+J0tyLCjcG5G5Bc8N2qE+1si0NqudyR
+LPR1EHF2sAgpwyKFk+NAd4xOB04/Fx6A/FOWGb0E8rAOlgqzPJRe7UnJ8pDTy0x
g0VEq5V+WcmSpBmnsGoPI/cIjsMOUSpJ1czysDKdUuX7v2G6OFMMZ481FRD9KCqf
4MzJ1y7QfW+OgFAN7WnhZwKgQEbmJoUGOTsS/ovwMw/fDRBEH6v3fWgH9gX32mzg
QIFpNnMEl0Bmvq2CkUHN6h3VdCneuKZWQp4lEcCrggZ6Mowak6ugXjkL6uxaWJ3y
Aoy15/IIr80pW0TY5sL0DkjlTYauIKEwkGt0UX/okY213zYctrVkhjcPuGt/kyX0
mX2oBHu9fSpW6GvlfDwLUn15TRSq+OxbErPHlGnF3KAvmvgTOD30eTEEB3JrUUnw
JqAgyJ5EpfKCkNn4T/ywGhdsfbVcqf84P7b0TZFmYlRL8puDw3iybaF9KLdG/akW
zgc0nPFeSjuq+R2s5yixPgIJqqD+hEIBDKFx6a5dS+RoZtmC1/RlzZUXujUTwtqv
xcpRqmJowkMbS9AGV3JGO1HDxwRdWBnjYh7WBK93DPywPJBAyIATdYGcJ24QLPYB
RlDrQShQrREE8kpM2qmuzqI9MZ+yVjIv2OswBrs4TaivQj6h7pCHZB4de7XKk4XI
Ib8ViwOg6SVGEX5inG7tJB8GEDTnw6g9NsYDAj/RiF6fnb6TWL4rdaLbWnnHjEwe
+4pYVRErD3/sAOTm0TM20IR1uQ9d3aJcJWywuZI7q+8iXaVNaD0mzm6Rnh9WrFIO
keV4WS81LCTgNzco5nPDftC5rnxdtmk+hIsan2eAb5MvLnormnvZARa07DQtOmHl
LvB3mbd4XNAUmPWkphmAmP3zwUX0FwHckT24ZH+4WTHIc7ROw2vBWQ2HOXOz9yj2
UyNApEDwdHB6wJNU/37uEED570683nOnIoldZwlEd+4brDRJqBusMj4DRlD1njM2
W7au5yhp29KqsLTnj6bC9YBUK31TVo16w9FHqTGDP6S04hcVmD8vxj0yMSLg+vYC
vBMELlobVAIsiVjpHDcNuZXkeAif30Ao2SZ/bU79xml4cA2H1Ur+3g/EqpoMXtVu
ZlLu+LRut24YOvGQjAh1ydHUnCM4uOLolAJZARtryLXvNT1A+6QpgERpypRJah3k
jBO9a4rfIEeIF0wutFjDosiN76YjvY8YhWGw8oTgNLl43D/ROZgHRlwXHckUTm+6
mOexmePW8PlTXgFv3e79Otcf8ellGVsu3OEwzW+CNW0d1kdOM6Guyh9yCbc23uq9
Zqp3wjVXZj/nlkC8glrQHpC8qk8Qa4ckRi4cFA6Xc6tTcYfUvLX5Ih2Jb9rkeT0h
A7m63CpDlPrn+X37ka1n4SvRTtHbtM7pjXokaWLhSTXyVfF69YH7w+Nq8Gg7L1Gx
AFBqteYp0844Jk7L7OOiXM32icnm0U+G9iGZ6Te5ECBzySOakyRaryXHEHual800
YYy1MBhnY9oKhQcRluwU9JKRxv9rsjQHjIZEqxLjKNAhYfx8Zo0qFjDZfeMX2xLp
FpMmrB8XzyPmbv4YwrUimhmUgdV6XNn8MEYtR3JqoqEibNIkIr2JZjCqq2Tu/UXg
l65717CZbuJDAqfojEL7i1+NwD1n4dfY6FTU0dwG3jdyOIu9Ef+FjDxegv0aCgot
haoNyVd8u5MacQtFWveYW9Al90Y4SDaW61PnKTrlzu4zy6/WgC5XrrIOzbqdiFvR
Xek6ZuJYa4ZIsnppKoQDLL38P88zt6BlR/vpOXUFyzoMFdQNp0qlGSnkxcAySB4f
sNmbGqHBMoSHHWJ6Ai4FHp2DjTvcSC32VTp1czcGmTZeoRU6RSdbYayVaZWv3HF6
3qDVZNIJXBnywLmWrpKI2nqJV+FWUvfQzXXuPc7wvZ86cmI+00Vtp/FMb2oMWmoS
kOUAr2M9frcx+UCKI8cA4tN4CshPCm+kMh0ceZGEwrdm8U8h5XsBdC2prlOrOcHL
93eo+9xHd5LHAbkYZDXEX5gZDt+7ge4tuX9C9YXNOZS55pbgknUdfOCePbwtMjHF
w5+7zg6DqF+7RDvx1GAVrRhlQ3kNB2sei9QSvnwjSjpJtAst+dFwcBXFhY0hspdZ
dfKDNiQ92+k5IjgjdVd7QaswGALNc/SRPCb1QN37MGZXNtFBYIEU7Gybx/5oVlvl
pH7f+4okjZCb85msDQ5TOctZtZAFFylR+myNU0eD81AF5KYt5gxI2/naoprjl7e1
gFa0EKyCFTxgeA1jb6Ud2lWPzPUu5f1hO2ofX4eVcABNlYBJBiBNZBVEgZJ9gdte
HtI5G6SgURTTZNZN7okvPNZb/9y5sWAzXxmQtPZX708ICmSPoQmQ8KViwOnVQJOU
P4cBJXclKjEHxyPQRleHe3KhT2ic9Rauf/ccKdKXjUmDVLlqltOoo/dbaW3sMScm
FmrPJtAw+9MWgmNCrgk2qQ5TxeJGwy7ZCqP87oJb1XI5L4nwuTzLEw6Ej1yRdXUv
X82vxWxllTVukur+epS4Q1MSWnjgwNsgl+0mrCQL7AxjgNpiUJrIItyiJIHOeo4c
MDrGNcevU6j0Ef2imxelv2aIXr5cyiz2yimbIJ53l7N0NBU0VlRn+cuxaL9c4GG7
d1cT62TQUGF8YIoTeN8N04D1+OYWu5xcSJ9sUyC7u7L79MIREPwcBLXbSjrWBrF3
s43icCmMoSJvcODFmKy/nZOsqAkVbc2whEtMyAlXIAdhzVM9f0yfVu4b4UfVQ3pb
GAhIgUSbeSwyFXMduSaVSjeK/2DMQt9QX+5xsmasHYZV5DHua2w7lizGExDh2rmA
jThTw42PLWv/K/Iw9R6M6ZfQ5Y7GRLHG5OR35QZSIIkg9UpPFektxyJqbBgEn5yZ
NKokqkfp2sdohscwT71MLal+CAIxnoiO/dd/uttRk5UQ6pEG55meUdKJgTfWoBBj
5RVozOFzjC0MO/pQacZo3yx2pnAGBLlwXTlUQZD0ZXD6nQMClDHTegCZJTZRqhkZ
/Lzuu785EQQnz87vIrjgMVtkEBYDCP0WrQfT3MIhijWt0CsUIoUd3L0T401Zthyh
AmWekYRb25PdsxA4nxPRP8zFRN+7zcL+pfBb0QrPQWI=
`pragma protect end_protected
