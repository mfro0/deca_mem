// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:45:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KT63H5m3n97UKytik9cZgkKTeQVFgeEz4fGz/CXDakcn8PyNI64y6JI6ug3us4zT
uw7r+87oIyWCruTDHp2dqKOo4VQohrJBXhspyQ7p9Yc/rf/2PRPEoEPvCkbjf83Z
qFMzxr+hB5FnnYI/oH6bWrnMhDjzo/xLccebjiv4d74=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
ImmztbpxobFYqqW+w0g06FutI/GtX4TGdNUY6Ts55C4VirCCjFQ9TA142pFtXSUs
LaQDsmjJ3ShQhZ5g6ckrIWYIhKGpOtRcwzkUYQzBEJucDHXRhL3U373iyB+Lr7o5
1jKRxDkYHdp4+D6W4cwBWhBPuuAWKfBW+4jd477Uc51ovtmlyKbxYK5UNmZ8/3ou
qpxXwxAkSLXYByrdYtbjQe9rS6DFXhHCU/iSzZ/VVKWtzyrkyh5fTQ5Rcgm7x3Vv
HeD7qDtxe5WDMokhMUXLWEoXrHaKbzL4FYruw8FRcUXSzreZfiUAlETSLGi6nVvm
Ty88p+Sn4hSHVyfWYoCAVD06g8DDAtsqdh3+0OJxCoRsqBvi8zfg9O3R/Vtlr51L
NWYEwN49xJgl2Lc+tWOe0Xb5IKprAfAtsXhcoZn3ImBeyFIWk3IWY/9Y0y2Y+beN
xzbiI/xNX7skqSgyhVT19Om+aZsQi5G7mSjUqbkBXEZ8v3CFU0x5U0MVGCr7HK1W
m9UDSUK9MIzICasMEhaoSF5Hxxjwj023yjzXQ4FommTGc/TQ9hz3nuwRSFezzIf7
fhiwko4g8tHMyfz6WBNhfGi+QImsh9/ZJKZMypoXH0n77rQm4x8pc1nmh2JVeuUw
McZ6GiEgtzjLp2MXDpe7uvhdm0z+qI1UohRy3AiesUCEee8ahEpCW/gwPVXjGAH5
N+EtsDmiv+UrAucDQ43U8VTZ+Sol6m+pAipEqm30uHhJCYuaoEfCietfi8/upInw
f9zuCr+x6jI4bMfQEzW82bN369mFcfURYRMfAnnxtTGdnLuD/BJR0oRNfUwPFbWQ
JLiiYx2aQinUHl2WVcg3ApQy198hFRIiM0VhNlNVAV4eTFNF7csRJ//FABu4yHUl
hYN4H4wIzXxPjeuWilvB+f8SMPtKMujAK4yXWrcn/Y6B6A1ZqWqDNu4V/C/6Wn6Z
Raka4WV4uXaUTXRWPjCUp1rrGZ9hPIFddrzFvaIRXZJbfBfLDY5vzWg4qdbq+l1e
/FRZD87U/V3x9PMHtH1qyGlQe3p+o7c7uaAsG1+v/Gq/c+aJwddQEWzzroSFv06C
f/0KRone8Ajgu2Os4mfVaim6vtKBhbkQ22nDdNz0KD1K5PvL5sIIckVmXtuwTHRy
1mhj2tiOm6G87SF+tauJQA4VW3eBUAc6sVpkJD4s4h4VhAnnX8LLMXuRCac6jiv8
34sQnmlQTgehRomN9G9llztb5jLS92LmhPLH7P0tzGg2J5Sy+dFqAaTEeWmoPXRF
JtJDzi7ZBkgfZLWZVNX6fAA8rs8ccdZ68rL+hX3FVw+MvX8tz2wSKC9vHxcDwSdD
M9Y4Kl9YYcYe2NdBzWj8A0r1HWuo2XtriSMWV6wGuOL0dTZnHd8Tq5uJt2wIkU0f
CB5DjwhIIJl0OOWBpoNtkE0TwfItTXJPdPIXvdt3qzVD4HjHRP4TJQRsXn9mwVkw
1bGkhuJiu6a7k81dyQ9oFdB5f///m+GFoBQ0KNV4WposfLDU8EEj/08o+xfz6cc1
t40PUMkP3XC+uKtPnfVx1GdpzxrtucZFY1O0iXKWkTgxOJ2PT2tVmU5LBYwDY1xF
3OcTzCpkqQUL0wlhU8z6aq2y+syeV0TJO1lxU+w1dQbMj1bblgfaMKA5F40xjm8H
XkdBUgalYMfJcDNMl95uCB1+WHA77nDs9o2ppiZ4uv1zO1Cm7XdJ67meJvRTYkhj
SJEmUTE5tRoyzS9SYq/mkEXO8+l2gb6zESFtblB4IV8M/XIWnKwsr7vMK4LjkU/G
nolv4tDdTh9e/xgtWT4KGEmp2+HApJDdzOdf0S2p0r2TzE+M8iHmErHl9/fFwsYT
opWjH2tURecakhRgCfayhkvfUy4B4en4FfmotJaXcuW7SrQpj6jRm7Jx+pYgsuiY
67Z06OJD1T7AWjb56p0XZLF1j3P63QNX3riwagaEnIaRQhUfdhwvszitmB4ZLf+7
W/Q4VDinKdZqAlGMflBtW+Cf77cMXw1t5uZy0Qp7M4U7/40v0toqfWuJgY1xfRQQ
4A/3LzhXRP5QiEkp1XZq9K0rDQATgnmh5vGPpJi18hq+7QJGqJHlpIF1K2sQ8W9W
JYXuUjQgB5Xkp+hCOGdQIFeUo61VVd02+HVCJT4RfBswhG+mrIZsdD6C+52zPKNq
8reLobuyMHXZhzwVVFX37oqJ0rdow+7ZzYXOqcxOzCCU19x6rolMAzkmgsvWLHiz
q1nTPnV2CXA0OtzGRV7mwj+OPyExX44qe6hDTtONnEhu0fteM1ZjIfUfwFQkfcX2
x3jMMnD75nSAy4Pto/Z5eI+krGkoVnMfOYDWYoCq/Ui3gFZ2gWvO4dNsYm7ZiG9v
lnjmBEmqSUsb0WzPAIdyN9uyXdpAx3UsylM8sAdZ0EjDERWap81iNFKv+H409F56
RWAIeamZNNOd8fWy2ldxluy894vTsiIDWon4kKRJDhjF9j1kFZJRVytuH2i8O7u+
1aqn4dqO+WeLWssXMy+GagF4hQ+JdBKBW4JPt58c/26qLrGPXQqjE3px23u0frO4
e4vdliunzbM4ga8Ley5Btia79BBhcti4qZlfTRsqFGCPGlcXeZjePvxn8DhC9s/d
G/OA1KaFSYMJyy2MBtKTHrPr9nD9sKoDCjNNcXTlU3zTWdwneCHsYT0YJ0GkCSea
8l5UYfTfJH8TAADB1ZaDGtxj32GlK8wuwGsTpw2vjO3i7SGAquzayGA51wHcqx8A
XqYTsii7WSoy029wwK382c1Arre5qSwRBF4nyIrw/+BCvaAfUyi2kr7fVSfRRRLz
/B1kg7YoipxTOIQ8TRy0eRkZLBSBSl/Z5TXeid+u4x9Pn6HQ+d52iBOPKr01/ooL
Ej+tObtlGCXC2RIGXJbrfd3xPq0zkkP8zf/ImQElB46CkqjR/hrVhqIs5iY0tN5K
arqm+xoOSUtT2ai0X3tUflFg+lT6w64okISZ3hoYmWgqp5QjCOKJV8HiutL84C3T
t3tPAwA2LUhbCAVGzMe4mQlMD1web57jLXFzJV8AaJL8Gf6qkapummcXkNxUPfyh
JLHbvbXwrxYDgtaNg5zmYQD+WsmV/3pbicGh9blSIlK3Pnq2SZA8YFS12Wt1m+As
eBWSSP4g2tLcL+azW7NI9Mq1IXYcrJ4i91DvhgFUgbYRZYFonrVVhsEecdWtbpoS
OjRvlpx135YPdwdzTDiZcccPQnPgpqxcu43aq06NIuwUNDEHIBVyDynQ5PnFrM48
HBPXmXNon1sY6ST0TjEkXjd26C2vGTAVYP6mI7YL5qvCJ36iX3nLClcHqn8O8Rpr
+nUOccJcYmtyN4+x/uCjxaSiaityKR7a2uh/RLa/+WP/8sQ66SzdoU7/u3qn++It
PUNS1lenemZemiEnOijUaUUipdagtLy+vAvIXP4ej3XUMYoTYN79bD6LtwtZrK9J
AhOgI0kFy0Dv/FP/HXW7QMRKb38HOt0h2FGidMphAv1IsbwHi8tw+HJ6unLl7AeB
YINLcX3vLjJn+c+lyZHzKDBG0R1hIC0t/MaccXO0OqU3+xWEKR5oHc/m71fCh1nf
v/MD1koj2D1qKCo7xByBChq15P1vvdYNOgeuHLKgMd3r4sulYDbnVJGs2//e0ZWC
BGzlIR1KMxgBK3Tb45xLsf6DQGS9IcvGhgkuLvvRBoNNOhGHj/dJjxKur52RJijY
Dm2ayOchOaCccJ3JsqhZlM8Od+TeP42S3XJ+zvfLv1wOAyTA2AaDqXS2EvjuqlTN
xHHzuRWJZ7hLd214foL8OLr86FlX3/spNin2bWHdWMdHKiY4ETJTbwyuJCJY9Bni
6CSB0K7NobNMF2ljZ9Q8m5f2oa4N64hBz8YCCqv8xkFgLQnvToTbiCMqnGRk9bz6
b8ZZHgG7IxFfAUggRJp6VU1fC9DWftWH0zdusm+k6iPnfpVi6xX4NGXdiuTBj8XR
wC4edwkukP0gfvyeUoNIXO8gtrvCGZJZ49mHmA02EebGInr+TbGnkZjGyYXKYL76
NnCnV55aAo/Qy2ntrSWq5nvlRu3CRVwmw0HlZSkuO+ceKqtP6/SsjRiRVeH2eurn
FzTPCyVh4Z8W+nSsi8e7McrQLNt0c1bvFe0L2jVzaHHlaURM1pi2GsmNcIbLlE3C
GimSdwgutyLUcU5cZS2O3Sp0GYB7/ec+CUvuWnY0YNBED8d1MI5Uf0MCsBn9SuCt
t8KU+9tLBKsgLFRnaShio4+H61y9dFSmT+4EHtUSKRQQfExIYc4rIZIVmIz/sDGl
tYTcu5E91QsWQhZnNB7IMD3Ot3waEmvrJ3U32EP6mwWGNHTd/aZCKW8vYgfWXTig
4haaFtNm8evMbK6AOVdTQDeKCt5DsxYEtjAd5xlhVXlLcSSamoX+8F3TijL9Boqs
+yMSy0gUU5tpSTMJBthM0e5yg1lra9QjBNfLUUgvI5xwvFPalGr0Azm6XOa9XE6e
vPY/Ir6SCNHn3YXF3qz0vDK8VFqfjVxg/AamImNXcGyf0BZPLxbBwkOOE7W6xO0K
d8YVxej0IHbJcJ8K7vvsY4yLmq90MHSFofkq1G5I5NcnYTslqzFsrG6RB7JDnRV6
csASWIVNO25+MlM7QKLoyDaQAUoBpp11Owq45iY3OX6EslyAAHGLECGMfUYEjvkG
1VUxj45IGIVGYkMsREJz2wyuR4d19adk0GojJxmFcE+EmO2NV0q5D2KdtVD3Xm9W
usncuLFCHwRcoVYcv+4jLHH3sXtcAsXzQepvMsGgvqt8o8vQFrhheCoyfmuRFW7E
OrkeH1stzIwTPfLJNZM4JSwijG7i7LdIuW3GsaNBn8Uubm0N+tEpzX1h4Ik+njHi
BEMB4AN/0fPhhw4Z7uTsewGXO7Lwj/77239lPOcyPwrPDg7xm+6aiGnUqZtkhTSW
cLNRRdcFftSTuef/kLeFvzkR9EpZryFA5mvVn28hyC+TIEl4Dc6t8KsGzzg11AfG
zizWsWuKZjsI1VF4Pzp57MBYa5sKf7JyGoqQzGJQfTstANpEFsL4zsvHZe7U1Ef6
Rs1uA2n1HrMWMb0U221967aczJuog5+GKQln7gWEA0u8YmwXneqEm9TIu3GregxG
Q3M6wh5mEQe7ohcdZl4o/3kNPPeVWQ7Nl7a6LObCkY60v7zsDVTRMzqjzNDU25rn
9DvkD1wUEcnXe63X3ey1sxLxPTECsyUlwV2AKQTLdzAH81C0FzFrFwnFn7GrxIX/
fbXLqG3zySB5GbAXTu4Q85bAqMV4e/YEvjqlGw+ryZaVss4hIFKXRgUOIARt3R03
x9hXhj84ueZa7fLMJdOCtRbezCiyF3qs9pn8j5BJB/l2by9SsxdXv1NWylF36YOh
Dbuz4L25NV321OoAL290hdYaivmFuWTUodM02TU0D0JGuuefFeDL3T46/5ztvh49
zzQXSKsqpt1CEveC4DY9NGocj//AUBJsSl7EzDKsKomTD48g9CsLUvcBcg3pWvhT
lng5/JF0ad9B+LOxpQGng4dvVpFRQdiXQTByVXu5maYQiTmdkHWMPDkWOnhKwQQ6
eOdMGuHSnzmgB8LQyUKNUD2wbkZwuX/y8Uq+0g88jMpABYIIisR9AZXzBN0lXGfG
/zWShfGVZfpYId5FaUPcnuVO2O01PaeZ/advyMHi/SuxWiRUrntsQx0TymgY2Uh0
DWykEsltl0Nml/2SSHvSIC9tIEOzmxH/lfpwC+bELcyDiuIGIfRlXCSdvURXYjSH
LpxL7aCArOlOhpZwZl8IwTjHlwDfJ/y6X05z/FB4kSOO7gJltAVCV5hE8N+eEMkz
F6PnO2fXgOx+/rX8y6bnNFmKbUCPKYm1qXPLpBOnok/AasqH6Ul2T+fhp9ODJsZr
aRnLW/WS0sPv/kL3ZfZWvQsuJavIjdrPwJEFFNVgttQf2wGcBzdpGYqmfn1KeTuU
2G/SSM9F3wgNeVtpsR8H4jEJNlrE2iR5nkpqYaAzdJjU5JxFVcJIlVAfM3b7zAJy
PIjklIDSkTfBuWVr66Gx0+W3sb/evZZIBZS2Y/KpM3U28tvw4sPfEnOlBJKk6BCY
tbjCRpbSuhA76VvW2s2jyGa76w6Tqlmm+M/Q9WoHNghZ+OtFrmsJbHtL5SPdx+wu
PLIcETobQNL7yzwkUFj9zA4gdGeE/mgBBYUf5MXdpO8novLNnD7booYe+uao+oUX
v+xE6fDKvYoRWIl/JbyOL92cD0hRdrtehwiC2/Sw4J6ECQojbU4oCdxQEAOLRFO+
IlMEjFz1xhWJxTtCnog5eM13dRdrg2Xr+oeAhcsT4qcD51d+mEs5n7I4q4MlDaqD
JY1Nx7J5v36WC13uFW0CbyGoNSDBWrDUnl80t32o7QK4gKt1GQ6Qhan63KK0c2NY
TDWLJRnsVuOu/iFH3hb03uwgLap2Ho8JGNde82LrLJwCo39R9tKnHvYfFu1JuaS6
5FbPhQzKmmywxdy2HZ3u1AMxfksMoatAKui2kZ3kzZs69xV5VYKkYzMSV1kmm7g6
Tvv/llm83oEgYD96G7JuCzOkvQWZdjDxR2hsKKchBsRfLZkS65dAiPsFA7kiU3wQ
3VO13/iRgw+2j/TjP0FU6Glczx0EUOUaLcAQ+oUuJXg+ChW7JbtX7pqcc41dzUoC
dDZTZRf4unwpwiXvlrvt5KgUSJokgsBr+ojUWtnW3ldNZwqe2oE5IHoVnRHw3OgE
dQhrmEg63O0+BEIsxpK152uPyr12DST1NKL9GDw4vcOYL1NlpipdMSfZAkOSrUzp
rfAB2Nk7tpX219BJ41DI3AnY3NdlMUfkgJW9LcdlAKzS0D2Sjt38BJ9vOlmBEvfN
DnYRh7vVwjFGWnLe0M8kl7Gl3kulXsVVwiCTAFQbiBI0twHYiSkxgX0tCc0cj87T
QxD1XinaTVzX6hoOyOxPj+cIDvocsaKzBzpudd8l1BE2coN6dFdIG178EcFQKctf
cwA15yyzCMIlCQuLSD0TxQ7Ex16vrveMIrsU/cKSSvJuGfV7dl4uOv+Lbf4YEqml
/dK2o6DaCLbH8QpuV5y6AKaSk+SelaZNDXRBvidGRUtuEG36RGyOwIdYTAgIhoVt
KlOdcFcuBnST8CS0N7/qQpwBI0kULV3lTVRXVPIVwPYfc2ScI625b/O+CGHCT+Hv
dRKpyMfEVepvyX82APHv0DM1Wsq7al4ikJF5rGXjXeyV2y6Dq15CdXO318x0t93B
BUDt6MwDpCPKnVNYUWVtUfi22aYmbOLKp6kY0V1TsR0VLdtJkQ2+He22upmvMWWI
5Mo5eyEi7kxlrt1Y71Y9AYlAmK19ZD80Pwy4Z5yudB6CbkU9HhWzlACOUyGDspRY
5ASwu6ecUH+2A6PSJy4NrUeChRZ+iWdujCvCZ9kVuw9UVq40awak3/5yZEpn7azK
OHk7QV9VON8MrOrpd2DElJtN5YLupErgLHHFMQgAKjcKI8NPuIMJ0VSnS7Y8aQPh
t3b93ZpH+4lkbUJQVRIzM3gTqQtrOZoyHn/J6z4Ud4agyNT3yAOOR+JEPgNBzSgA
oGjAHq60RXoN8+g63dgzXQEhFNsRPGhaU/5iE5DqVG+TPR8zXYI0xPG3MwkpNRik
13vh6xm3ItxmiRJVbJYnV5gfPjKPj9dSC6iJJlUw8Yf7o3NHLSM04xaJqPGn5gjz
5DyrIbvQRdBw8aGBcr2fGt0JtwYQvmJFue36HlMFnKHtiHo/lodRjWP5sfhwmJtb
JFuNflqUObe5lw/10tbkimnqhKKbr69n5UXRH01M+BJT/S3kMjtvZ31HNZedCFlV
llSJnYH5+9bWh+tAd4zB2phLEthWgoYcgNW/D43kgmXECiz1YUnT66NFkah2iVTl
KZ42uQSZl7RQvF5V+82rBimt6fWrS0kqrySOp3tSzUbLXnBkyOX66Ygew1dGhmgc
YXPkAEX8lWKNz8cQVKy5/ecGO0xYDMY5p7GkQs0AvM3rju9/XdNL+dj4yYStsXfV
1uHULRDTiWp+bDFDhuSUrLADdNNGiGumvKUpnA9AOLBsbIMtFKdH/xp/czjukmaU
Dn0BrddoKPjEmotBIYSze5CaB2X2/pNzRtvFkr4fAZmMMl7PVFdYgx3Xbbmr8QF0
PZ5E3DPTUbKKwacdCHU8gb8NK6ab5WclSMErJrwCcr+f7eJCKmOwu50yX1d/Lhzr
6aePR9V2zEJ0VJl1gz66QKgbwMIfmT4ItjfRbsUCYgDnu2cRjiX/Q3oOM/6E7Ti1
e8ucmvQB1p5xNuekOH9Qv/yvslW1fwTg4JI5WzDHpceL0JUDa9SpimJW1t1Q0XZJ
IqRUEMv6fRhR1C+HbFU8hdFE2Y3whs/LGEzMoqQ0SbG7Ajf4shzKbzK3ifgMpEdu
HlofW49dvmF33RL327lPlOUcQU83LHZpqSVO32t3Bg/ryU6KqTA/BTWpeK4M/D9A
xJlQ1v2SAsYkV0yn7V7Lo65voJuD/8fy3ZUAEodkDK0TJMdDg5lF2+qML7nmi1n9
+Z4czw0qTOaJhkWlvmkkSyjFAw0tfWiy4aSbR0iHWScKMLBbGiT1qd6BZ5uiFuh5
I7LZd9xnEuGPmullXtDZMjE4DoH445rGAIjBrURlS2LZS0HvbjnJYhliPnQ0oLP3
YuVGdV8iI/G0XPpZMBKXzt5Ez2+MQj+x53D5CKpdK7IMg3RVuLAwzo2yeGZ4tV6T
vPPgITS4s6vyS0nPaoSHCxO5BiPeUCkxD6vHNcKAhypPUPljlYrrFQgdjV4FegOw
TC5uY8SxgxsuCJy2hAgGWq0bShVAZq4QvnnzbUtVqFHCKuh0IzlbQXFyyUOxsfVG
wOKpbl9fNstwZQ6kkCCpF8UPBfrGMrhlbUK/yCrwIGrLBFA9F/dwuYOZrG505krB
GFCbWNyL1j8uneZMhb5SytmSIgFId8GmXJ7rcAl9LqeZV2wHtKThrWO1E8POhNnC
JpdC/nnI+IK9FgE5t6qk0qVA7KjbIBg6WS9QB1rkzjezRk/6rTcBAFnuXS9eeNzg
DMewDRPDt9RWbpDW0gDGvPWQw+UvXiSBfcNSvdqF6Ay4OzGLeIW89dGUVzKPe5nA
wSpH0wZKw+8kCgLpSvYuc0kkQD1plMzAFjrmKiRq9ZwJ/jstq4Y1a9vustUiCfyL
TijbObS/R+LBt1IJM8hcGSSV4X438KQ7tdAuavUj8tMM+TBbgVsGWXz0KRWRrY3p
efgqo0lfCLi5KbgrhflPloIZenTob5/j4PdzeR1h4LZEJkhsJmd8eMn3xgcsgWdJ
wGUW8/2SFnqKxu1MddJrVUtTtQjBc1B6hDq3sGxalB3v7nz8ZIH9dg2QiGPLvGiS
FVUhmJPqQumVwcOfPgwyS7Bl9XCtWG/yGuP/Aa5hv1zT3+VExgwEOH4mrAhF8HpY
2WF2aOf1tSL1uy7rghlJ7gX1x53NaWMgeojV62FzeLj5XBolTgv1Xnh1twu9v1E0
Q6RfP5rOCTRgbcErfSICo1er4udzPkYUe2nkDieUwapgMZw3zSn1tPPFUyhTwR8E
sUjrzFqv8pV9ifduJaOG4nFVe2BF4yumid8ygvV7X424caMtJc1WAQ+aK9ll3NBA
LfIzTcQaDYfyrCGJMuB/dAEGK2R44oIW5nMcLnALoBpJoAtiwHqcsZGld0MTeXy4
aaQOTnD8B/1w1Wg80wUIPd/76jDS3HAnXnZ+vYUtJBNCC40RnUfqobFBOmWUAkGn
BXAluhuz6BipkNAMClsYXH/w8kzCVPX6yApvqWZPcTuytpkZN6+nWr1hci5aHfgd
XRrnUR1mKQwKvk0WSKs67sSA5AiGw9qjzIo0ZT3wgNBBnQEbElAlcMKkrb4lb00g
Mpff1jr1Ji1+3xdpNQ+3vkrnIaEKc8VrPV0EKk/URuu1q9dlHAhImZVNvK0S4pKV
c3W/wo6nOKdcT6IWgJmMWAl6UFcPrCetLlTfW/XiL4Gkos5eHTQvv3uGv41D0Rga
9ICOP1cX49krEF9/OeVrPDh8Xxx+NOoxcpYYJ1AyiV8V9d9GDMwZiWta7U69R96W
PHDoOuISFF62Qv3L6qQORlx+78F6LY5r/pVXl2xPP2jxwFA+duzUcUWPzCwXvV8K
6+spwihYnTEBb0g1AanYd6s19BKOFt/+HyATIBclGXWXC0DQ9DYYF7Z3RrBXn6YX
0af1vLSwj67+NaXDZFZUf7ONdtoevbJVJyJUqtfaLwS+WxWFyXSvdPH8pUDj5yng
ekvLhldVU7gBelCAzZnx5kZ5sxY2rpmwWgKZpmj5UNXj/2qSA+zSyN1rHMquzgqC
BIKia8st2PI43ANAjJaIfssEFT6PVNOYCnUr3WwXXqpRwOiTCEa/GBLEzFOV5yvs
tyYzKGt0/9Fm8EBI9NqGzLtIyheK3UrSQ6LHUb+SZv3DS5UsDYto9ASkxzsLdIBk
hKMzm57SnncNxG7qw5WXC/DUiCQ4bfYluIbP+wsi+9vpyd4KEJ0KA8D97DHKaqem
YW+WBgY+v00kW0z8C/9OVkN9mh2X435V1DcS3AG3atAsYz7Ve3URmcfNfWP8ANcE
w8Ap/i00A/zsqDqKeZldvmCEw9LY6OJVQehN1pM7e4lcLNpkDYLG5VJ+arzOnzaq
YI3S5Yw649beAgutbG21e3IVPQLI8XyrhOEmlxB7mkXK9SBMD1B8qhWp76cv4M33
hUKHgXMQsrhjxbRD+4yvURVGJcIAaOEJYoon7sCm8n5Dc4615bgDbE/61fw9A2+q
P8L99UG59Dc9hED66lcbOSD3uHu+XH1EleaumnyOLvHLhiQY9GC8DWNSvNEWVItp
V9ZFXEZ7lSlyG5T1QtJxoeBzNh2OAzZrrhgTy1RHMSlytF+8FUZ8fL6KuQWIDUu0
nLqyVNl8poaY2QXEpzvqvSvKm0OQ/KuSm3nOsvuiAY4IlwB07Qm00eb/j513jt4m
xwAmrMkx3IVlXfGjmRyzAFEThkihFgfm5sT66veuO6RIKYCbnK3201gvmQrip5ef
1UPXYoON4jr2VOvBvTemY5LQ4eYlrEjbKUjS/ED1fHF6SIYoteFF+/qmQr2g4uPH
PiNC14Uelqb0315BRWur4rMU29c1cq14Il1J3qLlFeKJX3CMRZ0S3XbXpw7ZARof
QajyCjzuYmL/mKmUmdy9A7Zzs9Ahp2wgnwKORZy0/1cSw2Ye+fYO8eodTq2emyfw
JG8ApoLSWciaPkP9Y/JUUhcPa9MBwn+0dNiUriEPbeEoZpaU45AwvDCKBOv5rzej
cKGaku2fky1p40/pifKqqVJf9PeQM6CoE5PgMtP9pfhDjwyYE4CeFL6F0a1gFXPP
UnaJOzVJfwhN91hc2a20f8O5edtfOm13ZhK3Po+YyDoICfcO1WVjHSOoDh+4l+H4
lK8EbEaTjhiCSe4GG5oPmTLBI0AHJqvfbmMVjgktUR+BisJ/BQGRdaYszPRUOW7r
3w0He/FLfzjHb8v90V3Hn8GdHFmOxpHaRA5wmCISBYsIFi+IUsu2a9SIy9cC2cA/
6HJRGvKNiUDohIbktxalsH1YUe5PEKVLjnShyfo8DISAbkdhFoJ7jJl6KiCl3dIu
QAPhacJ/C6hsgYemLQrKOYlL6E1GTcgGKEQbXLN9CHpx+IoBQ+Z2/zAOYDZng3Yd
qlGDy/xoI1Kv4M0829nq8Nr3Kvcu+ujlzVRdIZU8ojh190cPss6+OnBkVyXlz0Cg
WGsFSi2KqB3N215f48LToiI/ymw4UnEj4uavwKJ/Af+MM1RHf8nF9TNT9vLJC/TY
Yv90nO0vYkp6e43jdAkHX6WRkKtyIzsIIGSzXSCnFMDjczDL0wUQpPeVhS2sVH0q
TUUeoBFdQoDzFiUODpEAC7cq5AeSdZvE7NmfPsWlEWSGVDPkhv205OLdItLocCxM
g/cAJMYsV+3q6yWdr1C5Y0AtNHCtb8P7+Hnk88FcTqXhPM8WdCUxJJrTxoB6OHPU
h6K4zdGJOOqYwDMxPtvkh9LKzAfRNFVV8jk1bnFdxSc5VVJ5DmkQusuQy8Yp/N4w
BEsNxl0VIl+9PfQO3+B/K32SRjUJLoEZr17DWehk2Fprzn6LMcVHH9nHpzZuX9F4
qZUVjbyZNF80AXUyOdP0dhORItfDgj9hA0CkusYB0dO5qo02SU2bnXn0I+dedTTd
orWRi+KjCWSl1zNVnP8+dKlG26vCqpen4d1PaqMnc3gNSYq4AnjrzonfW83DJ2W3
hKKXTKhaj6oKBAvvhF6WTYmlAngqGMnhOZmBFLThWxmW18+Z0qW1T18G6B1lEKH0
pCki13bIkrRywaI/uoqqss0XmQEJmB4XFmxkQEJsG/DLPGmpPIprQwL3LrATQH9R
jpph3DBQkxcgyhLaDmLlcxwW1mvjqPWiZdptqep0wMxZE6KIHCget0DMpEtg0HDE
HPoay2TrIf8HxkJ5cZzYifha5sgz3FSGiIbXdYQfPCo8nB2RIxGVqM5HcYBf7sUh
VpAeklfk7xHhpbyng74K1LMfjPYlgDM82HMK60xnfNCvFPYHfuFe2YulqRZQS2nD
gGiLNDK5D04gvkFF8os7950neD48d+7oZHR7s4AnheWM40qY6YIBE3BLIgLDP2x3
h1uBdsbZbC/K+abKYHd5oKP85r9qNLuWHHak7PVYX0W++39reOQhRoT6QtbKnTyC
Chafp1y5Vp1ft7Atd0+ZlGBudPTg3UTiOPkUf6pjAkl+TAEjM5/oUSa4gyUkzfbs
gsbhsGge6EdBlVuu7ga+Ap/hRYeVEGhDyJz6KlymLbolZtXSIzpFD4m1O/e5sKNP
r7o6oTBaW2S4wtwb3jm2erbHOxACzdk5PWotNW8uUf92mk5IqzDeShOhUJqX8nm5
NBKeG5tARTS6QrR3yNmhuXVGIq9MVuN/31pkA09DAF7YfN7/rBK4yapQiA2texkR
bE+joj2E1k+pgog1ofd61q2Qw/qdEwdQi4pzSfRKDdpahqbadn2ZgqRJv94BK7BA
WGZj9MDCncJzR55hQyBFIBa5NUfqiGQSg/HskJqgjk0MTW5Ja7eASMyW9ueL+sCT
AsZq9nKomWnoWGu8lt9x6QypMmTw6Ctec8HkmYzhPlqO/2FQ3Kj2DovU9rd3jSvF
tck/dta0HY/bHVfMMoHPrrXGIcpgqibHpveRXLYZzPX7fa/S27bzYb26L9TZ2I0+
XP6Z9U7ZQQBEU8jwr7S6rnvIlccJ4xznJGsbbqegFV+Wkeu/8aZ7XRlFBzLwO5rQ
xwmlCGRzUuzckB33yrvMdODBRl9ZphFEsiWre9dc6qBw4VngjmFQqnfCwfIpCq5J
Zxl1KZzeFhJ4Yyk79X50yzOBDaC/UYHXXhSj5M+g+Ovdp91FAaKTwfzq+qb2U2zb
rKtRtbZYkoXiF4DMFK4qgjmw7Spv0t7xdOpROohnYJcIRKH7VB8fqzmLEGhmHJrv
9W3K/Ig/a0miOP6Q5RSK79sLkKisYS56GESuF+bxCMIuF5l435uNWtBOFoCBoluT
n6e4nLO9POaRASAVkMb8PuLTKNTeyoqpo6t3VkkdzrfA9ONMAh2ctFqmvjdUh+Uc
XNu2sRrKLhOgYpMG/QavbCwrYMHLy7HuyomGHD1MHhj3AaaBCjdEn1hcegHLL43m
OYgg2WfJ9r4YG13xTvhAgKHm8OksanA3fZZKhtlIG1Iv4PCmrnVUgdz3WtSQ/vAE
jZUEcoxZrpciBFy5PuvNcgTRq9WuMd5/Ouz4T4D5fjqBjqhY7dPlfIbq6L+Cmr9P
cVHotOUcEB/tDOV+HvQnU2QVHnncSRrMCTPDxJyRLx6hTjlGPlW3erV5G6+7YEwR
JeDHNF/gIe5AorruScgY7lwGNW9xjSJUWfQjSd4WxVU8/UmQl4h5R/08I3i01NvW
R493oNZUgXVTnSxVTfzDbg5A66Eg1T+nhhjqDGIVyi5Y7bVbOhcMYi0P/RVhD/k/
MQYF5mhGI4+xameSKpMECpkbDVLksRPImKLa+ZITni1nMOqlFAJR3YkMGtRNBrtr
XRe8G59cJubh/9JSobF80IE0gfussmF0npbSVD+SBHu4heAPBbOp9oD02BXrpYJK
6lezONSCPeLw5nU7meO4re/3xHQ3wB2fX/3NkTjmEILRRWAgrKP9L4cOdNyuwM4U
UUnjUS3uPip8zQc+1K8c5hf1efGGGAIJ0WuSrT3YsO99d8iP/LM/MpXvyLdstvSD
KRdww0JDu/y7U82rPDgAlXsie4OpSCMr567TpqSozp4XjJql71TS9aokJvxt5cYK
ZyOxCmfSMsYQ66VEDE1iZlRBB9BO39WaZRq9fL8dKssO9j+zYbLkdCA3Qn+kIW3A
6/v490TdGYPYh50kuL2KcSBHmGeRxtBJtxQFVVk8xCfRDbgieSnBVbuSvOrzahOE
xNRG272J3dZKgn1dOFdXB+cGhBOPC14hkx/QtbVeN5HJVL12x9+GFJJicINEXX9z
T4tz5H76eSZbDr8nWJkA7KHNFfVLXjhfr2JTs16Sb+Ha0BLw7olH1iR06oJo4pt7
Be7T7kSRQTyn8VmafKJh4bjapZRPjQPlKeV8sdI4sEVx5em5bFpLh1h9dJsxtscJ
ZxqTMgX9SsXNk+Tu2ESHnESmxfWar3AzVnh2QX2PKr2x9ZK5gLk42Zq8OwnDebpf
pC5IZflIPTCht8bYHvBgFEsf17OAkQR4IUgCBvcqJ9cidgZQbzFPwApyHHDD3sHp
Fu0BQP/TFc/zPavCdlE3rxX9i+W7VNnp5R5LeWl7SKVLGwV/GcIquo9guu30IJWB
XPZ1rXKpBkw3cV5hOmpSMJZfjCpX058yTk9+gaqBPaLrx0GfXvFHWZkX/R/+8rZH
Yg5faIyQTUoWrrdD1bLcHWDIUg8tM2qnxw58EJ2uFtrsdYG6OxqVBGcqkb+tmaF2
jzNff7t3WQ15Ds5uIDwpwVBMBtzl7JCpB2ygwdt56on7PZDoHhUDbbzZXTjDyKMz
nnUkXoYRqcs4QchLz9Udcmceym2tk6vm28/qy4I5OpXaaL61yKjByR4E7EerD9uu
SXWO/d9s+zLXkxUfE/nf5JasnnyeBic2hHXBHiMJMTdPeTcDMBtGt12TJHJtjQNa
iaU7fkJilFb27CZBqDpHJyJYMTVhooMTDh4yQ4DNX38w8bSeuIgLqbN18KTdUeoq
Cx678d09FEJpC8bhFtIJ86KPuiq/dI7c5rP395+zUwTPwrTgclKIcZpkwZANorwW
z9CgajV/AUHfTfZB7kt23vKVAgsP6g21VqluUzXgOlxuegAGyD6Oe+ePW+Ue2lg2
GHb+KnYs/h2wGmzLfHLHow==
`pragma protect end_protected
