// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
g1Avmu2GJN3Wo/PkCBulpRDC0TR9OCkeY4URdzmr7iV+YvNOB/WS0cgeJOAACRfxXelmK67VNAN7
yJfmdfzWJhGFHR3Cyb58cI+OnRy1LQPufJnptW+MjN6Ep9dnSg8Cqr3FXKhi3lqtWoj2n92SF2qB
VOj0bFzyLjCTQ+elzd6rklRMPWkgTY2qk05GxJvpzYxdhrxN9QQLKFrMzgjJhjwAuR5AInvxigFn
3SLzQfMNJeH+lgjjFevI0ceykmwQdPnd2197CGGPI5rsOeOrxI9Ux0LFDyIr1F/g1tWMpj0cnH37
Lu4/u3F+zH3RszzBR1WVcYZpkhRf9vTc5YXJiw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29408)
VKmsT/asDigBRkgcJ7YpCzC06bhygRb6Nc4+xYkUgk+J462r597iGBMudasKq/iBU4QEQbP7jjw8
upzth6OicINtrJkLSveSRPKw/Wjwx1KjxwP4tcG4KbnMX7rQB+H74VWbaf92mb7mlXfiAcbwwK8z
YkUcVYfJS3m357lA9U1xv1XKWKVyzafdbwY8cxNk7yzLVFblSZTLvqBImtCDuhsLbtlR/DG9+ErP
0LBShF5JZvqCZM5EAQHBI3CloYvg1YJhvWMSNJQdBuZD4+92JKKRb73MQnxZ0C06Lv4tzeuyxBMb
asrehxFpZhsTZSgipmNIMFRCzBjkZ0J6d6q9wMBqqg8ZVi2a15qWOBV7HKyV4mfJjaGGFzSO8DMS
Emja2S4laZPb1/fJ/u8ux8aVIxZZdbVyp3m6Dwc10wc24333Cga8/YMSKDgKi0OPXJISDp8pqVhF
DL45srqBSU3T8MKymxcikXrgWE0XT6RmByzWkWVj/veLk1Tg3TpRp/WrzCTAtV7Py5sCuQH/+7f7
A+Pm20EFeXwLTjJSjyfU2rEwwUfDk2sxP4ThtzMI2amp6+9ED4KMbh5ujBwCHV4dutEGH4Wm2JPz
BgfOI3Y4ZpciEGVrJgJ/1RKK5y3Nx7hONPMmeIqUal6TG86AkgAkNeQhrL1+l8vh9ky1DdR0qcNI
fpqbyHVUlasc09b+fQHjm5VI4rySKFzypLKpsLVg2HpgS90isgMAXYzzQED5O2sB5ZObPcJX25q/
BWWsQSlgc4O663kqYUlkKjSrs6zH48E4UDrKJW7kiPIVvoz68JX1nW9jWgQIfeRZsquo+cFEy3uU
KqjUHdxGqIRLsJe0io+RrJj1GKk5ektvC0ThE7jA0pOTaME1m7JPggQCu64kr1mmRVnOtO0V1etA
Eqz3mnsStONOza87Hc16r8iOVkL4UXd0JOBkDPrRk4jtquKfT+8oeqrzjd3oiGPjqYLLbxljns5I
qIDVV2coiVrvCN9Sm6ukLsnpDUJMGenoE5I6ehWsD0GUlXeoun2sGgWNT1oR+p9PmZ2o3HpqeuxW
Jy/64jzhJK7IRR5mHIsaYsU34/0Oxj+3Fx+xu9e7dO5gXnPzxBHB0Sg+zCev7Ts+khQdW9x2UorT
H4348lfxkKIFYs0vOo8WmZbf1pjf2Y7/n1ZH3iaFp+hDQ1CljfgZLkfr5blw+3nnhrz67+/9eTha
O8PGKyzl6XGMEEwvmGAACIozzsTYN3dD/N76Qe3k8XxqhGjbyM8C17urTFb/XC8Km8KrxvlEKlOS
NAMsdIlIusfbQJG6D/a1ji6X/SxYEWzBc4gVJg3L6rEz3wTc9TpPSCKyhjbf1jyxcgRVol6yXuC0
+3lq9GUUOMu0ei6yMOPTrjNP3rZrxjzJpVOFDf9tkH+/zqHIkTfz5z5eN7UR+fyLr8+lpECMPI/6
O/PXVtG/fuM015VRrROuKQ5fsPNwxjLbreo3PssCx7wZBj2CTIO4s6fLZyLs3WI2OnuPy0qAUHsx
Vj+don4lM/W/bvj6i5oh9JjODhec9/xgb2Lqd5w+O16e2YYzoMxqmY/oiDzHOe4oOhW9D9zAhsQb
ydC+0bu3Sa3CoOPR29IBINOTU3fauguhMP0sUCiLNyjBqTzEhxtbo8GzBcCCJwYD2Bsqq+5MaJ8D
Y7eGxb7IK1AurwGAGBWYc4HdE7qIN8HyO/FIp9eYqQghQz1cadm6HTirsibflcnqN1LP00q0fQ6i
ojWs99rhiRhKO0zv6asSUqYyGaDGN35nwsw3o2Gx25Wu5NTxmHvAiPUVpaWigqRNJEIRXd/jlym8
55gCrj1pz/VKOZQBDmBurynboMnCqQyGp19EXGLDXBeEcxBbkkAnHGDS3U2pXh2uBuKaWxnwkt/a
adYEsQgQCPWlL6sMCQWVb+MqIYyiQOoezPVT5wjOEzdsbX8/b4IvmDoN22LH9NMwBgyy9imWHYNe
MLnTreOLycdpT+p3jisql3rfP3xFLTOaPZ9O9z/QLEcScqSMZoknIp0+S6756hCw+gVce17rWKzo
OIEyEUcEppMN6Vti86wShapE81sYoWO5milkSJhebV57xZZH96rgXlTMXzjS6r1RUgy8Wpv2pB/I
oyYLryP/FFWqccNlugJf+fPQTFHB0+h1WZPpvXPvf+KFyQjv8PAOV1EdAPE0spoSckRwqQu0rMLS
g+uSZPekzylnXa8c4GvWmeoJWZoTsBOB27X2gmfgYn2R0tJCJpH4elMcu/adT38MsJtZplpbizM5
dprcEwxlIvxh9xaujt0c8Oxdm5+Rs+I8ac5q8CPhvTHPtStWjyAKWbqtGPZlgY5eVMcHoTiyPLii
2NVAHbusVvB1ytbtWq7I6B7ZXx7rCdYI/yyYA4UZDBsHxY1wOJP4OXhYFmArbsXO6ogzuxE4oEko
FUZv9vvPV4L4y8nWUVHFlM5JglMoG95h4lzCXhubgbmucxFHuc+7a+UrU1NC1TfHfwrCA7sPuV1n
MrFey0DXGiQRkAp3JflAUhlP+SrjHfWpr8C1mqE+UIc35LXMqTGkm6EZQFVKsJjGmxiH98mmLjdb
aUXorssOfM4bGjKNpf64um/DpjVoWD9Ll7EAns4zo/GAuvaXSbu3hIirygYZaQLic64HYXorj4LF
751sGRXmfAWoTEhQrIOmL1upDUo95ESN/3NjBx7Qps5P3mmNlsfEVLjK9EVNpgG+qKLFH3eYKMko
SfgCRE8v7mF/KljI8YNW785TvLx/uatf7AYHfh4wPmwzkIyC6/br3xtDyXE5Ewza3N4Ei+G5Zh9z
6EkfeMrS0fAczRNjxHChh6KiP8KYhtLoMsrerT0Lgg8aDTdNlY3bW1ZETYG+wxk/uztuYN4BwWTt
zc4EVsp1sfxTR2v5XP9Lt84j04ps8vU9fmlOIPel4Hc3kGfpnoMqIL6nQs+gwvGfCstBFKz/zOrh
8yW4qS5qN+DKLxXvSWqNc4SVXWhm/4Bzn7k4aiX0RvK2+xnsbToTpiO+E7aJZ4a7QwOn0J5FrxUI
Z9Bpz7xuAraSgXEnj3NIf8m8kv1qO1SYfbDH95kRGItNxirahNGJokRHTyCWRZFp5NYO3TtvVWcy
mWF18Gr7w8DcyDEp/lW3mBWfTkPsZEY+e2I1NmUkWf3l5yN77YmqSOx8PBKs40dKerR23eZ4V+g2
lkwC60LIn0vA71YdOg7iN60Gzraji9hSJU6oQXU7bzLRvfKYyMUPDdpOYOi97iQa3OxsZnFOCWga
fwj/SvHqGj3/U2T9oepohgsetxF3N0r3iDiarOsqDYF3qcsuyNwdeW1LNwfqljk0srZEqNts1po2
Lh1XgzEldH1+jwW3eCXUpwH8jceNYzH9tIecpMtVy1ucgRW5m0tXF4ZKJLGrk/EMLtPphVD1Mg5T
nKRP85DZr837s098PmG6dJZ85yxCLWQyFI3/OzKL4BEDQ9YUi6m8fjGDTPp73qwr8m1IeDM63W3t
tyibQZF6YmaZpKfsUEFAWPGKs1AnLUUbBudxjiCjQjym5Ud2sK+UxbhjDux5JUeD//SbgdAkEYrm
k3JoRA3cB6nsfvBbOpaut9CFGFIbRDTCPvlpFo4VcVvGEQYCgRUgSYKi3mlqTi7aM1AYs/E/SsUJ
fxJB9XhooEyO2gNTQWhmHW4Ty80ej8f0pJwQLaFl7Jne1P/PMCJwKaxOx/v9kEHS4GxexgDbjAUN
GUXXT8Nf7nPnKptre6xTlqBLhDx5q/vyymkfeLE5QwzXnsdW/gJPtbKK8JhYF/NpZfDqzRMyJrj7
Fyao5IKT5lCVPSkqWIVFXsg0+Cr9r2a72DWHDbYNwKRnGuaaLiIFQIhitfOfvJDAv4JB8/lIso1Z
S00IHrSTrthABU4eJB5RnSuqVGfMDnYJbbRKCB/BtI7y2PI39eKGJ+KFp4tD8daZsWNgSTpZm7Mr
502WhzDL1/Ed8ypDZYyWQGcN+teEQVMX6Fa6D8NX82kcztC4N4hlw2aEH1d0Yuqlsen0VOjbxH0J
Mbe6etQeS74Lzhc1G31LyBGPOGyhFAO3hAD2IATT0H3RfcuTbJz903VGVv2e7MGRmq/7lO313AzD
RdcXH8ouQxWBUwBGLlzeXebYj3246RN3K72W2loDLaJOAhHiJm/q0p370WMY5C53bG3O8+5cGxCz
IAng7Sy+lhPlrIOHp9FCoEefNMC90akw/0bhQmxJAkHVZKnJBD7uo76Fa/VjB8CZ8ZDMSeOhFuAs
yIzSTbyreR+YbeFI/yrubd+ul8KJ6YYMuyGVsBAx6eVoO5AvDp1CMLcwOM73cqvr6eZkkFoQjIu2
FQ9DYZkIsak13LygeUOwyZs2kZ3Z63q/EYsHr5gKRfjCXRt/X2IYyZp3rVFHqZS623XsYxHnOUxk
hQHDMCRuJfkc69EMoYIj7qYPw44ZpJJv3awCMlRY3cBEb2a+g/8XxKagReR2sIJDqUwS5opuTnUi
HkDesPlFrU/8N4jr6PrnwPj0z8J6msfqmN4vFCZzJo+zP40Q5vRg1pZvE9xtG1WuOykxx0Br5Enf
yBy/6KJ8AV46EJcOId3HdBMIPjML3TeW4KTtK6OsK2AZUu3YUArQxFI2AKBpHt8sCtMSogVgEr0y
HaH7WginwpNZp7fse7t9nZ7JSuiwwkkfsZwB0/9/dwvaEO1XofNRdcw19priS6BCgJOS2w3x/g0p
35qCPJnrxTV1jjeBS+BDFCX+0rE2UJ7dV9NXui01POInXgYv0WnOCI53SlmKLUY48QtpfPgJ/Kw4
+mWnCA5j5nmAqzYRuvfI4+c/cxUhgUXIem6fPb72skvT0A+g2PuR7uXI96Cj1Z0j3IoOhiXM2Xl/
2+ua+aRVC9AsEKZAuXwL8+73TksasoBu82OQGpIoPWMLK20YO4kA78mYKm1g8/B1jagRQ5CzwkCz
NyrOqGO8SRE0tsl6AIgEQ1jeXA6dEVOjrFJ5AMnbxY0GtseDOGW2WhBeuOVKMD14GOPR4CDu9y3W
ATrz3eOjf2u/qioQtyhrJ11NQjyxqZQ9RlAEbnjS3+0Ch9yDDF2DSgTyZxa1TzORrqHItjFf9X3T
4kkap7m7tQJwSo+IYaEJtVtC1pOsydztWfyScaKbMn8KhFBjoM/xOFLi7l7s5eJGuiY8MW6PtS3F
ywbiR7ChSIbdBamFugbx2SmtZIf18Mioc4JehtySygvLlg5hvT6a6mO6kq41Yorig+RCuZFiSYX9
WM+7U20dGJxKClpr384f7AJAIh5QfzHH7cZCrLFa6vIgMTVpWQhZI3pf/cgo0yV+rfOaAfu1X072
nsKVw119/D64M2Zh1icKkImRF4zeq6msG+3u5hZccNFIK3SOi9PrcBoPEjFEHhEvi4n3Gnz3huMN
Lz/6OOTc1ZZy0jH3AZrBXNCOO/pxmdGpZVHNjbrZ0HoO2vC6XdVwHz+SiPiq3xleDppf5OhHAig8
OxjWl/nQwyo70EpJ/IhIP41j8jmy0cbSq/eIH32nln9ARVGBrgxaQ13ge9S5MWKU1PwgrcL/0d7x
PlvyXwA+Z5MUE70yZ3ch6Ln/ea34jQGhakg5Ft042fMWPkCwvqeNFPg5jeNIYiGbMOvVyIXo6/QO
bNKgVMi2XATk7i55g8nbEX1iW5lrPa2hCl+148Ao5ZXmzLbXa9Jmz8w5ts2um7dEd4pAUFKaI8H3
qgA4dnVZbR6AILPJfnNs8lwPfZ3DtSdLzmfWh3EIwtIaqd0bUHcHSu22sqsGWR1l4kCiRWOIRldu
p+S/INvx3tp82fMaYWe+LWPTw3tOCmWE1rbkxBSKbbAJRtud/sl7isUmkXcGwRwps9da2yZXTh5S
o8I39Z5QzNUXMbpAqYDeLq0lhT/7Sq6crYUxrU7BC/DrYRxq5yV4YNn9LNPH+a/xrDYgoKexPHXz
aUucMqLmpAeIOf6nKmSeWdgJsf/HMume49u0XSZSl1srFueFtxyBw8GjOSwByeKhZDiKRJOdl7ad
aMJiUxFxWgMvivkSl2ao9Y0XzFuYbg3vdOaCSPMVb+3nAXCC3g5yUa4+CZn9i2SI1NGFv0DeHEfY
hslGUoj1kyM6hsAXHSES+ygiqCMiJE6OWIfUJHALIpDuDRcPMoZHUALuO6j0Qu2SaR9q10BB6nBb
KzrY+bmniJUnXvXnJ1iMXwu+n1fbEA9BYfPQ6/m6U15yA+c4uKcSEs3rkeD5QJKwvRx4XZlQ+u7z
nfCJxy8C1HopugyR7yOtCVYmDDbz7UJOBsdZBZLnjD1dpPg8vQ4TYArhfy/i9xK4jqZBrP46xkgW
PBSm/b1XGq902CB9W8YOCQaGYBuB/SE/dbINaczXGaGGFr3B5Dj+FVbZ/7mlNXXlZP6AF7j55sQc
TZ43YagulnCA0Mv47L1xp4RI5Tsba0afBiR41/V/dN0Vmh9lfSL4oor3B7hHEDwSH21Xp5kZFcn/
9GaiDMqsubGZyyRNp6+p+nhYKTvTgXvv80GEAkGZjdPqgsDcaqvIYYY0iyyjU1Glij/sCod++DOM
tvcx4qHQAAt6kwkKpIs/+xxK3kwmEENN7FGkLrrNaWQ3kTZflG0SlJKK3ALICJygrrpYMxmOgC+0
tjMJuT2Lb6hOdKBDjt2q0Cukr+gv2yiCW5FP84YhTpApTfcCUySVD01LTLf3QOC3O6BuCfcf/S24
A+Wy/rxQ508qgHrxUXZy+hF+xEAweehqIh+gpzBMFH555E73feGNdhLnZG9pDcVlc0nCv1Xt52d2
aUmxL9H0/1cPfZ5gJb9fZ6gJ+u+6ga9/Q0tiAYKhK0fYLbfJSuJrUWw+EU67jIC6GFJvLRdevmPr
vGmQ9pkChqkGgHma8hBFU3YRdD3QDFO6M4gZ/HENXImF10yfjCClSxdA6WsidO8DjxD15aLu7ocR
aQjNj4vBorrHlHzSxx3n4OXVTJ01B5ymeHbg2RgHTlkKDmXAmarSIq8/awUm5V8u+9HgxTlPD/1U
cChrAQjG61E/7MdnAdT8+UdS52rD3LuOmxwOi9k0syKP/8C0DBG9Vu73SrqtKKxUKy55wbN8aoP9
LlHTrEG6huS4awtOGx/ao7yfWt7oKgLmBMdgoIFzHq2T6F2TY3mz9CeTr2NSZWsUfD/IxCUqlXJ4
7YvLNDNiIEaYyQMQGzZCMyXk7AT/0W1yc2LqoBHoErQR1yltbKcY6ojT10dSRdv5T5pof00dAeN0
/pf1VLnWyfRmm9sYOHyQn6Yq8eH9TFO7VlPSn+z1azBPL4rC/RYXnLjPSebqHESzSAh4HoNQN6WD
cgM++fkLvyhxkCtZFIy985f+XEHddv0ZccilXhK1VE/GIG6dt9f1qAEYf4BBCDmGOi3GAD12T3b0
TeGGySmuwWOmWe43djsJfB1MEtC/HnKDJSh8KLMZOwTRJafYGug5Hm76Aj8s9djjwlZgla0wgtWV
UtdSQR605wsnG8F+MImWxt2lsSsVrJL6csj02W0ILSwhcLttblkZBGjwyZGWGbQBmYYaRV6iU9EC
jiwCQM5zk4xrqk+uI0LOjKcPe+a5tqw/P8vDUg+9zGBLspsHCkHGO6Wg2gj0jExnpgf3563t39af
zJD3b8LKM13H2mIq/dULm/KE9+HWNoK+JTpyJ2gOtj1BYBuheuOKw+ue1+WiKcZzoX0nLo6M/gF5
/E8etkGT9hnEK6mj9VuKmtgK8ss0ZfAduSYyJV9Zd0wX6+Wai9ABLOsp9DyP5/gxQRdL3QovmsGN
nRt/lAFNqnYpaYEy/mtFFQ1kAf8vH69iA8/o43DLV3XLdltx0ox5ttxFFzI7Qi9fR1hbImOg+00G
gEIzOsMcdPhzNHQq4ufjCaJJ95P5Vb/nYBOAIgzw4TZ/7smN3VJHNrNILshQf14pv9BznayZZuTy
BlwnCnkSEW4DpffcVlOxfsBbGg36HaD4hM3Ni2MAXPlWfmH8C5bf5igI3P1RUt6+saigI5kn1C2S
55W154M6lHXudkVibKkNrIeKlDZ2WyF9VQA4XzJAO+fSCpOcS7ak1P1ms5VIE3GvntxQEZnfrXQE
9FkVlL8aum/ebwSSRqOhEy24/HRHpWvtq6x9sIetd9ZM+gV+JnZ0p8s2dUleN6jCyYYpgokRPy1l
jlmD+S2IKuJgjfz5xbl27i4+pP8poUXeZ4eLUG+BqHcmoITpUY3C2kpHf30+Ltx/XmGastqlEMuY
c/9sn0eoMTLbPtopwgqB7IeMCxBkXUKs0w2BAVsigDTypUuIq8ejHHtmj0mKlgf+HQm7lEdvNhUr
opThbUe2QE0WGHsDu1tl1wnVxi5l2DsmtEc8IhbS1Op3pfoK6frgpem2Tz+iBDleO3KitAXYaiQZ
c8EmJZ1QJ95Xqd406iNR98xqMkoChKl20LL4hVILRqlgnE3rXWOyXIJsfjBeWsTHHjqUJ1n3O0OK
4KQc5PCMbEBx+7agYnA5RwO7mAe5vuQssDvH93OXwJy4Z+3Vyo7jtV3cO3pSJMtbJ75B3X1JsF22
z9CQNjzFIt2PpkCNkmOKM9sFUOrKrrZD6K7iHGX/iHtewjU8wVIMdzwXEAYYuLgJPFBx7yQ/ec85
/lfcaSMNt+iNTvmS7EUyulQpq6NKpzjV12uiBlgY+IACfZ12XaRSwwnQSwnQYqTdMDQmZ1ifXKq/
H7Jeeef+w1sttHEcXjtxJyWDBeMQA1aQrPJTJLxAQt5GgF5ia6Oo8yyXxmWsqHtspCt+HdMerKD+
pta4/tpwlyT5MxbBaWNSVR1qT+6qUI7qBrVwNgfosLNftfKxEw4MZ+X/XYqaHI5p05nsqdlKFECj
3F7mkhsGu8d/GcgdoWiVCfCiXzxheT/+26pUFfKfesmLLp4PLOXYKW+gQ84q2GI9IEd+h3VyhVIk
SHVaqm8iq9i+EmEWoJoONy/1W/5KLc4gzKgvNh2ixtSVEb0RWmTVOYE+6ifGkzVcADAHfBYGz+cg
2s5PGUlTa6LELIzCAOWEFHCDCG2eAMe5SgbFHjJRHlM6jwASfg+orBtdsMvnyer+wq83IpClpu6U
2w5ylSFor48JpB8Aoz4Pnmw0qWfwH22Q4TPkbAWw4/wQY2z/CDb8bEKxxzEQVVYeRcDZTqdUDhDt
V47t8wszJ4+DkU5dG28Alzz1czOVTtgBdf4M9HLGjFXcNs7VfWrAh72ic29UfVi1OcxqLHwCR3hD
NY3J7bGkkL5mdqtAOXYGvgnIX8ex4jS+n1Xapi+yhNdBorIEmvKmSFM1LRTy0wdX4bHJgWRNLF2w
aMR2VF48oYL+BvPZQDJWAAmGT6w0c7mUW/DqmNgBdDpO0ucLXFefdnYnwoqxossj9C6GCj/InvbY
f6MWPGnKbW9PM8DknkU9//0mlVOQ17B6UpJgWI7G73bXiidQJVl+zV7uoad3g/6OwkgCnvBGVvA3
+mkFLJbFIX8JNUPzbur0t8Dku16JiiCkowAGn1CF2pbETFBiH4e+8uamjHI+7Pty6IwCaJAwF8ux
1dz0XF07W0sslPFybTwpJ6apn7ZVyY7bkJdLWUeBYCty+2/73+y7WM7BOFBc8oRCc0NS6O2epxT7
DzX7PfWPzV5WKAp4Ko6mK9t9J8oc2KECUJMJEqSGYQFcFxxuoUdeNY+XD2wmb1fcthTP+8ZJccuv
im966IcoakvXNEf2UXXCQ1qlqzb5xMwfse3qVvGxe3On87kdcU2nc6HAJHvKT/C5lWr3t3pNbEzZ
F2tsQQuvftdtwRpFEDU5KxW8phkjOd+XcTXF7W8Q+/Xa3QuFyDM9B1hmh3NmXNkiJCB1471eFy10
w7VG/kqsokmYI1qVz8QYWXCYWs5EX2cm8bMxft32a7dPlqKbjaxASt/2ZFUCXUJliEoWETG7gZ97
kmmKRgCPkdUNUCouMANPTGIUCUAdW5duftL6w53efqBQOyCyoMVp6Pv4N+Xr2lsKkR0VZstGOLpw
GA/mAj3ocA0U44989Q/JV0xNzOB21yV8zfpN+Jw7qtVtc0ZgUEMcds0oUF66dPWzMjYa3xHaUTEe
g8BMmA+PsMFRZdQY6UvBzXzV4OB/qoQg7iAZH0Ex2/lp0u/WfZ9mN1wnK2OYD9azW+OAL/ssL8JT
/Tw3j5pGRjlA+fFBAepfkuuI4W+FU5aii5eBy0/oS9qNz7FLEhDKmkKZ2Zth408EOxowPtcufkLu
TZ1uQe/RTTCc/r5ko88+BgpNndaKA1vhEBQ5szDQbJLs0HcRdLvFbsrsNyxD0HMEW8V7gxtc464c
Sxk30Jmw8WqdBkGgAa5XfFMG8V88H5LdOAsOpg2q/w6eLGEUzX7c+QByvKNPizudaPjJ16vVpoG/
dHCtX7D7kBH3TO9a68lDDLWZbkuC1eVdN4u4ZuUHRLFr9oNoyusByF76qBWTNiC2r7a3rnLqEhXq
lgaAdQ6bjJADAAldG/y7Yetszk3EDn0W2vngRy1IJN84t1yVV0IuVUuAqjmFzEEiYfxOb0VeBuFg
v1JIbjGIabsd2Y1L5kcdC19h+OfWD1eCR0CMW7d7EOK4eiZrWuC7l6xk1AgoRmQdaCrhRwRw9ekT
ecX37ZiYBwGzv1J9x8jN0dZiMIGeH7Hfg3t2BKB9Rv3akWFxVzxVFxCTcXTcwAfBbtX1DS1v4eMl
xbJ3nbxXMEdq2ns/hOIRPvTHv9LMvS/sRFcaU6V7fsQ0/x6r4ly+7cvPTNkcxVSw8ge4k8PTNVbY
V+du1x66By1hMO8k9z5wDjkbyrh2qvpPHdIz6FiOl9crb+b5gabXyZwGQCecT6W2d8k7tEQbZXFl
VZu/BXUqlpjxgpt+Gmww8ckmGwolq1kd/fdEkpVfmBmUKlr5jyNJ8DySKkE2pLatoI7k9C1P2Y8F
2UsXjS2wJU1t4hm545fk9Pd/U5oJajk+KbRbkuSIjR670g/Cp3HSt75wAk68bO9G2xl3RZPdiSxZ
IF75UPhQR3NAEtXcjDqcJJ9sOJ8m6TFw2aK7r+El2ESmjiB1F8+1IbdIOWMz5ZJZ0dfevhJjGnTQ
Ts9mjPYHHya77UcB9ixgSO4+4C6vCaQH69DIuuAIk8auonhjWtiglNShGa3OaLh9qJK+KJpXaG6H
ZLjypNH0wdVb73XSL92qiFt3XPDzRYgpY1xtBj5LuMu2618Z8mGRaD9tzaVYD6G5/SecMwDWfZ4G
9O/tP/xqQpMJp9FsTsacPPZIIedwgacG2/F51YHBol4cC7QcVzvZ7sEW4XA1jUc5Sw5j/+KTpU7b
S+zb+2JMO2KSSM5uS6O4Z0iwk4pIMWGLSzjjN6P3hOkFYtpX0e9mIFrCNcVkOJfVzBIr3F9XLpwD
FEIdgfCiLnOcFjOU8WV+W2P0wOryhJJcjMu9z4JNE9+2Rsqc9gnIOxsmW7Zo2gpoRYpgv+/3ojbN
hLaDlKkUEgnm2QWWu4qj01Rk5c4NdtUHjSMZ8Dy2D7lx8iYqsrNARQV4ATktnp04tW0LwJCva5w7
EqC4ucjxiegyfRkKRXf215i077R2PlTDoBNz9UIIS7pzBPJUbLRmNEddnzBayLQI2HM5jGulDxph
zosU8VtNWmpgg2PgPnOI0SC7tHLaJqPMbReKvmLIYxnpcPw4cfU39XIhOZ4LMT74NH8KUhNJ0OdO
ec4Y3349wKEyQT8P85oSdkcrwaCvIVG/xKNO72TyB9oCN07OU1LjjSN+cW0UxqzNx6coyNKVUdCb
eBQof1PQjoOPvxU7S/Mb+wIwVGcgD/ZH5NbnOMfkgbQE3mCxNUmcs5kYo4THcYIABYJeDC+tlLNc
VMp2DD09b5JE96rd5oPl9hizlU2G5RFp457XDSQGYVFpvD4uosZUS/Q/wq3oi4Af1aiplKxICPAR
eAX3iX/C4HiNCrVEyZL9En9Ok3TQ6FXQar6TvbTWvbWDkVqO0MIBStOdSqugxVL7T10TDw4umwnN
Vy8m4v0WjPnUbb8MyBicdJfceVKqzvmbBwV5upGAxcSrLhxetEgVg9xwevmntXQXLzViBxAdHBNI
IMdnIPhX/REo3kPeT/Kp9TT+uiQbSSnexl/v8IGpbEfrjZI4GJoHVqK8g+NGGs1OyYLdiYN3r31n
UzxLwni+3S+XRogqgxyrkUQzWMlzv/pQoEkeicgFnxjq7XPO50ucUjsaDDn4hKCCcx798FWFWhzW
/4VBGUcWGlzI/nEFRgiiCwUfVN1fg3qR3EY/ylZMAY0SXjsCrQrgsIlChUUOsozaD1o3TCAloxAN
k9PzTqTCbp4bpEAZfAN3GtQV5EK/wGjcm8K3OU8ap46Me4582mssXUf3SS7HU107EoC0d92jZRGz
tnTALRYZir46qJmkhcn3tf4UdQSSHcyvlGtlK/vkkLMGGaTeDLn88V9CPC5vGbCXZuqHOu9yBgr+
MlSfAf2bp29lfHRPwVrCMKC6Xvyg3oB97PPCudVD5Nqxs+51gNQR1cq5zwqAgEFwOSbK6kn9Flzn
YPzc3gho49i8FWhryrqEd+nmuRqp8eMT3HhLYdYFae3S8+VLB+o0mlgWLw+jKpFvBENDPRdCAQ8m
ekhOudOi3Nhyyl9+yeUuUH/v93YPsb4KKmfBwHFzI/uJUfgmyUfYs/+NMIGCZTaRikti5yuZNl0b
LW4bWsaOkAFOmetwpvlyj9xkf8TJ0ws5LVJHuhxlGDHAx3modR8H1SIWN68L4Upn/21WFITfsOmP
S/su1qaIL8vL/30Ay6h6WKUyHhWRS50dXQRS8lODLcPwRC1vU9PsKBaoAg+m1AN60XIGJa/d4Zi/
CL9DwJ58gAfN6437pJaltZD9Lo9kOHo37DUqLk/W3GnVdXGLLFfmUMUkc+tYWaxCAu3nJIiqE2NW
JwuKUrjtP+OqaGBC9eSeobwlEshpEZXUkcPrMxgyACxteSy2ScoTLHulzB6b3hJkPO0mryo91gFK
CPV2DDFPIrSRdthU4puG9svMnWUbdKStyuUCD1atkz2qnnU9seJ8iaQLzpe5nZD2RcEPpOiuhO15
oAEPsAqki4sxQG1g0Ipn8Uiknj+T61YJuYIGMITdDhy8umfO84zuSvnglInVXHTzKSJIyD2aWOlJ
BuLsSW64hStxtsA5EhkSgFTnusByv/QKWF6HPNBLBQWsCMrQUMAJ+hGlzVTNNp23J4HL7OB0fXAL
7Y4tLfAoYMwrms1XxtZ2MHu2SIsjuc9XGDmRAmp7YafqkL7ODMFWnBZC9AzLKSyvSJKLQANpkze5
Gl5vJhAvEeSB9RC1wfif+Pe9/trAWAwII2GvVyjJ8Vkq03vQ7zFydEW9DPKeuKNrLVAFxHnUtYB1
Q1FyoZb9/wzkkp1wmZW4E4dve/kwtxbjxUtoIwgYFgGVSOYMiXvK19uToZsSKpVh5UrnE6/Ntt/2
ryAQmGlOQQraL4ZdqI20DcOmL11Xqi9fkyko/7NVFliFLTZAO4gTFrHD933e1Nt+J4KrvKR3OEPZ
EA61005tYrYSLQBu5AT3ZrKwE8FQJsybvig6kJ4+TTAdcD6limLaooCxrovMVSBNo1JMCcNjn21Q
II9/z4d9dfITvuDL4MtIQraR/X+1GoPf4OxN3SDE41529/1WUdweRhuOTKnjS/0sPxgNC7MbEKYB
K1tWqVtAeQZNORVjWHQbOo32r1BTz4lUAvO7WQjkBS99gRmtv5P+G++IpmXdjowXySfh09EPf5R4
Jtygy4RVDJKoGmVeG/XGVgfsBZ1cRp1oAtg02cydonw9D1oYWHmaYCkPz7tN7w7uXWIdyUJQ/XXA
6EJFHPwEseFkeI4LKdq8+Pq6UUkFrv0KwLZNqzNbtXiptokE1LMUxcCM0jK9MQahplWQF1lc1tII
8x+MDnbdGA0BdTonw3tCBaINmmFnuE3Nrz2W3oJysXrt3RGZn5ufKFl2qysS2yG4Eco1C1ML1mHx
qTlOgjmO/6WlQgVaSSTFF7VlQahynWaM3CayitfWyW9lYXaOMDYPERhXKyEicD2d/z65joIZ3K0O
/ZQL4TXfjdyf+Vlwa88bD1hpHwAeVmj56RW/FHfYpuBRVNDxxNCVAE7c3PtlCGJNDGuHYGZSDrmi
Rh7JnXvL5kvbDVrSBrTxC7ZzQMbNzARC4JuGFZob17XJfPXCsWi8cgdRObYm9hi/F7vIuHj4A0Xz
UrvVG2UKySY84pd3qQ77KkMU4Cr/sSo+s33PyRjGBxxxaLiCc/t9MrSi9N+HRmDny2GI+STUCXBe
8XE+RXqoyrPyQlfim0kV6dxuv0J/vufmEj7dYSXIELIFyVYfV3PouU1IUokXTk+CL4fIRlF/J27P
V+y5IV9FlY8Yqqt3mAia0GUFRvchbX3TsSiFKO4YiuIaYc+6p5pRSDBCoinRuYe0KPvT6b0fi89V
XQnlP3hMzEoRPgQMD6uzFCSiy1VS2ifa2ugPxg2h/rxTf8oxnWnjfht4xW3TBzxsMHM04+wSHeX6
ww6UNEtoEJM3xfbFFN8vEgxCMo5wsKeDL/cLu88KYw1mDHfG1U/YOmqN3g0yW1+4H7bkGMQcY28n
Os6EtVl+OlkbPL9btMBmZpOMGdYzRzvKDtbTSZ08zoi87vpnezO+HOFtGK7wHVMpT0CsC+tU/eHo
9QSRlVXbq6UUtm4GDza1Nso9Xf+zg6PryrZmSYaFdxq9MnH5l+ySHImNbHTpbUkxANBrb0a5pHYY
iY2cH8376lqro0WzrfaKZV2aA2L/2mthDfHw6hIb739rN0Jjj0rBGimEy2JlqC5W53ZE4ijiAPkv
Q0U3qf3SUNe3PazGQ1dL3l5e1mvKNi/WLupKsrwmtI0uu11+R2MQmQa8hX8vo6a1iepWRzfkW+wk
anuL7wx+nl2JjH7f23tXqyyuixtchn4Th3/PKIrsBE8llEYWemtkyIYwT2/1Y6rDZySO+JqeIdEI
vmib6iZhs7VvF23Ukh2cdPUkp64kDTi27DkH1+ONOfccIh4ND3UT6L52GjFvh5KDDZMPEZpAOGRR
k5QOJShjKDND6/oVrDO5mEsPOEkAHCicJ+bbioh+xDxiRCRvco+2c35VBjk4XNFndyixfUgXCwDx
Cg9chk5u90GhTCO6vCYD71bOYKMGi0rkf6v4DDIex9CuESHhtAgg982gNANcx56LGKRJbvvZvN9b
oLP4uBPm/Zeov7aUTnaw+RpMTNo7TiR+zNHVBFhbW+ImedMt6YmAzdURR3tQ6HdgG+r+imaRJNEs
o9nuvcet+ttORMBrbAPStF049gmOSOe0/E42WEDt1+1hyf6ewX3bFGQZYb0AkDMs1q33K+7vQH5P
0QOxgQVLr07slqTsdnHr8K7nPJo9v9pFer7YLTYKsPA5AuRnC9m+ypdFHBECIkQY5CefCW9FOO4E
Z8lpnHW0yIEClr7atH8UjEOeaylkhDb9AbgkttOeybi21X3m0KPtG8KOc182N1RJ6EYHremYal38
cMmpA19KjtdI9UNKz4f8WUzMNsVDZDrKdng/jDBiUH1wskVGhw9JGXdoGChcHtalk1OHn87Yvqu9
ZJvdEZRTadsfJ3buoK5cQtLE+nyY1FYXLmIdB584d7Qlv9RBgg72rUavC2yOnhsdarn5gUPFsrE2
zrFwLVSjAg+FURXVjl5yt+Egvk+yZxwzBdeJ6dZK7Kqu9X+AGylLycBQojbDnIe2Qe1ujek5bfV6
d6c9wajb+LjA5z1cVmGsEMF7xq2sQXR0WGDbpOTlvX/DU1FzRLvEmavYxqJk236vEiw2AIbqznF7
uyRRI+B3AjxH+EcxWCCJUmZ+cgnGWCtMfDz92PkLiz85DJBzpCFp2WXJJfXB4bJsf0TLvT5z/Lmz
wqgO+N7LXanVd55AP2VLzdKxgl8zPk3HTjq6WJUYNpgne4H0b88tHPrE/AdHbGph/eKXnZIPY/Jj
vMt5HF2EaADWY3A7ImSCViLbdjWmHVaQLuAP7D55bDIznXFHIhtctYOvGhOyXWkC4k0KwVoIVQ62
wyNT9ZshdXdVYdIErcYdyZ+uh26LiqKC7PwOgzt+Kxz1SVKvpDtUILbvIGqcG8bKa5GRSC8gVZNx
MSmqdHLAoJARQGV9+J6UP9V6yUes4rkJncRRj9/G3n84bVAqLcbfn3yWadyjWogF5mDUg/E/lohM
1nBD9YGoqs/T4GqfUPRJ6iugfcfWZZNBeW/qFvTnzSOX9k3mYgLlDnFhbV5ul0bTaJ16gcS3hGXG
l3pjBZoJ9XU9TaY+z+t24gjj6yMxWxy7ew1628ocZCc3dbCb9dpcnBzL/KmcYOt+Ho8UTIEx5Tu1
/uMY7MNAyDvVL/2TAcCsEpKGEmVLKG/heWzkUjUT0YIAI5CRr5pKJkUoXmDEr5wVVTwTREx+uC9f
hR/I7lQi695onzyC5pdThpC1K7vhQ7yC0Aw5F54QkbMHhtu80XJMwQDX6D9BGwQR0F6xJzXpynp1
Uh8fTM5qXeoTV7Yk5iper+wJe5XDi9YgU0RfqvFrB4q9HNosv+jCYIhzAOFp31Pnkxiy6nqMTqgi
WWv9fSLUG3izbK5zVp3KIOF0VtaOSqkHhSxVpYSzfOJC/VGX5wN7uPZkE0h+wdQCqTxT4VYo/ltI
tw7bYAOX2yH8CFxhih38TxhJvDwoJppFAXpnn+hRx6BPkYf7yrRktp9WpTt5rGbfDiiHPU7cOT1M
jqISoEzaXCvP+YAl2hl7QSCyjebfmMtVUTgkjpcKIj2oDYuBawHimw2mH5JegSXfpPfEdOWYLKQh
QgUYEd4Lw7Z/+yEM1xD0SvWzUvvNohKNYyvtPgyTwM0HuGNhHwGLXuwbmIA61I373OBp36Ba12Cb
XriH+e8AsUaR8OKy8JSw+zug5RBPMC6lkwF45c8FSa9+08hs+yqKSip/te3N2J6J7n5mLiAOfC8V
FZ0RlpBttqWlFUtJacOYUe+mcnyf82UPjKGbOayWbvS5d3xPi0hAK5z7gUAAxyNA4dfAKBcTl3vo
LyOs0pVJml3xQwHCvE3zXJIy+gp+t/dMNJhNjmrzPwvmOVgER63jW/e9tkL2oTXhEAM+j2xBBVUr
5Cpr7UNrs+2qICH8Syohkrg/1XJql2gpfjgJNGJuFuJeX3UD+yC0g7//kT+xRPSJtW94aeIayRej
bcLIxabkhMFmrACgw3LOzzymltOdqoH1xArL2HFWxe5EET//fIEp5JtHWfoiMd8uKa50zecmQqS4
yPcFV085wBu7d/Kw0s6GcBj3P95fqPXpTPlo2mqhKr8/ToqnzdG4Qy5U3jXDnotMlhtNQLEPR4s6
6AnEjIjK2neJD6zDKpiw73PhozK3BYGo9BDB0XVWxo9KM/io/OfBtM7LeeUSdmYMxlWspPIDqVSV
a/O6J9CgU50/hin3m5xE3ozNEGQfccYFEv95y10b3Pds7gIZO8UsW9ZCY/odAedgtsPXXXNvCHGh
FgNZeoOb9mmdEcLPR6k/Bfm+O2nE/SylOYrfwVtn3n93X40zojb0B48L0B1Zj4rRqFI/ZBq0BpHj
VvlOE6OUpG0vbFZgZrpRMxk7giKP2Q6Bh8N/5QKwaH3Wu9ukcBz1ZxBTUSt0u6VJ51V+iFqk6Dkp
QH+G/LI/ZvvLTwYsF1LBK74EsbpKNxKOoDfWE/yUSJjBG2CRSd6coJvS0eP5Qqk6H4Z18XKG4pKR
mhDSmTdED9dchW/HkiRpOt7bFv1UAjJDVLYZ3kx0fWC6WJVC8d6KZTrppz+6/nd3ZVHxWeIbAULU
3t6DFpQRoB0CPjtMWz/sqw2AprfDcMbmgy890E1lZAiSVK2L4JJRMkg2zR6iDP26bQXeEV7O7Mzm
EKSusMFAh9VhsSTp8+PO8zejn9HUVR3k5RBwTNA9/t+90uxxPDsi+xxfs3GPcQZpIc3d7rcaGAfp
7dw+r5CWiJE9usMrUnmYnUNW7L4Re9OtCiBCqUNEMfS0Dh6rAZ+znGhPfANYvleRzM6emr+v2JIc
uubvuSX7rhNZyWAyzPaq1NeYzt7cxNQL1rzOpKYfC0K2HaxoI95KPtJbOHSvJk+hrzKzxsinYZDd
nqzC1l9jjp1aLKJHteFkVzok9mXHoyzFdZVtw1I0rfNRC29UIzuP6AHGWEASKwlS6mz90blvpdIt
pmV2TiAonFNAAKg88rnZhiw21nALv7ZEmSRix2mLFR+NtODsPifRuqPMGibbu0+PdKO4oQWxD/cW
a+d67QZwsMDaETw7X4aXsFG3UfPDbP36CgOaDAFTGUNdbjJZuBH1CL2ElbRP1EKNkTs61QaLaNk4
EJvgARdHcTCAflWgPov6B2hjmpj/+yDmlND9k4IBQnY7ILTKHwkOfPNgjbO2o5EMJ54GFRgw7ukW
uiFpXU/C6coIxX4Kbl60dLNPAPc/ZLj4HESlUo2d9a7wzcyH47mkVXqpgSityjia+CjUfScOjp1u
JjZMScMGMVE/r6I/Z25NV8A0oKo0NLFJhRdGxroCBg7ru8x7B8WtHDZiw/uoL3aQcagd4L8C7lf6
P+lxeXJAaNNNfrfksfBFp//8M5c7ESzVMa1NwK1lmJLGRtvOFGGdqnWcoc+n7/S5KR+lEkDQs4Pu
i3jhBb770P4V4YWJS8xBIVVR31pp7RFJ8HkqiCTJiORe75HKjaTjsJwmG7Zw6qbDMiVgLzl7Flt2
Sy6lYEqcrsBWrsmcSW+vLxdeutTV/HxMOoIc0WVFgDzJ8lJn0O0g9C84GdDDjR1kiaKPI6Be9q/P
7Bn/Vdy64g/bkTqYs7VHIbt+gUa/dQp9ABk1IYU3iZ5SahyA0bUc/g65ic5zxSnNa3ufhQ9WQ0If
Z+zf36fqmS5UicEr7X4nepmTG9m0DL5MoP2nsWvjVVCoc7kY9OXy6NS8HbIRjvUfKHcY/w9ZNv3e
Ah0p1T4K2LX9ug1F5Mpns9E9YgUQPtxwEgxEX0qQtlCTbaB3ObgZF5F+KYybf/b2IOmNMbC9/EU+
3RuXwGjKw+rxcGMnb5tU6rKce3iuKHIrbkCxcsieNF/qOfDl9QhAgWzqAN2iJWtVvS3AwGdWWTyt
KwGUK7Ex+T+IwblpadgQ2wXvvuk+5iDcX11QtS8V0f6KnY4ZPcDRn2DylPygBPkWCwUWzLxnkZz6
Fm3X0z1efRDkR9Y+4+EK+0MW7kniHFRWNthbChP0sjShikD1qFwKIxCQqv6ZEJ0TkRu13jiGCOtw
COHudNWyAguU3dH7QbBwD1KUZAjB8st3g6MeTIXKWdRBOfGewGNYRv1KGt37upDOkxOy0IO/ILWd
wEHYQ948C2ntrdiRqkYP8A7omYgxMeL8EFFF29zkZNdI2BChbCENLhDxPrDoL41fCZf381k7wroE
n5hK38341/Yz+GzbKd7vBa8cZeqEHbli74zC0w8Ca/rqcCk0aNwxxSf4b6FVDP8dSSuQD3jrPQfo
H6Kiylv7/U+HDJsVK2NqDYqHcR3PRe6STDFYRd1X9b3pcEW+i2qkPnQeIeSBOoWCtxm/A1tXuZTq
KlNvCGHchizLQYU/80nfRSCU77A+ZXS+xzx+4BSyUeInZ8T2+WYPKmrgRR88DHBXTNqirU7E60HC
viifrNvGrBoXBgOmVcdnBGupL0KhqDzf6NCXThgZ83wn/p4CLqF0SNIINNPy60Sq9AZT/UN3jZVq
vukSiV+fY/kaSKCloNGtkHAk98RJpSNR5kwWK+nZZCkWMBXsgS+m08ZZMs+zRAk59sn5cqIEMR9Y
4FKznXkcy4yPDCJT5Sx5V7zUM/732eKB1Ylgv7DBDaGCYOT2Q7AAFAWH36VLH89EFUnncrd7U5AZ
g+YjYiafuynnuyxQS9nfzjYLyY0TBD7MHs0aS5+kfehioCyrcbJofLPBWyuvKgviZNqvXqv0STWB
lEtYsp+K/7ftLf6q1y68VI5LHSAZcFMbdNKmGNGaz/JDTWyR3xEN52wWNQIyNFl/Bls4P1kLvG1m
G096t4q2BO7faERIYBfj9da9xVz65UzsKoP8YEcoEXk11Nghkn0tjw+zixMzdWEs7r8V6dwC2N5V
I6imwiWpKjbw4XsHJAOfkGwe/zI8r0952ha6IhzW5mu5CoAXleZko7I2h8Zf0GWTF9b1Kf1J6Kk6
GaWPAafoCVk5N3aZYWYY5RDuIuXq3hE29litznsUCeI9B10daDynvo7Au9o1S9eIca4dvH6kv3fp
2C6yPFuUuhwhHeyrRhHccn1NC841S8NzKjiryfmXX1DWtGQF2XehjimWVj8VrV5g6VgcvpcGJesD
jno6mJMz9iP+JqU7ZiBsNGDjBKB7MLPZEC4ek0Mnv1X+VRcAvQx6VbA2lou6i9/fTM+JH8frK8ip
Z7bB/4X0dlHQZHLAeKVRHpbgVOcHNWjpad5BonJRAQKOfcXDqj5f5T8LzywMWhxTPQt8NoGgy3h4
UlrN7hTaQRi8lRpuZgvf/u8D6PYo1zLQ9HvAEfV5cNYwDFADHtqsbv07KE6QUn9tEcWtUlY6y/K2
moJd/ZAQ1meOLnsCmZDQXGGKPtXTzveYdWyoeL1UHBphhleQmNEWDo2y0z092OIyXtnWJglx8z5U
pvt4PVOjihss3OtnB/oEgiBFwLwaQcF2zVPhJNqO4K/zJIuSeJj6sltmSZV34BrFyztufurl1cZT
ioyNax00TyXDI500m4OvPsnYA3JRUQtCFx8i3NSD4T3jU3CSN+PgcyhWi0F0VJux45KHmKt7iKEF
PGznG9ZZcWdZGMWACq+60mz99IeKm942Eo5ZbaWURAiYeaY4WbRnMb3D1pNueU8t31wyv4YTuMCW
iV9ygcNTy0gzb7X/y9oTIRFs0BFJMrWMylRMyTvVwke3kXpo8fPc9/ksp3UNwRm6D4Qf9dsbSl+y
m34bB9CZHlaZUxJwsU9TNH2jrjEvyiBm/un52svZjKQpeND1Tq+9EA3YpQ8+RBUS/HpZ9aRNtDDI
ohg6jrn07McaczfalQCX4RgKN+CHOZZf8Jjys/zAy+Z5vhjXUsp07KOegam46Xu5ynHz/EqGPU0J
HOSc+nJ3cekXjdtc9oI7rvzO0NHsdyZx+N6lsifriqRzmIrkE8N3wUdNruRnUnqsZ9RnjvWeqFTl
2+tMs7xf5m291scwVmBGClWKUK1yccKN6xUlZ2kh5KVA/6yjaSxuibVJY/lYSfLCU2Nr1p1YqCa0
Fr0nxsgKEj0DKMijuhnzaKouLJ6z6dtdGFgCPQO9YG+0m3g8pvGGAeot81hcu0VOgLfgB2Wu4Nas
6LE3hBq0ZvHWzUnYOvGjvIj4NpeSfMOeyKZuVVr+RZYnU894eD6Y9BkYXL8ht6VVatA/x2sQVZQ4
PbrQbnHvrvbXTm+bK1Dc39f6JxnUK5jnpPP33VDR7m9g6RB0HTgwxRKj4S9YUnUm/fvh7m/l1jKA
8oIAiogr+V5prNTsoJ7CUOjTDBpH/saY3L7uLZ2sDmJJMYzDhW+O3Gvmuec3x1yNfWYRBzhNMVze
rfk4xOv1bqE/nhPYfyOyiwnmpCwHcR4Dvnmy6ChgGnC1tB5536IVlXhvRkUttl2AWWVFK46S6zf5
GCQZ1kPdcYlM1iwDZyWFVpAE1aPQyT3bWDIZiGWOTqgggaITWqmSUuNA5dPH7w8TDnyNBX4xGs70
ZVu7wVa3D5m33PEGjlq0wLGQOlrSOY2l4k9iopFVcLnDGReo/C8pDtaFSGVRL6jIsLfFy73ItHZb
+k/a09TRjP6DFu9/O7QJomgryXIQb/4rm/YqN3YGs2bZQugaGiEZS8yzVE07+Cy/eH3eMgQ+H0qg
C6p8/x8Q3TmG3zJlzjA++Kk68AW54MEmHI0lGTzovgPdXWlyqbeNBR7sywo8Po5ATFdqJlvkRDWd
L0bR2au0mXf9jQGWFMj8Qe+FHKKSoT1EOyOROCeflvw5hNEW2Rlx0AQDnTzItSP+/0Wq1hPaMTvl
dS7GTGN0b4A5FEMg7grM2mdo/n4LuDnM+Kg4ngX/55XI1jyC9qs5FFrAJiFx3we8OAAv/2cO1ob6
fSsw7sPL5YjCa733UaBx+xOxDCSmZ/68q+V7Btx90FgeMFF5Xy9VCAmx5BbZbz2z9OtR34lgTcU8
KbQk6Mqk/3biuKUBY2Ezwu6jHS6gzfJJF9x2+qIxA2zJci4yTpwQkBDqzzicXyNjF9d63QQ94cbG
sRgJSE8cRMkV+heg3xAhkhDWNJ2rAIGNM4MBk0SnSAOdvnXOPyjDJdVrIyXfOnvX+fmnZR387UXC
MxEhpWfQiHqe3hk0LfpYP14i8QCXd3DBPFJQXG4H6PrYxu8bVD1Q4qyQJ68l6A+rNOecxQLRkDsC
uRlQsiEHLN6NAnVGYthJZNUDnXKrH8BzbAuhZh1HUfBQCxsOmntcIfEQsLf+LNT8+z0riWAeuTXJ
+P9GONeNxylFdZtv5uHoPCqnFUlw4FXiFpXkd4MKtK0zoYGTV3APV0maW6Ddr/pfy40sSr8zgG0L
cFfO2F9n+vId8WDYv3VksOO+wh624lO/jXtSDvhgWuKtrt26thBEKwb5GT9Kine+kxyg42rUXUyr
mm6tRUN7Og4p39vPzBUeEtes+TUU5rf2dYlfGyyCr9OmQwpoUiM4ZX1WSodPBc0OadoRWFtMtmkK
Dwvhip7C0e0RJJ63gugfW+91YoWwWIQM+XnfaM2HOJqx3z+r4+vE+SefRI5+7eqisp11JnehzAgE
rR5yH6736dm5fS/6Dgsp/nkgTG2BBxZ6VVcVKBsEJC17OO0CsIe7faavqi1VztNdHKKSlHhDwthk
Uc/O9/emyB/eXWOPhScznBjcmROJkzGGdcB7dJDX+WCZQPcrD5Ik7jBCGZ9KcO9F3CFg4W6fA3yB
uBFB20ioF6Oz/KO8S88eXibtBZE4wFpsKtjEeF7o+5lE+g2YaJhhff6ifya8Jwx8PcQr1iTgfcG7
hzFf7pcBWalYZHc8LpTXLztip3zWMhBWuV/vRMGpk9g2Qhuw5DbEgQg7nuzdGFlhD3mT82CHWMcw
RH2kxLORpfLZHN0g4Ftw75cfu7pnbuxL/zI9EbkxfF4Mxd5RN8P3oIXm46IUnJX7ZeDZPIdgMDqV
DLeIHVRO83InF0zqAHM5sb99lVIMceOBZQElUchOp5gJr9KV+ZngN4eYiWL4PuBnaj54F9ox30LV
QMfhTZPjs+APOJXroPqmVv/cEJt3OhlklRUJzdKMdtx8BZVhJOQErztP2SiQqVrqeEvWBQxLvXR7
nPYzrTEdAAigBFhdeVg4OG7HyYA+eSRzkIORZzA5x4HBmDeLOsq6GOzJZvj66IAKZDa8gJsuNPDw
L66BmqXok5vVa4Q3+5rfRa4qb9cb9Ls/IP+pvq4fa+hzoKogo8O1alpkDT28bqlXDxoUpn8aW0qY
pHIS5TlwPU1A8D2mkrD+exLFpLYmJS0WNgtaWeFojcN1n6f72VS4hRTHzNypeVLzu09IjApSG7OY
l7MR3YMoaJ5zCMw9gytlyrYIl7oedVyOM9bXhumoKRDhSwUDnXdcWLnC9RgqrilFILKaGJXUKb+i
iYR34jhFeh9zdqYMlSx//zZwpu5MhXm+6IAnbW+TzbQMRGYmJRKVKJIIZ2qUwGVfdz2IJQ4zPsNn
hDHvZcMnd8VKFAiues5BIQUsLZe9mHrZOp5i7/eA3eO35RRbMGm+v70qx9o8z/Ehi4V+7q7nTsDn
hi3jVkv25AyCfCdbaVLN0og0+b8aU2+7S1KPyDNA36JlGvg9QlWUsYzUrYJsBDjy+RItk/u1YWUV
YZCApmqzMtL//eE1vEzGeWFAL68Ft5q8eB7vRE02bNqJKaMzIv3xZ+x+m1t7h39XzucOcJmwSlrt
x7DK+cNIF9JVad4m0tV3A5TwmUQ8dkCftsqigzupLuX4b3QzwHc5I5R0YBI5PtVCG05slSBpK7R4
oFIOXqvIhRXVUrLNM4XhSPSeq+vdrQoQIjIVWR+c3TXAROhNw+DoiuWzqq4jZBv0LeMrxi0e01+q
/tA0nug4EQJzpPba/wf80ZRAN01vI0wX7tsugSELvof/Q71aaAFwtZjbEdybU4t1DxoVnuj7DU2D
35C+15b6h0qxE56ZlkZ+s4BquSKNcBim9DNrXe8hEe9xM7UMQMX85kxhsJn4UMrbj65dLhk20VLD
D8dlj5M8K8saCPpd0hdbgWb4+c7dTBPRJTYA6Wv0Ukv9QT9vDgSuNEbzzn1vOp/UaWTQf1D2W6fA
BDTdce+ZX4658lVmet58tdIbgfU+SPxfJ0uu36f+fUc8JBDq7bFT+EJhZ0+uxZAQeRRDG4oA6rHQ
zrL7wazrrLQ1mVqbY53OBvNvfEEd23NLb0eImCPNLhEOYJ1NCbWtv1cWJvot2c8oDFxwE8C4WYY0
HbeMWGgc8xATIjLaTWgF3993v3e68RpGYf2QEQV2gU/tcsTu/jah6u38xR4647qgeQ0A8wLcH+DL
T3bfT08zTnQQJBVTm5U1UH1KKFh35G7FaXo04zPXqUrvMYDyXlaPrS+vbIkB1mGtsxWSRXY1vgpH
m6XFa9/+6apDxqVDAbnJxmTg8bzp5PvD39r7cz+40kcclagHFVi6FTiRyHaBbfAKox+7B82RR/KV
3/JFJt4OnsK05ojffqH8iEPezwPEU3BTW7gnMbK6CWXvOl1DUFf1BeU0PHlPNdbHz35fzCX1FMvY
oL8Y9adK/gCoKpeJiZ1fCdmYkNqqnw2BanOEdZNgH+xbMzJCr8A+0VmSgrdwgupbvqzVOA8t4AwJ
3xfiqCC+LS9QPrKoulebQBoa5DGAXshOIzBTWJ4eZyzgfLKWhKBm9NRhQCy5A1vMfjbdm1Eh28G9
/XNPMlJmqIs0QP+wyppzFcLch7c0EyrQXj82cbTqQL/BhUInz2KQnzkVt3KHuJzlNaYjg/YC592T
HPlIAhmvsv+rr76PiUNpZFXxFvslAfEP7KMz0GWPwHd7yrVUWx+q/FdERE5VR7MJv/c+F1EssTVX
rNVwb6CzsR7xSdWi9egn/xTRXRM18TuN+LytaHnDsk0rEWXFbuisfpv/YJW9V2yspx2kx9g9M/u8
kAEvBq65P9c6EO+WNvyDcJSRO1MFJiv/WjNds6rPBH/GBe9GwxaboxeKBXMCxhtMQiB/o+kMEpc2
yasVkXj2Ol8c6gKuPaPeXuHoauTwNT0OWU2JMRKXc3/Jpfh3KiTorCFqURKxgi8+vHMB2F2jNoCL
XMcjfen91e4+lRdqSgBBBNjgSU9wMLsBtq0hDQCpUw2zF+NiMLvXBJ+L/IZkB3KHcRh86/c288NG
OoyIFeHKH7mPiXUqtp/6cBVnpQg2KHCOV0ApULmJkoV/pjoDfSKO4Eop407jIZgd4+ArLEeuIVPP
taj8pJi+/Qde7GrtZYEMl9t3S0H4OYJ+3eNFwCl3bSxXKQEU8l+YQ7qy3lPaTlBRGJDfQz9v00WL
F3cDkfDAJToy9Tb9tufH2TubHPWmWKN3qv/7aLXDOc8QMRXd6J5JMivQ5W2FqEIveUEGNjPV69W2
e4rsje26j9xdzX4T3zruFvLpEAL+7Lbs4J7mVeNzCR/3A8Dr71N9CIA7qHOOXTOJ8bOs+JKjKwkQ
TcQh3Y/CUVm7CmcO55HLcFMXEZuOCmIPTlVqARRrjjXNnP5gSr2KQZBAqHTfd68wpZUW5a8NwiA6
qPRWs0xwny4jDRBKzY/fc3WrKCACZKw/AdLHjg1A+xkm+VtvgZSFozXJ35qzjdHKZ94LP374X+2e
TXPCbBMLtQnqbrUdRXsBXAc7CTOJRZiZdSyTsAt6/myesau73QPl9ht1hUnqX6KC1P/ymjeLggzg
ZXYeKGc7g4/CoNl3EjnGQ32FrQiZmKjE2Mjyi/RVmkHVkhUaBNVDorxl9nL/ip202ljpSg6V5wue
t1JaJffAA9PIGHQjQcwx+tjftzZoEMawpjEG4p5kj+XxuCmTmQJymn06wS0Tj6M87H1vQBBoP9kC
BuONq47YjgfNUBkYbWi9FIFf73qSXq/BsPG529d0vPGuBkRGDy5m/bWCL5sEvv/YVdWZffnwhhw/
3TigYfDdyXPz0E9yPsRG7YAkcGkrNynFIvyTUmXKBHv8i7tGkh5Magjqy/kMls2S4v6DbFmZwTMN
2N2T7v7bn2vKs6M4imZcdF0pi3ya5t1VcsGuXtdcuiC8NZCknOkqJoDaF5UqSuyzfoz6HGjkLA1H
EEwKovYEjU52XBRR5K2bq9I5bdCA90Dr+OejnQ74Rj2cwgSwUzuRf+KARX2jM/0TL2JVlVPCU/nA
ja4Cq3WYgWxlrMHiClnWBAGRyi6x35798etVAVDx6kpRmMikKmDQ7s/7+O5kEQzzEkfP474vz1Hb
P+sgiN/5TK14xKzPUyyJVP90lJK+nM0vzCF7MV0KZA2+tsXc3JmXvd0e0vnLMABVCVHqISArBUlR
JP+27XxgE899a7hga/d02xL+mPEFOJ7QW1R8ZJPyJN7vY9xKvfREUsZ0lR7cpnQG3LAc+NeqHFia
apAwTKx3VU3LyWwiF5AKEeob1vIZrZJnHPYJ4/tq4HJrYh9V8gcyRkC4wfmpq4o8lHGF0goK7Xmb
EwgFHE2CMlgm6H4CHyhh5Zjo+fpgL5HrRt4GvPcNTz0UpljuVlg80Yg8Dh39t21Thz4MJz8o+xCd
64DSnlImfJWqhO/FGHVQCbHylpb7EpxNC6E4bPL4B38ZwdYIk1nLeUalVRRsQ7huBmoWwMMlwZJ7
CZ4Qx+UDB4QiV7+WcE3f1JrA1CIN2Dq8x5+opeE+Vp8qB88HkEmNQLECf9giBMw10RXFMrolYU+w
07CIvRhTPUX8M/jp+FI8JohoE+xJ+zKiHdARUON0X3ZSIjCNSD1zubBFg0kv46DHCWtySUfY9sN7
UNIOMwmxtx72cgKd3FaX6vaLeXTCeXea3JRVkaBeotqfhRfiQ32Rtn86E4M+zglg9ImDbaEWjOZL
FA05ezO3gJP4Fv63SBRUw+Ivns+x7smaNb3+HoFwdMS3YSF/5cCsE9EqDjbaJjxtiz1lLlEmCLAQ
gxFZRmzN5BG2BsR5aHPc2JNxE42qzjPLLvX5Ebb+4Qo0LyP04qNTMW+MSCVIvgH4HibmrCnMizM7
s3138tVOTDV5OAoOa0Doz1xsXKQroAny4gLJK4uQDYIrXNRf0QU9gbW0mGVbS5/pyb0A64ta6G9A
qkw3mw7CQHvqDU1Soymmx7ECisDsMPNWctXK1qzJlKr+ru/swEHA0GrpEXI+TsWJEPh7CdPmuAf5
XVxV30IR+Mp5BlxxgBbWlZS8f9+juxvIbwBqYdmiTJUVMt6k5n+hNhOATJ6Bfuz1glBCozrys6zD
0kc6/Tt8fkkc9JQUmz5UxlAzKLFsFndBAi8ybwbU/IqDcbPoRVtSc2sIPuWP3ibKPhwwGWmK/d8a
2xRdh4bd6cW4M7TS4GayOXpV8oBlhP1rpFyKe7kqgG7sMdq6H4sll3S0mTLHdG5uwKzg4Fb6WyBg
yFzuuP0Dv5u8qjLR0qZS1dhTYBtTxkCVSPDaPdw6NXp1JMbg5r98lodFJmQcsRJNkcdgRWUPGqXx
/JtWJXzWGaLnX6+9Ki+nwQaOK43YWBAVPVs32N4UoI1lkd0tYxunMgT9lkFWmjeG/ZXIsnD0YWEm
libQCRwGWC9QZYFkSngrMhMFM02MbtnveSQykAcgKmwl4d7Q60CcB+SgIx4G3mz/rnFsrpNkJ1Ja
7rkDTyyKXByRqVEYz0kd+4O53nBUrf39yX7mSOmiuTf8SBbbZSqx48vnPi/0CotNdEX22x5DQtHw
xlDxjsVrQ55Xorewt6Z3S6ZkeuZxdbVEigDwt8t1V/T5nQGj7XP2FM25TXDulQjTeWmnV25Sy08m
gr+rEi4RbkPXgC0FQtjSKdNxTNhnu2IPfkWRQwmaJQndXXksjUO9oy6n2HWm1+LqY4qN1WaLXsEw
LyUUL7mcum/hP8qKzjptlE4UnTuVZcptAxkYh3T0CF7Iq5CKvuUHFu84crfhq2vcM7JIxo+PoHgM
JLTQEBHYyNXfuVMjYFbFcuQbwHZsyfii94hV01es1WVH2NzmQ06GPrAeXZ8tJKbh37X4886RxrEd
0hHSfdhDtKgG7VEXMjTR8L05IQA8Geo8CqCr/JhwjGRhgkJ1a5zkda0nGjkIjxcxjdGIU8tC+Uuy
hBIu6IQ7UJwueuVBqc08CLGkpKWijBWH7SyLjpSsh2fXfz2ugZ/Qan/g0tHRILwLIswaXUtYQ1LS
8U2miGlT4w2ck62JW6RyQiYQijQS9MlWZ7cqvGKzq3inkK8JmJqYEbZ7HI4pWgP2Uuo7zKS5PSdV
92mzK1AOqEL7DOanJJFbuodg16rH1/ptU3D4Lr2XBO4KzEV4z6lDUPrMsHQb2d52t+gfidgr/2JF
zjh0JcmfKLL4SSDUcyEUVvwlF+SSfU+8xX2yG5fHCXXGV0/cAhtUqFR9Mr1bl34NcWi9lQ/1q+O9
Cw8F+Hrm0HHTs5UpuDCna9linNBGF1p7zWrXyxtlsL9RDF8twpguj8jzlFjdYUpPo2Lw71LT368a
/1KCqDY1hm6TsvMvpRj+ivdQcVLmdBIrWcsUCYcYaJb2q1/lLY5pISjQJuEMnfdcCpJ0GcHfYsTF
A0lIROwNOM730a3HD9s6N9QT/JzBhbGkAGmxqUlX8e5XjrGeJvq10AQOcWZ8ifBPzuqJbrOU9cK9
Wvc7aFPZ/+JN2ccOp4kwkZAY1dFHpXXgUCbao+Eq9qQ/asNv8tng+HpvK2+/UFu6suCbpEefWSYz
fRtlRuti/5EfP+OwRxu8Sb2afEAJDRT1Tv4LJzH6D4rVhzKR05qcHHFQfEb/vvu+YEj40khz7Vv5
acP/5cTcXALE3Flk/My4foVwKjIEbnK63y2ya7tSZuSqPjozFKAyI+DIkdQ6l5KCHuyuRQd94MfC
PuihIhHbf3X2g56MajjSBv3IwHtq5R+9n573THGoJrmw4BP52CGBM+IEna51bCld1gOZyVakGHCs
dlTMQKwt5RgthjLrZksCNq++TDELB7zGKHdGxtkk6mw4/zZwe9jkvYW2UCl4tzEt9lgJdHqjqQ91
Hox36LlZCoR3ir2Z0IclNhUsgg6MCmS2msXZ4D8dPi1oUGs3DtqSckDavt8OIO/AueagELWiFvn4
7ITeRJReiP0CiXyNXfOzz4uKn0Ff/+B8MA2Co52ZNgjWBvbwfufvuCckK0SgL+1A2X7N8IOYPzCW
WvZUDGssw1jVDvuEjzkh9tps5HMXl8pYeqljumjcB9spqQvgAzl0drNkK7dFCMHtnTaAp81t42iG
BQ3khk7ub7tOjGM1GAIlFTzsvsaDLRy6KifBWWZlNkrWS8DxEnqGdAAqHZkA1F2vYLICvGusjq/i
gvNY84/RXHdaiMFNCswb9U9TzYPowOKL+AH+48JkBhNkmooBIin0B2S6FrqzpUr33xE/3fSY8vtb
PPamx0gB/wr2XKRoRgXPlucBCOz6irCr7nkHcuDFtSV/Io+dT/ZMIePanADMmAYpxBSbTdxb8l2O
xbke+CEyjFkkn7fCRmsFbKbwuw+2dMBstX6Rm/JW5otDz8Gqz1CRap6Xf6X6l5W1MtsqKG0Gidbv
fF+YhkyP+lq5/hm1+SLVO7O8IVMiw/UeX73s3wzU0aGSp6XJnbQul8avmDbaeWY2M3A2/PUt9YNy
JTu51DildyHkoPZVRqBqTjmdRnZ1/bulk3r7Q7vP3/a+vI/P9Pj2vidIsYDjQkgRCPv77Y1DZCv3
d6HjErDD0xlrZDzG0YzEWiE87ZpwY5FXJt4iqhP0foMmhj+Eza0zyxqOJNTbquXmglVsHtdziHPQ
KW2pbP3wvPlJ3pb95YrIW6Z4K8pxO4nNy56HKMSZV1bQGK2+5Vzo9xW5T6RckbvxUje7WPCxzevE
jMGGf0MKaW0Qp17JOxCXvf6REAIayXeppFYf8yIsbJ5XvpWZHmMQMtJ8WgJ1PbH9zg0MhepxZpN4
wCuxvca9iVn+tGVCNh1n8NqfpQidhn+jGIYFLXYCRdzYI+RGReY7/VxKvK4/A2zLhtq1jtSczbxi
fw/NVeBD0O2lKcmZhJI4PB7Yuzb+nBpBU89VgdvyAOPJWH0KAFNEI5ZTI7mfqmtKTNBAa1uyMqpl
GHn0F2cUy86ly+KyAhu43ulArQYTkOU/dLHmlujJTjeX2FhI43rzBKmx38PPZUfdFTFE1SPdqMmp
loYyo5dnKxv7AcOZfs0hMmhsnO60/83k8xTGxUmmWqW/0ZKJWTuptRaG88D66KcnYDxMYvL8n7/K
Dk8cwnt1o78TCNMsGQh1WzUV+s1jzdSjW3BqGSNs/dRdJ0fgXSnlHmn/vHiEV3EWgHTm2M4I5+1r
K2RLy8gLhpnEWnHikmQhGeGxT0Wljl3NkD1fuom0mn+1VBi3goQLwSi6DS/XQ7fUAeXz32rmfE+n
c0dWKm+idG+VaMuI/ibnbAmH659fngRDfktaWdpWru8kMhc0lZDaCEPu5PFGzNdptTywuPYCySr9
wUKlv+mG2nfCh9EtnXdu7Cvbh00bk44iJ7axQFF/1Q8h25i6mQtLqa23iAYPhCEqgz8JX0riEeM3
nz7GGvpXOi44KbHlmcYUAAjCn0cqvRUVVJqf2egFJRsMapQ4ORL/Ki4P+pQ0eFG1+ShMwHcF5m26
zT6pk1h42XgiD4vkTc6Mt4vcq+Aiqq5n4Fjs6A2g/UzAGv0qSpQp8sqzznkgwlRwZAfMid3qZlfA
+YdOUfH6vTeZjmmBTroHfpS5mlxYLjCQU9WsT1bpbNq5DZZ7OkLPj0CypbwkQZR3C+n+uRyfQdKP
UH0xduBAMjQnjO50Zm95HxzJt0hlCkys3OVV2mPNm8y0aOX3g4NohLWVoPhlqKDoBQbzUx+X4Y6W
zHQ1cInUrU1QERBCKGOhMHZOZF0Mg6ZQR3ogjgZBfr3hCKFkTp6/03t5Mu12DSd6iWDJSIHYgpzB
rp2sHee0veYXfR9wZN9XGpaYlpVQWW4k9a6/+xWnZsfOQMgw7TbpBGWBxWl0aAQoOXN2VUa+jJAS
5xo7t+67pKAfoohthsZUXcs0sWwnqkD5YPtX32MdYJ3GUSDgXp0lfRXDUNrRlfNwcW6C3gNPKmi1
FUgSPNR4O4DsBNIZHJE+JnQJYbNgcHrhN3YtnPYpExh2xuIJzapzjIigrmucnF44Cj1qjwKbM+52
VnLA53l69mw00W4A174hR2JTDk+9iPR195NYVqGBwZazg3BIcoPPbeRnTRAClcKt6lDE+7R8VrdL
a0ulIC7DJZwEpnz1AKrEhfgTvZX9yRKCxHm3fIya/j47HHz3Nm2AvFSyrU5nGhvpl3nuS4I8hKu6
ErnHIBz+d8JXeG2e/Q62FY6CyjnoLG/Vp8CcZdxfh6mFXpJHy+3Tc+e3vxf+Auq0iqbW6nxtX+8b
S6cE+3VVL6KhhXXKwT1Dzm+PWqUQyMMlSNbbKmWI6GZU3Z+R5jswM3aNtIyVqLxrhkZQKvadtHHH
PGQ+G6e8cJJSEAa9tOFkxI82JARjBm1/W6tWlZeD+tlUs0xQsD7YNFDYhOpRG054yWDpGCqrp3ig
Gf9lAybCTTMtO8ghDNCucStCUle+jufkpUpXgwmjSC6JhqK6xRe7Ec4aZIIeJl4g0JQGZBB4C5tf
54vocrMi6t1z4eb/YmFEu50U8cPQPDXRcOOoTRF/Gplzi6zczxc0Qpfzy7HoPxQK/Axkr1mpwlNh
cajE8IPGuT/1Iw0PLC6hVEIni4MMvQVBZo3o3dW0EWmJP9InLduXyCiNAqWxfavj2pv9+I3BvSQc
QBJqG69ruqXVrOqPm0BWxhZaaSXWqy4D3x1nDGo1ty1Xm3z2J9Xk+2P1+2D8JuU7Jsz7PYgEwgMY
fpfcdVaFZRHphyyPXrzkBwTukp2QoDr5YhDJ36K1yoMfb/czjbsDr+mBoODppMr1IfgDJ2JqQjEl
O4KlYAEAQ3j+ykZ27v7iu7pyIKqsmAXsY5KDoDUEk3hE3UYIcQoX5v6m6MUbDiV1P48gB+Y6anA/
oJBaFmsM1nTTjbFaA5ZgAI36H3s7L9p9QKfR1sojCWfmSaOhOsiMQlUNqh5uhnI0MYKuvt+/SppV
KLXyj1537SCk9r6OSHQc48J7x39KjmFm+bqt6Ms+LOWaKJifJNMTEtAWFMrr+CKmiUsYKA391bli
nFksljh7BhC71lwB+56AZbAig9q1avqwIQvM9QrNir7LK4/g7IooiL5/+mgRh2flfvfiq/Ms790k
OVk6bgpL0J6yfmCkr3JMQB9S7NjGMfdxh/802BpxilFhn2/YdGOnXOffk61i+x+Whgvu2CdaC8fP
FFIOedptp8G/FVUxIMWOeMJrzutv3HbctafwOJdkB3VpM+AOqNCNHMgzxn0vambCubaf8Gl7DD/W
6TN7xfDieP6kxjwhTXOAirPzTrXe0TD93lEsykpVsLDSzjPRlMlktEKY8r2HNAsL4WmujVlOo6Z7
NJtoA+I1VnksMwZQUtb5j6GhYOeH+M4Hv36fJHx569eNyj3Xk12ASUtKYvpIIP5te7FkOprRgT92
JZpmwYOG2aO/ktq2APu8UgqOWsAFK1jJx7oIXRacBma9LBIMrCsu7WiAgHBaNYeddDfi1QE/Okmz
eI6O9B48wjPQ/TNvopvRCO1EUFWQ4P6TY0A/37itBYDpckZGTUSTf3alCTZMyRZ6IbDa4ENXXqqG
4dVGciuJWtBc/fB0dzqTmDoL1z3/Y9SKUT/m9v7HfYCwIHBybINYDh5cBw56f26fLLOV7kM2kkNU
gcrW1LQeFpOHTewlf+phaAmM4TXqP6GO96hfCdJ2PiiDFxU9oRxXCVdbJEEq4QVUl2A51YhKMnTY
5o9eT1nte/ySMUXF+S5IWKPHnd+vXtA6RXNAPFlsHIEUrQAdopKmmxr/fct0t8YdAff3R5Q035FV
HFmnZpn+l85vQ7z683bYjCmvgPRM2U1x3LK6uX3fTXtc5x1X2DSHAho5mO9KZ3UWbrDn67A57KPR
olnfezbvBChutK2PlUbwi9CtmbMLGGQWbIPIxTwvW5zDcVOOa3/5wIdfD8A6hxuUzQ8Ouyvvnc/Z
kq7NK4JdobNaQ+90UefOkZ9R0AgJ1UW3kTY9xAHcp0UgzFYpCVXqfE96AfMkQv2WnWL0OcVZdrKd
8dsrGA0ff1vUnvhXdmxSe35GA/CnuHjuz1M0Zg8fUJVbrho/CORtB8m/cqCv3m5QSnQaYa1SBX0C
hUHO+9lKrJLgmxl16JwWZWSA6ICoKh5WjYNaPvgjwiqxV6S6DNw9xvXZ80zBAOb5DOX0/JFFZ6g6
AeQvsCzVvvj3jJ++TPWzZ9o+cWD7YWJ/VS0Z+Roq3dUqH3xUMY7u9JL9aCY7ruGppDcXpAFYUnKq
AaMxj7fp/DO22kLp66gJ07csPt4ZIUgxl4trs5nR6gK0OcB9LenkcIJSOlG2bXhQBXAgn8t/EOgV
BB48B0Bq2kIx1rY5rleJ82ByyguYqyFL2CrZcnrooOSx2RnAJ6Jr5ZrQl5DY8ThvKEkrJ7hL/Xey
r52iLaxaOaG+pJWYaKXaZLwVZH3vOcCxhg8fzajQEBwfaP7rQS/Z0aWbcOjapk2QXjib5YpoRhGF
TGacP6TFxl04vd78ePv571wjD2KGYKxEPG3SSVWaISZ+vFIG7Nyb3KfdGsorWXMcD9oOu5M/RyzJ
u1xz5RACWAaN7hKAcYsyj8ckGyFbBL7foKUN8IkD+zdYmeRFkfPguBHKXx4LmD7z39JbosWOXgqo
hn7yEB9rIxPkbw3NeXF8lgLFS/2249mlHC7K2BWcLS292X9snB70xmSYIvU/xwgPtXwjkO7BXWLg
C/oNUnqGLg63NLPgZ02vs3eTSfueoVU+etBCUNXpFbiR2LGEx00T0f/ZWlwSnffN1vbHu8PpAqEe
xflyS/CsUwvBorhhwTFP38zQMquYiCyV7NuCkLGY7Gs3C5lfdv6vor8wADgN88//FJQ7EGnsSusl
YYhFJS3/tsY+8hVBZx1zV65b7EAvwbggLR1OwI9Sf/qmqzTcOnOUaJ3c36+cmEodxfTAbx1yo83k
vVopqK4YNTBjHMR5gd0pu/ySW3tm13tMcm/QNxQNKlpm2X6tLdTK8YXvyI2HYA8BVQXuE754Lp85
b7HeeOJthtB5yOX8XT/usXShB/F55gsOzGIqy7E9Gucqz1qh9w+okhU4NJmK3p+UZtiHeuJNGKL3
8/c2DFhDINeRRv8FYlRZyn9WtniEnXx2LebPEq2lNFiYFYeepmtbGMxQvHplJmxWUMhQoOIa26xr
ra/DkHusManwZzJiNhKuUEt1c7+GJlN4gsHX+saILm5i6C6m5Wc4+FRh28KqrwF6RMtCqbzPu/Oi
82aNuZWfNoXEUBYZ8TPsEB0/juqW/jNr6mYqlbnqcYOwCvfj3V6gm4HxpUu0rEj/M+QusqSFsI/P
EBZx2La5RMSK/07igCF793QeFWLySN3MbRABU3TsPpMWeuae8mS/UcqnqHxbvyCTGJ4ZnAhdwKRf
eTC/K3qctw0/IQpDYdeuXF6ZvdBDvsWr45U9kHMx3XAmkE2AHOR8lxf2633mfZkZmHSb4Mk4eh12
J1Ep0Sd3RYLLqK6VdhJq5vpYvDSvjLuqZW+zR5nvO1+COaoEPvWgTQaWOHaJ1c9cyNObH8jM3SY6
GJJlRxp0lYdj7/HXKIEgNtL0UPPEMZ6eWn/Djsp8caYx9X1jAbzwFOO0MGPwNkUAoII9YFLBPPES
X2PUnVhubeS0v8bR2Kof35WpwHfith0bKARgSLTG/cJqfwiT+Hv4znuukXZlzJYTYH2p4vO6tGKt
nX/pvC5AZ+/n4N6wVJoEKh+QugrYytUdXvdB73LvJ+jZx7HlneC0GuX0Uhy7Fgp5J9vaBzVOCrd6
VJZbOGw3pHi5p4SQWVpKFRypDUW0pr2A8Qa1n7zA4yELzqH7pch9SUnxRsyg++5DqzPrHOx86grj
/QPw1LqgMLlGkC788yMT3AwQjAyTMuCUt3RrVYbmCSncnr7D4AtF5vOcGnSoLt63Q+GpwjlVRrmq
g8N5xq7juOpDwau0jZ/SWH6lHu3iK7lWn6DrplpfIu8NGFexL060IjmEZfKvEfd7E+d9aBa8j3SY
cHqyAVK2MfDKy6bKjaD6inGRbHRuJJv9WTscbU2u5V31Q/oB5IpE0njpmvem2tfAvka05v8WptPq
hd2ap/Q8m5CrD+t/Vkkuavi6risykPwLcUgYcYCbJZvfZ2AujEBBh70Vm75JIyFtDCDoIJCuWqG/
dnVqvX9XyMfbr6T0lwjdOGVdMVxrZwp1AHnxA2RLkZ9CBQwekdaT4E8nmi1ykj4+q9RIpTdONu3X
h6kPUJvouXEylffAzKkIxIF2g0frWBnvYlpf8drGvJyltACrPrUTH/mcjtKmCMrZ4Buaa7wPpnN6
QGgSNZAiqvyFoGXvcruAE8HUtqinpVxRw9ZFFmmY9uwA/9gEwyNKkO8SVEWSv6IBYfz7mL3cLTyV
/fgc/Ksp10rd8O5Jq912sIHDTak3l+hIRpJLUcr4Y4iXoyfpQ0L/oCbjqTeMrK+rwlw8159+dfQ0
PDw7MCgeVnAPArRVQ1ZTpL+u22fU0vHEZYS8U2hs53rxqAo21flLti18BVjJlOx3UId8DxpSIOnk
LaWfv0u4WxUIuFBYyDWYO4alX3+9IrjPHZKLxFwQ4d9iX4MkA/ySlcrMDXSQ5ewBzusOSjHRutmu
tyjnMyTrYNqtE39x/1kgEqSMEcN7Cz45Dt0OmA839+eb5Rlsr34S8KbIkHKygW2kFTZIvULGc/cg
kofKs640BOkfcExwva+LnXaPa9WNwYLKBINi7jw7XqoNNte4KcQxcCA8w9dGT+JxYa7atDM33H8i
5Wtgxj091XINxEwTkPtlJ4FDk2OCsHA6/qa1s0Tn6HsIN6QmGmfRZGsyvXGzwtV06JD+QB6lGldM
kDGcODpeSmPym8vGc7j517ZDFqYjK0uBIILyckWZ0qgwlrcEZEWuAe4oZhMT6pFm024H871JzEIz
SUfxlmoobHffrrVaW8LIWB6t3kALVBQTOvF1PMM/4dnTR5Q01J6/3NMD59LrHP5Clr3RaIBOAp2U
fo/1TG0a7HFT26Dx9E8buQZpZluwKxhKzJvHGH1h9YIqhQgqeMUzmV/zhM1gJquKoBImtAJ0lDRi
fdyuIBpD05ipjOPBhEDX905ZoKjeVqfctS1+80pttk29wHJo9ofoImQiTdQuzQu5nH2NC4Haw+iU
OHGdz/LCDwz5S+B9a8/CjbkuDGESeNBwxzBIkvUzxxEKNqAaFooEnRTSKTex5KNSFj7v+gLj9zcs
W0JfvTqpQRbmQ8k2kiADggJxtLDqZD5m4nMaMnoa6fisrzbgpPUX+c/7lvRvCL8twNQ4umqx6tYQ
a0Nv9UovdMQw6XqZcE3mC5EXpFNj3gZEjBvaMaZZbpyID5Y7P9Mqs7XTp3UH5QRRIPL64RnTBo3x
DiSH+iU7whDNgSl3TKKGa5QXPvufmNtoT4UFtLU0/YLA3zUwUnFlRDnpXSV33/ScLpC2+ssE3Wvc
pvD1nTywNTqLNNqjtZ7EIWjAyEROYb8AtlaiLE1HLGN/YNBantZF14cMx0joffxQtzzJTi6I1O+n
5lxKH19HhR/ss0DPe9sgcOvGsqHlEVYlzoQxY0kETokwlrSks9ok0uhKsuqlr22nKtLHA7ayvZLR
8XdGy0sBp3zd2cOfj7T79YU78p4wGbFYTXBShryyKzH3R/RB9hZ/hiUmINPwzoOqh2s3LoE5sTQX
oiAoaAyyZ5nt1S9A9Z0W1EVR7VomCU/oQM4XfPd3QAUH4ZZ362g/+T7NHvv2GUmvwdEkDRuHFPnB
MCc3sQG7ZZzKzVjKXafTT2KUi+qAz6Mt5Ti6o6rkTd249JthpkvxXRqUaO4XrHBqWS/ZmCv01cSY
C/bUQ11AVn4s7oXzyGptjRnuzfmbHjEo5z8eLKqH1oTRI2KF0+Dx6eClWNH8zTAWR8cLcMpNkorz
toKFIfcZhBXwvMzOBHEgLYGTzPV4s5Iit9kb7YQKwyQ6J5wiKyfIKubWSKbZm1hNl6BYWcoQPCiL
wOvoDHhQXrR3a6l/ipCTAyeBi073Z2ytXPBiIpNMeA7561kkieKw3eapmY0m8a03olK9M+tr/z0I
uf0iblIpZE4ETRPrcuyTWJZ3dwYvOfFFhFeioC8eMHVPNlQYHMT5QZdYboWFRAtKkrKhaVOFGBdd
7yk1ndVVzV63WrfgmVbdfJDed3AN4YTrUDp6gvIDm2impLxLydft+0q4HsWt2sgQUSaQwDn+R2Up
AKAR7/2uYD/uqkdp8gLqLfzGJjROKlx6QllMlUcmsaSQvsYHN5f5TWXeF49WGW2VFJXanrHGIKgZ
JXlHX9TjrmMyjHHc3cgDKyrc6atkXVBSdGLnprIBk8WlSIg826O2Zqm0bH/pZyVQSGjIvJRYTv5j
43mdMj6FqZFpR7yJfK8xMzAR8ESnd98uwNDzNsX6RLceA5Wb15s59vlM6ncDTkayfU6xfT9GoJpu
pjLK8gC+bS7CIRSicvPEvCv8C1QfCERm2cFu+Uzw40kbsTHhZo9zvn9QqFVoD1C8sZ2RaMd55IHH
UuezVnaFM5UI3JyL/9Mz2T4L4//K09+KJMD3gC/+zonfkoCNjwStpGp7jdu5g+NVEnn2Rzeiw+y7
jn89rdXFFTnGUYsUyVAUngdfaiy609j/uM+CyRiv8nSXtgsLECzbaCP3HZ1CtDcrLkaJOjuBom3s
aGAnSMVQl7ESm3h281jQDxuu1/hGyn4dqPHCr0GmssHQ6yQqfm4Cse5dXr2ZGRCqB/Q+SNzFlqdA
VfI4/qQqPBWGN1oVfAxRkuMrH5SVGO/RblIAHoX3zBpQNNbs2xcqTwKeuIvsbCgOJKPaqWrq2Ox1
Ty6OAyrE6smE0kAyH31oWdzofeQV9J1spDfNUOm6fo8v2gUnLaDWlz1Ux0yeH+qA1RJmkWoACHSC
yJYBWwMWtJoeWzOJgtdD9ai8w+DTc5/Ibkv+OrbEY+SzMFv+2d9yj567FWlbyT7+Qf7Chd66uq2t
mA9QVstEXboFw02SlvNxK06pDjibcRQw4qacmeZBFRTC/wTvWfY9whiGuZESflWvEaSXJNRkpxAH
CCZfeNw2hu+g+4hj48wZcPyK5OT8WqEPBn9Nf+V+NxxQedGMRtzClNrdhke9EN55bbbErtmUzXjk
erOgA5x4lfprRSHjp1aeYluEwDC7FOTF9iAQLChsJUlLPMfED0hm6qbEal50H4J29KlGVjdOAjas
UXmb9r23TvEaoNgVoIXdgwNgukQbx2CYtRshuxhgKkIExII+H5eVZ+yDWbJ73B5yvbYeihBizRYM
Ph2z4nLaBY0399YKetG4I5BzW5/zPUzn//+BaCscy/z09ca5mVvn20u9mUkUMglEvBllBp/cT+QY
SCu96ZtiNOzyYx1wWeuDpwsA5CJzihoHjkdMky0syYan4PMAFDpx5fTxM/dTpPn918ZEuVz+fhBx
lAXrDN3+jRNxCft38JamERExq44sCBlZTMnp5NqjU3XsO2YKp8MBJhEkW7nMEY9/GVlbDX6TR6C+
TbpUSnv1YmM8qY0KZ78R11Nutqzmx7IdevMEziCzGhuJUFkw+Be/LH4gs+4JIEDfCb+dacys7zTL
1WcFJ3crenGf/ByHF6wTM4rVUjdrsIINulhgJpso1PSoeKZwR5rbCBcANiz8aCKuYyuxTIdV3WQx
TKQnpGxLm2vWr2QPHEvnxMjdzt/Ae5KS43C+OW4JJAUkA7UaciFhlCdME+zS8tDmnFeFzWDK/1UY
zPEmzxbVVF3SgHe2RaxSnz9tLKPp2Jh6gfYLEO1Sgw+DWEWZULopYiB0NCmL3kvacxdK0QebsG2Q
EsWoujDvIYZ7LAWkU+iSHhNGaTPh8rjCRaYAl8iugFNQe3cTYKUcfUvHQxOrWAQaFoWlYQNvnjcL
hNW5ht9iYc4GfP/b2GEyYT0fzX4fb9j8phdtnWpkqfkb4r0zZOeacDXjSsfZiY+dWMGUjj4e6Etf
D8JSIh+zl5gx+eXDZX07Yy2AO+Oej2Zr4KVGqedKQmRbSQRBulX+KkjBWZmVV75cRGsE3Gm3T/+x
fb/6LJfq2yBgXRid6ZQ/Hv636L2q3vGuLEqPSnv56/uWTwGye82VZHT5Rqk/HFyPqFCNV6g=
`pragma protect end_protected
