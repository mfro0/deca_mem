// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b2A9D5kmXDYzkFgWq/gM4ejQ1vdz+iBsG4I+Om1xJiYhOH6Z/YI4piFm0ib4KgQ2
yhPfiyn/q6ZyJBJg/0Nf14h+p9nEiYE2soCuzHWToo2ajna5B2biokV7h00es6+j
WLjOd3PzKzNBIE3Vn4wLdLBI0r5B8D5Z5wApEn0euNk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13536)
h3YGs6LN31f3wqTbnsum2LsSwLfqM7QUzgqYylYMOQoAy1q4/3ra0mbkRizgWeHH
gdYygj51+GqpJwoFqAO9ihWN6iy4qIRAiuSFZS8kqhKj4buWR4f1iOmVwbc8XuZ0
LilqfqiU1UAv3phvqjfMPLUIHBOPaDmCBtF4hyz5bCt7sSBsR7aI0gehuBPVZ5LQ
Q3G4dkie0L1uL1Gh/T6eTmq4xnA1bnlkpXjd97FaLGIdHxdDARUBV9Oi5gStzubI
CfG9fg76LeuJ+rXjz9AJdAMW+UgLqJCoyN0ylwVseAW7wnkFndh5mzb1BBUpVXyh
x6Z5KpqKYhE5bgiai7kOKDxjFe2zriGJSfbBTdWsQaB5BTK40K4BCYDW1RUtNqxR
ZQbgZKa2B2lJD6wDeTiYooLxhgMccE/4+NYbTKPJUhM7K6iMfq7k/b9vm+Xd0O6u
cJ1HuiSzYkCnqOfHy+C+SchdXrm9PU7OfpLHadaDwmVH7fYxwHGqsh8waMpm/nX8
aa5o7JXrxmVp8CndYqOyzk266bzwTJz0BxHZSiExR0efzoWhZrtho5hy0iZCuLZj
bZLGC4LR2+mu25sk/EmmRAZBPAvx/pb3jci98p3aqfy2Copf0glH4f5GgtYwS4b0
fI7RgclMbwNUtmJCACC3LTSk4ML35WCN2Jyswp4cyd/zHVIuq4ubVHQXsstUQEb4
xjLPn78MmZahcoZ4SWVqcUW69Oz+cAC/efFz4vLWrRALDX6o99m6WoYbzeZluIeM
bR/chkB7vY1EesqlUtW/un81iQf6PPrwlO5qOJDzZJ2GPE28mTDdmiwEuxF4lo/2
yyOLjVbSMCkCY4MzDF3Zm8oA4P/kiin5TZzWiHKdiNhQWTwVR62oTAibsrOLpdW6
L0GVMPlhpsQlSz6dncfuM9FiRdze6IcSTqGfKXv9il0Ke8Vb4xwb8q85heioYolQ
R4QJQ77KJTpoNsEVfKCmuntglZMSv1YzwRUFmVGSUI0IL02nKsTOCmxnmPgF0/H0
Ucv1fo/LnPEV30//9a0P+msh3Vop3D4WRRqsm+A/KOGIY1ZnknSRhzCYlxunW9W3
fgT2iAQlg3O3a6rrOpBgUnibJWi+VBQHlnLhNmH+5ISs4w1FhY2v4wxuUifUVg66
EO7BnOiCTP1wsyRiS9QgPFXprYI3GSjQZbCCFYyciObx0n6AStOYV7WHPVPciEVs
TRFdzvaZn02+6XbFJlorquzJ4c9j5urXNO6NT/F17eIcX1ikp3gX+w7VPq6r3Do4
1fdQD6X7gIhATT+AZ3eU3ZqUIxe1klB64rIBtBhqEcUlBu0YfY1dt2sVuEKkKQgT
c93STcwyAk/oBfuU6p5CHt+oHoATRJbj5NqbsqYDKJB1mORVdICuFuGmTdI1KKBH
oEmImmhUPuTE4UMojbpTFBN+NqBPSCt0PZMLFnLfyE2V4+hanGs85+ctxPCNnqgx
yxZ95s3Z3f6ZCFTGaulN5mva4QqmYb5YDZyvPIV6uuRbYM78IEbEWdaou2N0K6SA
Q6cNnmJyYwe+hK6CtUh0tTkWbnxh7GtOP8fWWyg3LOrBlcIfG2hlC3BseFySwl5E
nrFQ1rqPCYBsdbKD4R/N04rj67wXU9XOAyNLq6u0zoH/yukLx69bwopXp1tHVLXG
MAjwbVvMNan/YoGz3iogbVtagdsNHRCeAZN+GA6oX760kyXzHhtAOLSypFKG6Mki
57vzH2q5NpDyeuGaKCbbRmgQJJCddrx1V8UvURcb1YahBLmDXL5OwjQfAvulw/T5
oD4lc6ZziGeMh19vl/QXFUq5ornfoT8URdecbNks1MsxbgpNBKvl1MA+CuiAbiHD
WqnBk48CecBvgJvVdbLquDanCaJjmX8meqe3KYf5MQoSHRInjw9krHK2UmvHB5ly
D7d3GjGVuazzVtx1X2Vz+mQPRz5JQHx5hjnvxF/VYr59W1nxflYtI9BhllphMsyi
BDElu5L0Lc9gyY62ig0pppQywK/buvT6GIdDSrgoc5VOw+8GwVBXHx43Gpbx5sZQ
HbGgJvRYPctXpz7lm47UqeXukJJFTHvmcmO/j/qquZbhIDO3cCNIZRGNNwaQtB9M
tMJ7C3VuNjOVtrM5Vc4sq7Pn4RJYwFtbn/uVYqL74I52EwGFOO7OEFXI+aowlL6f
j7cFHst+cMC3O0wYDVEdeYKhp5x5hrYzzZfkyY4gXZcPDWNp6l3faUqO73DExXJH
JDPXiCDZrtTB4R3WanzOEQ/QyFW5XjkO3khO1id6ldeDmvziPNj9LaXuqv9ANJbg
yLdcsP3OxsluqSATkGXMD5PXCiTrDLg2NvuR3POaM6Zd9QhWWUkk2zCiT9XXh+Za
kFfdZopRhLTCfctRvfWWu+BnKahyhI/eRaIpA4xVyzSrTAdXpbzhIktvF7AMVtXm
7qfdT0Fw6UKfqmYmoufC0yu1NyHDEhBnhwjvE7tKzzgZrdCzYPsvgqbOcQEd/f3Q
mq38XcqlTVo6oPjawxvhMJtFnQFIJS454IPwkLQeqPtbEfMZc4UYf8rTBvPRCq94
wrIMH5dhi51vXycAE5Ydv4NVrOHnxlvTktjkda5Arz9CO/MsX/2upjeyhAw2M/TF
pXGIS+BFiisz49lV2e9WQ/cy28lv2Uanv7b9twck5bRQy5uqIY0+AyVePW7HJGq9
/Fa4yEqFLWm+9if8eibeovCQZcBHMbqm4h/W8niJUpswgZujaS+asZg831zKNElb
/SzNaZBsOe67q9TnTJx0DQuyylB7IaAaTvICZfwkvRI9lLbm0m2pIevykzbO+3Dh
atUIizchQrVSBKuKGbR5jplRi/TnvwLqNqtHrkbwbdf2oCp1dgsxOheHqgyymb82
bRXhpedZe8aVnRnb6kLT1uc8z+2hozNv+X2w53hGUr4e9GlephYVstZAmX4+z6uX
Jx7MhBgsgb92fG9qZNurugLBnU3jg7lHNlmB2BWThcPpyAHQ49q+4RUOD4ADkDQ3
TOdHu3Ts0hrZStJ1AAEXihZVvf4zVHNjOWM6X23aEYqWd0XjmkfqZFvntly/MmK/
SQUhD3aRwWfoqsdONzskOaoIGQvcTqVjl2x8bMrkecm4LYWOanxTpuf0xV8TyBpn
TkraAlbcfwPekIs4hpdR1o8p5Yoe4c7nd4/mBD3vWrcTRaIFrFyWM0LcjjVBHnxP
GvnFqtwSsbKMz4aTub4DwSrXKc0Te2c6Y1dXSbf2gJpmz9tfLqA1DffFg058HH7I
g4K+OgzOZtqhkoaYqws1rc/Kjea2DeOk/Air2qOT1R7dM+XCN16Zst04lt1kbZGL
IKM8Zp1ftITv3degdrk+pS41IqB/OP6xEfp+4bhOKCKqIZCnrXzzH3sjh1iIHDux
4G3YxzZix3Ei76N2psowToIYql9PYoKY6DGItOGS3pLqT7j4n+/Cl7CmOIqzbhJc
eizxfB729Krt35dhTCvIBeXxCZWHHBQNd2b3IsS7V6KxmM38d69IKosTguLB/u4M
aZ7heCYQapRzpgfb8jQEe9Mt/XwA+/1oOh1e2H8ApQUMQSmqlE5h29g4gNxJ1w0E
wZG1b6ZbGK80QF/GZCEToCJCv2mzLRE8MFhlAr6PT20FvG2lu/YFjIAy8HX2xMn9
edtanZL7Nhygt2A0kJrxAsr/3DlPSDObMXgpcwBZfbmfxUu2u960iXD8dI76LNe/
ZjPgT5EQI3S8k9lOGkVzJJUPFBIrOk8R7UqmcBRWxuci5Y0fvKIWSyoifKxJu9X0
sfCn7Nzq80GHWojp3CHF17RD6BHYODKhbBwnHmGAb/YU2pYHefxZDlVUJUEqGPy9
wn3wROlXf/dlGdVozBfvvOiZ5N+onE+Yu/afJnj/e3DOBci2SrxjvUN/kPzowFvq
nfB6yRSkDEkj474O9dnKvq5Sgo7NJGUWN5RXa6xyo2yVkjJWX6VAX7JFh4p6zmt8
JopOEqlIt4CH/nstNMwsSLeA0Xud6TjAA9OVJL9k9JBPzdYrBcgThZG89O6pDXNI
IbMcaU2G5Aif5A0q5Yju6OU2aKCkaEzGUnTp9J+3YCKypOq92TnHb9rGivvdRf+i
siEN15ntqkwaZAoL+PFTsfHB2FQzgvwfojhCOprgGJJLcy6roVeR74oy4gRxp54i
bBkxqxcrhCTGKtLkeklwHsOEUI/ZBeFfFb6+poadcxzmCndQ0Oc4DT4x84JnvkEB
JOpdWCmbZYMSEmT/qxkYllkI7DiPjyWCUOzX7T7CLUP1fjE2rdoZ/H6LJWofWTMA
4KMBTJd9Ee+ULqgsDCZKabr4VNZktNjZLiz6RXDBe6asgeigHCrkYgD0ZAuDrUjE
RsorXmDk/yFjcQpvnQRP19PwDQl1/xpYeblVbkmSTpZga1Xhrk2tqcOV+TnLIZoa
p2WlryYNEeMAgR1CIvWa3VbOFp3l+tIS7MYIXXdjc2Gw0jNpLqYnTyziS+5moVGX
UDo3xddt4mrPaQs/UsrZIJF5iZnDR0pUS9dsGUNet8BVnwnQkrBW2N2avAOJIPlN
6yNHK70mBCCjThH71XSzJxmHd6/909YepKK4HWVDG+gp/uOoZIClwp97yU8mkldf
2A2bu1fEciolAYQZTo4WDl2qZtLjui/9HRi+xyewxJReLBffQbY34KMHEWgmn//P
F9xBXqRDReVbFVeySFJOZUCyabBCTNcBGvKv/M+8ZUICmvhZHJ/6VMI54HjUh/hL
b6ZlpMosEGloOeHL4u8vx7Uj6tY5avk4HvLoQIZF21cs12eYFL06PSmhCVFFvFJi
q1OA0JAOITwt/mLOovdXSLbeIgiFjJIuNdLYX35aa5oSzP+OulMz3XVqgkj+XUjq
w900KKR8frrL6Ub5JIiYTKRRbJ5w/cGMOQS2/dYB6HV5fFs32mKV9wi1SPADXfpK
QA6FuXf2TaPDTyVHhmfg0QiGJeVWpMz6gOpIxPnK2EqH6fIaqCQABpoPZ9KoOiPK
T2PTcjnX5pucMZ4xKigXDp62FnFdTsc9tkhqg5merr/YrwUjAt9RPKzuHcGazwGv
5yjukB4z7llMxonevM0bsdFADhL7ZXqbpYfALK/UPYcuRXc92r60KCS0iE0rzZf9
4G59JMQDNOylrRlMSgmyRZB1DSRl4VkNy1tDhjRq+CNowKeEj9jNCNhHUPnd4lGc
TtINxv6pvgXyUL4sD0RYQaAzutwaFYWDtngAQqOWkL+IR8TUSe6teAqL4tw4jOQv
nzPTgQiUjduCLZyAv2mWBtOqLfj+hQemOnGACn2MslY5oq6L/zqoWOEb6nJF1sCr
wdDbYWpkUzNem42LuLI3ULFRpDz7v0HzulrJSeoyfoG6TYp/2Un7juzPwVE0xFDZ
85Njy+ikO+klfVoQ+2Yadpw8hh0TUs9UuZ8AIVN9Eu51nyzy/DHR9d521wMtSWM1
q1pRs9EzONSqZxht6ECvI8XCif5JZki7NOZyaxnWlR7JkUu9U5CELg9jKuBcgKc6
pIY32BwowKh7lapeVAk1nEAkpZtsSd3ZxwkSaoHPAEshNyiVTmnnBf+0KvSqwxV6
xjUveJbboHjeCYZCCmCowmlMLZ7eTzJeKb/Uwq3MlZBcLIqSnalOc+GPNB2+GkvP
SvUNyfYa0G7no5R22DZMeFSiC++MCvRwRqIkRAsMBYfHsmMQFZSYbG9b9PFuF6iR
7t6F1P39/tGD9c/jqY9iYBtiln09b87SZieLQ7TImMMkoFUCbQDjOq82QN0PTpWr
2JKcl2SK8kDfSauWpUEPhGDsF7tROIxhsQzan71DPflLZAUN9soeME/DfQyRPBKX
3YZMJGT/tE6x2DxUO9eJvTS07tFQZOnd7gLk/n4xj7wA0cgBWFnXvPeGNteJMdqV
o5EJXBekim2qN5mUjj7xUdpsh6KmWODdNJqhgeLDbyTYiii2nPadZygxYuLDyowI
H9ZnlWjy/Ve48owpb47Znd0GaK1AntUNPV7WePZCiYXYckP/8SzfFQBDoZk4wba3
psPGTGpaj1+t24L104fRZ5PjCwZxa+Rg2dkUgiPgFrnBSD3DxblfCrJEQgVaKs90
B40VjM3ULQNVTsUwSKtRlqgY7na1bOMK0OzeJ/Qgx37pOTe/4MtB6e9tFF/KnfnR
DGeCUUD17B1sI/SKU1FA8yP2dRNgiEa+gmpD8HcobCFh4kGRJOiKepYNF0P81C9p
zEnu+cHvXO8u/N47FLvaNCHnHC07aIeXzSnhA3bJBUpxBmGHE5zpdMde1VrXnAeW
WM6CPHJd0RkeU8oBJ8GlUq/XosdbqXdXzL5AhYcvyeQ6nzCzIFWqRK5tC8fKmv2s
QZEuLrMwLMvqEGInwYb1qfChoRg48OX30DIMjYQ/zc2CMvDYvmPlMGMxlVwRfAxj
fRgONRleQjyYQIPYGJ5FKS4+1jFOpxocbKxheWJCLLg1xaIsHWEoxSDo3Jnu7nUd
lDhn4J8pcWRVjgOorQkTZUpCb3lqRr2v+f05RCeeXamhfI/0hL/nzXv+D8GJhCGh
eAS1heczqw5ptdotoUlkeS72NH2ewf443zCO8TcHEdpfHGuItKpU3CXJRvQcfeNZ
8H8oJB9yTMdoIXEZ6GTRz458Cc01ekVwe6oVpLS7/J2qAe+PTdbdUyf32Qxbt//q
ocwL9gNALkvX/W4kHz/X3bHCRwr6lwaKHAQ/TEusfkvmD/CzE1QNhjdVhHrlm3vI
dimYOUpoAehHeEaHU/gh6y/PAr7R3mPKdyyuxVA13bFMcCpSqdlqSWwwC9LfZyxC
aNLvbvA8wUMGWFVko8oL9GHeuvIvwOY1ekxZYGFv5dQF+orHmrGTQ2Wtm2GrFw0L
pNBrr/V+P9g2BR5M4Djx2+w42c60AmKXX508CAO8XGW4y+Yol3FCSn7sA1ZGJze1
1o+3bkbsn+FFXiPyuAsIA4IGuPe6W2BjP8I4Ih8Z0mLUYYIXvviUe3AYcY+zKb7N
Xr0D2rz5oYXnznh6LOz20V6RCfxEPO/BE/tx+6otLaDy2Qhcvl+kcpraqqhb719+
gVkoFxwbFuYsb6Hk+pXTx19i1JdMokBpYWG506F7AoKJWG4uY/NFZR32nqEKPf2t
vDFjqF6BO44WuskV4oZNR0wiTjYxpuhWHsh0zEoyHn22pTTy8KeBmzk1rFMQNMSx
2x3O67OCJaLBPh+2QAh6UIyZ9C4nt1ChEeky1kj5j7kcP+pUmVyukf/yiTLhT7QP
aWMDAPuL80oVjaGu2ks0zKBGAfMnPgMcMLZ7Hf+Hxz0a3KtQHwyTvsSOe6PoPsCC
pM56hYcy+mGoDsl5Q0pJ8Lv4s0Z9Epa6cHsWIXp56Sn6KoH6bYBB5oyOEe/M1Xc5
uBY/GUh/x33X1f7KMvMH+RIZVksOoxF2WD45nDygCZhWHHrc6KFZwVfRhWikBsk2
Xo3H0LFCOHAw+JwzOIitFTJmY2rO6lAMgS1gPdjbtO1CTjrKxoXpdIViz7bN46Fs
DvWL1ZGTGLY+VbZL53uaGh52uMgmfi46WucsrZec2P9Ur1DJLCxhSC3xFi6Tts/2
XTfyRKqXKbItBCqDNtGEjtBTfvUhrhWFiaqn3JRcgdBAyZTFkV9+a0Mo3F13OO0v
Yatthg/SoMMAQQQVvMg0Z7Ojf9PBQJotmkUwIQNQza02yEWr/yiq3H8kwXhdvuPj
DR6E+PhVOncvVngFsvb7kBjYSqqL+JAbGaEWGmRTOcrAvxkh1LeYDRbP03PgpMbq
wfEEo80VpKG41cH4qrp7m5+24mcbbawPLe8uJvaNyoGKb4tijAobQh6008a8X/ZM
fz84/ZZbUsBb5gJe4jeZduNt0llP7hkiXmz/sMT6/T+UdnrP3jQtr24tkpdkqBKT
YAGIy0kdTOxrfSG/nmxTrl0KHm/ZaKmqJdTycia/yVsAnm0k+LHE1pNEVIu0/f6n
T3QXxWKgMOGQXX0ATTfibZQ3c35YWWysVT2TcAZDxRUX1z/h28/CA8XAVPLelbm+
71/zcfssF4fDx50BHY8k1iLlBIgapVYPADLOKoiFxGr38L9HICPeO9McYSP9RXjy
f+nMb1IqkKM6GqGMrZJ/Rv4BsOJwjwuibNIDm7QNVdrHPx/JN8nPbC2xFk/vEmbF
3R8f7lS9My0notD9h5WjSGvuZvt7X7QEvvSbNFHSBpUeZPli3kO+aAiHxC6fR0uK
eamYjM3l3b3YSkT5RSgZEV8bLHYMw1L6Vd9wmF4bKMLR909AnqqhwXULa2jKt8Ou
flsH5ZjpqmIqF2U5x3mTL43nnlf1mR6LOQVho/CixI6y7ou83jndyblaw4Nd5qGR
1J4UbRqvJ8b7tBI6GTn6l++NpZy9XMK0gXYxx+dvCxYbJKUforURY16FVpVyAukl
yNjeBMMNzaKhDLX1jEj4G89mbwjDTpt3BQMWynlvjb9I/gI7Nnek6G5o/kprTbPb
fYDh7oUFso6Q2bnGPfERsfAAf7+5qneunYCy+8G6JcL1uvsWgXkh2RG7K76yv+m0
49p/DfgIPou55vHaWjnJCfKXN/gfsmR/5zevSAokBIqGL+K24w9UQKHfkwEsaH4b
qF8Ubv6kU4wMGMQWiLV1cqo9onNxGFiq8PUAggsk644xjqRmYV0YvnzygW4I+5vJ
1UoI9TTpqJEKpK+gzDkHdtAM/HGrc9eexcx0IbTYaPba6VBB7a5b36VRVdubElkj
5VHtz7s41UqxeRuHVUI+k4lL9mezKN8+XSfg52vmdBisg/Mz+b+UxW8UtDvLjmIg
wCJRHoUKi31CsuKJo19Q/K5q4q1S765bxjI+gme/hANuxDWQbm2fIaDE8TPrUPNE
ToJ9FOhVXKdd/318+2TaevqIzNLjRphfju8iArJSuyZMYJXAGCimwgyEr6Tnesfw
vEIFj2j8dV/S8pmrarSCZy4HSNDbfR/WybMYTfv3y+iShlTYwTHbfHu+sRD2J4Pv
zCqhSjCa103OMRMAM0J28pTLo9o9uIRMaBnFdabO+a3WHsFuCfM7BTJ/RxIODSjz
RgzsXdC8gjUIkZoUE5W+UbdbSQRpmqzknqS6tea6mRMUJ5HfuJNwZRH57bmsqOiY
FDlFXJXswTdFStwwqtdPaHr1T+SU71jrsudIqHCMa21ZaVzfcVgzxQM1xXnRkciC
NQ9f+q3npls8SNP3tEi523SWP2Pu0iFWTwLW1eUFXBBjAYpXCxboSbBWJv1PDXi3
/sJh5nrn/PB7w/wYT2J9jXloTo+zJI5ICvmQmB/lq0Xvoj/Uc/7YxkGbbV3RxAoZ
/+XhEsX2YGd3FCI3VEpwyjn5sW412xSr2Ho9Uk9AkcTnwalAn6Xy3ESxBmfkaQtU
F1DbTDjrB+gCLf+8+uziIVZjcA6A+bTLy+2cBIEW/846/pKyJK9wEUIy1EKo1zTU
YUQEGyRL0a6qjb51S6ZZGlOAhkhosXex19CMDpZqV4BAjcRcX+kNzhHtOxvulC7d
4rQXNh2d+6shZVCfbINyk24BOzoy5R6ETxZkPFfub+tbWI/j8vDXt2fs1boDDd26
ZigknB51E69iTK8Gl7KQiaDggxsvwAnBhjBZ913jMJhj1x3NbJWSUnSf9vMFNJ9P
bJzZdz6jplL6bpg42jYO+I8CI1NIq1uqULaDK+/khOY923HF9+a2dA0hYv4IptHB
iMC+aAbJ5bTBG7FXY3U7rgp8Yx93NZ+1JbEniTr1IUG9Z6w9U3UcrxW5UZbOUQQ6
vgcBhZ1PCCrTTKU2Ne3qYVNFPthhqd9c6WDmbyo+TqX4Py4RJi6gSQqNkn8e6HYl
6OT0QGAb8qU//Bxm1PtRUmMApJodheNOillao8TGyPIHkWtOz/JXfWkzkAVRiYLe
87yOY+3fD0czjknS/l66TV5ajgpbzuBEqqT0WfEc69aHpmkFjXdi3ojKw+DKM+wO
Kvz3U8jDEckIwd+smybR/kCnR5oVqtGRvCWKojkuf5dvsmS63IXC4W2CLMPN1nmh
rigdVmVzgA5Okvj7Wb8OFCJY8LMfkOEFOcVRnb0cambn3lFwmX7NfpFXlLgUaQSn
t/RHZ3jRPM9ojpVuG+32e0tARvFyjBb/Jw3iYgGffUW2G+TNO4rnMEfUD7kGJ6b7
w6xGeozHt+M1TRCWst5V0v/v/JJFLc2MbKnF5VmohUo9OGqIh8+5UEPBYHz2ga56
BtChqdqzLHXRzwEAZSAJF4FRZ18+rrwfwqVDRsdNc8NV9tX/MilGbBW6T6R3ODH9
DVEoEHKA7xXJ/HpqO0Ie7PpVrZVkBunYzlhL9VA54qsHNCW4hvuI2ZRa/gFilfQf
1b7B6/8cIbvbhztbtr2naq4Yz3R2N0eToYTR0/4ZE9VLQjV9oAJHuv0Q0QQ4nvww
YoeHNYFLHvcU9USP8Ac1Ft3QvvaN7ddy+3GaJ9wgaOP4Z5Rk2Nb70tqkmdoxw2eA
KSx+fjgqMWnTAyWrOJP7BjmuoNMcqqPy13Uoyax3b/ty1Ez31uVPPJUY22KTbzsP
YvHM5k1QOFmN9eWUTpXdfxr7MyJKBHQWOP4sE8+ACN8vovFZs8qBzquKSLEMAck7
mckgoG6wbE08TfdXFHyMZrtYGKjbFJvNgnXEMRFSAkItDecQGQ93Cgyl5vsb5zqG
ABfAaf8PofhZ9W+1GqxyTtsZmzSDUUpGv1DvGKRo13tZuMu129cQqugLe/7QbqML
90jzdaB1NP8p+/A2j3N9BcyWDTGwgzllyHwwo7gUnFF7k5pmvuQUJqCJedgwVvQU
y+0UTS3EFj+pXfHIYqqyyGuXnPcNHl3xcOHq7zw2L1OeX2bEd7EaEkzS76ChQ3Lv
E8zeNXjlTR1B3CFX1qrekylaw54HWE08p44IUQEtXU1+7FRwB3PRHdaPFheoqkKq
Hydr7QdSeTOp1iq9QHm4mPi1nRp9YFgRVbqcH3TqAMI0Tn3W/wDp6TIgxKkxCG59
r9gxB6Bn0xh236s0I4eoYwmyqowO2BeKdTiZ964V12GOK67uJuDPQUq31uo+7T+C
kU3EwVX2lsTefilBrU+nnsRSqqtydpixsZbqiXBzLcnIDwxGnvr4wwYJFK7Qu2uy
Sp7lFMhvJHx2idtYaGzFdrrUJz32gPpCrElOQy6MWnoTp3Oh7xQShmmoAVKdALh/
sczmdi7B3KKlgcC0alSnki0fXq05Ia2xb2DeXfhtUq1FGbX4BEhe+9MThZMuYQ9P
7aXxVLCMjgj+gnoGoqptvOuNB4aX2ZnI2Bo329Jh9tq4CpEwdwo1fFZynKNIFHyJ
pU2564GL7c3s1C4Q9hTTY32yG9tqYxI1la+cwiB3+Cox4n1RlETlN9qQK81fIEOU
OyjsyxPTjWC6h/ocUhj69lOtuWwaJ7NlWWS7eYotEXfD6ylanjtsEfIqIthlBlVK
HxBt7n3ua6qL2V3i84KuIGunZIGxoK10VMkWbH1cG5TCkH8TA3+iIXZk7ONhVy9w
KR1pYVocuh5kP9R7VFzDmCPVgfEEKH14cbYN/su8HLtDVnt6dFI0/DNJAU17Mrdh
NC87030f1FUJxAZnUHnCRmbiLgsGkcei11GCR9vTkc2AGcNxRrHUUIPYmV7WJCNu
877WiLgrR7y9J4MPLiYpohyB3w9i6p0KxQBVnvf9p1yH5KIO/2jC2uPYOMBmAvW5
0tblDnEy2MjV8HuB+1XixqUBbfci6koxdgfpUBvaHc86k+CfDEIZY6t3+hrocQSn
I1BTZrcxWwar6Sckde9+Mu+mTRpeiAKzMrrE2RfNS58Z2bx5gVLCLAIif+869CPa
5KgJIsMF6XF4mkSA4KDDTq4c9Jur6rorUhcQ28JAa3g5aNRnoV3Eq541tuhFyj2G
e4XIDBhmvH4D18T7qotMzCLXcPpCFNfhQ9NLaOabwmLxmLXmMKo0FxtatJP5VQog
fi+fdDrk5xSyclXIqyu4ZJUPK8/39+FCmgYAxOJm1x1k3rimWGqqoNjw6aLoikfM
7rNA0T4zLfTGm3Ol+JrPiu8Lbp9vSxlYwWS+yRoBrNhAjpQb2ZQ/SzovxMNrfeKj
fFobvYUwI/sEi7JLQLNvkvltP92yAwBgCriLRAT7/etD7TtVi55ChXZ+D4+cE+z/
BPKsiq1G4khcOxgOImFsMh3nDWWbh8Gn2RxSj3km9/aTt3F1hVnl8zf022lT6csH
9hS04m+ktGOgu3c0Ia5ibWt++WvzHbmlvRH/owrkq56dCnafReB31yTwgdm94oWc
JxKtKNx7Of4QywRdfJPvSMwhU9BA/nh0pGN6kzZFsQ34XcL0GUehgqJ0OnICrPNV
ppn77Q05kVQZ6rYnIA4srMZoh2wrR9Xn/771pdEWFqxMx2dDoHeqKBN9lxhwj8NN
KFylDAzYF4dyqiWOPHPx07LMDGgDFV57LyhLfHDjqFJh6ipipbMeb/WmWS7G8BNO
v6ubvcMMmiOSSBQV+TQBzFDHBJIxvwfg0yiJuVUr3Ndpa6n8HZOwQrmuj8ylWVQv
urnueM98FFN96ghS03pi2ccKa6kxBAIHtKfHFdzdB4vulc4vfVXdbCRJDWPJ0k1r
A4UgDLuILebQ45PDvCZdOJmpQ8cKaQZMr0md3kOxlMLCiXn9poEYQDqVk1+Q1YOa
ehbZUqwUjk7KQidBX3SvoS/d9LytIcxWKJbe1MgsK+0BCiJHmxIXAQpBLVg3SXvK
SlWOt5tlDtDp8B9vMoZy1SP5FCDgHku7TiCK02yn2F1w/BADdwI0nVEmPDQRPwbl
JN3WdfKNSUszfQWyDX1UN+PIJ5m2ZHWqPTyr1D0HV1NLGIZ8cIH71c1txgVeVEKv
oMB0dEu5NdAuxMnd4q+wROkuKXifA95tVsDu7yBVtGtJYVk6wP3tO22p43J0czMf
qgW9aVd4J2LO+B+IFI4ICpKAvYRNUkQCGeSpaKUUo9Pgs8FN95e1sNpByta1oPba
gIn1ACObPWRgL3Dv4ZrU0aSs9wbWM55AGehkQYRYisoPq5J0B/2PvEPyN+zahhFO
ZdDxwp9uLlG+nL7tEMMM5iaBzKOMMndmqyEitgxcKGVLq8WHBlon2ugOnxQ0O20V
9p4D7UDhgEhYh0Wr5I7GbpAVznOZsN6o9RA1jpKg74MHJoQmDoDZUb6PfQT/+TZP
KSMY+a7R1NK3Mf1q+UfsymASrQOMVznoN8OVlRFbJgfqXksFq8JLDQLLqq9WGN6h
98EwCbo1auuypOIHQOOE8s/gUxpOHEkBhxNMPRitEN4s32WPHpqFk1rPAdUyDYZx
g+7jo6erw1DRmDJeuuDSBZBudFnF0254GTzHdk2z8dMn4EhVK0+9CNnV9Q79yTfm
XGbzdQwrOrlf/sLlTV6rQubCISlig/FTejjolOMLpgM9Ydzcx649XByWKjLykzRC
OoS/bIP/gTi6OOcfFqDLKj0zbJC+VjFkd0Ca22p14rhmwtXIo/LB6OUXf3CWeVE3
yw52/8SfU3E/qTUT16LH36Szx0qCHKqSmkDM0mBXwVUlNqDgm2N8ZJOMn1gftCz9
vrxUApbgTVAWiclwZHxnryjQMnn0HBka7uGvql7qHJz7dkF9JTgGgsBNWeBJMINs
lsIfsARqsunnaejAv/aaf2664x/ZAD7KWDQ7rqYAckXMCaNDY37ALkMZyUMk7Rs8
kxQLRY/zBu7RuqpZOwlrg2ThlJSpdr6ntgw7aWEiAB9zxGHzMc6DL+enp1Qx86Rv
VRhchjBE/QyNGsXLq7gz1z0PaPJT/WPnHALciSRZ9GQfFlYm3jACkwZthLbz2tdA
fhSsSTzj835Nr6RjDqQpQ46Y7eTehKjzL5LcT6kmDIlrDZATSKz5H6ro935NiGlX
uNoZpZUx/bqWI3W3A4bYfGByh6vBClP7OEfudxnyfNl+dk6Zc3Vcxm5YsPweJzCj
m248ms6ajoo3Rs5k7NzEbxSmHLXYnMVugGaZDAtShc2FFtbDeHro07Qk1nRJjXdY
0DA2Pzwg5xpUvs6UZolMlay32wC09r03hkA9JdV4k0sYEeLnwaGkksm/6cxq6L5u
6bpT8T05PIx042iHmgPUMqJRyJZ7PeV87aJxIdRDFwlt2YTp6aWNtjLh11oNuZU3
L9yOcYrJCA+jQjUC5JBei+EmfMgTH+TIyIIRt8tIofssMyTBUxn+k+CxeoN9mkUW
I6r9690d6apVoIYkkJJmhZLjAlSDSM63Y4r4D6CFeOBKddZZmfDUvwPB8z4qtrce
UYmCxcJkI7lsbnEJG0AEewuZvTZtxly/ey2J3h60wb5uGF4Nbop6bNiFy22te47f
bnxyccBrk8j4Jcu3hnkMo8gwg8wRMtbpQmJOkiQNyUipsk0nd7N4dmR6k54080KQ
3r5nxNH469wlX42Zr3YhiCTn6XwDizGLkklLg9wQT4IcFwCJsyUmlnUnVnaeLmpq
EESU9ciTxy+WJrjfooxsFIGoafpo65LZMRkahIPATb6FyN+KVCWHKJsuQrsYbNLK
7uzwvIrjAJDSlXirjTC5s828HWJHcFFq8RhIAyN2Z/oMEO267KTyVzJ8vycnIfVq
GCW9eKy8gNK34RdEGZPiJCrPbfGwOkh0YBwKAeNVLWnPoWZ0Rl2j01SlG1vszdgO
KY8fnvrioGKkTetyoH4AQZ8tLPdEuO7cLyV4t1woJjH55ZDFG0pDncM1LaE5TN6P
CeUVol/WBZSIIva8tnIDJpLsDJV2gLg4FXNRItbXkN4+qkJGWkZyAhEb3IBncyE3
QXH1bI8EQ4PpmkEVz8YR6tLbWLXmFJzoSZcmKNXZtIBgm7kiKiyU/7G/8IidX7DH
C1YLX0FiLf5RS6kDZV1QbMGq3KiIQzBQ2tJNWHstG5eSqt1DQO6qo8BPY69yIL8w
vP7pyTD8XLU4SK0Li7oORs4J+K6aSsfQeQ+zhsxG+Hw3e+LYmIVDSXbLPb4WD78j
YxXM/ADaWBR5rmGSISmXkApwWWQlCeyh5tzF0u0qfmY60g/u9mgeoqyFRt/B9w2I
z6piOlEb6PWxYBYnkF/BF6J28dKxLE3TxTZWH8jhS7FyIaU7dI/Xae5tENVUpjYM
6zItOgiAa0wJo39kPqxb/jd/VlZ6TDIZLHuyJCc7bJwtu1xEE8PlP1nWDl5TA0WS
+4ZP7sbSL8eT9ogNoj4hXmIAmz+Gu5ca3W7igQ0GPIVG7vseccE1EMZxEgVR3Dle
4NHaifwyklQ0MRibO5/6mGqmeW4Y3r+HKAjZluulpN1wfGZRncp2nxE/I8lvhEqd
PbuisrgQgHkgja1mvvEzZjM3/4a8U/nSiipImpDW2A9zAxQ7wA27qoSW0QIFEtWP
V99ddsVN6JJARBNNDZAkJ0irPFy8hqHm4XRS0W2zNkjui3nH9ipDMaUfodW2Vyi5
gYft8GD76MLf3t3rgIQooAsh4Th6t8GJfUg4PCVEa/oe21bj2oeO/ssFbp7kmOIU
0omcK++e7i3F3/UF7ldLcExM6cRtwe6UnSJzx3klvKHOLZm1XCK3NLpwhElen7VE
k1zzeoBXS3cUfrEr1a74Ua1VvQ+FaHeHiYRoKVVozNKmVJeRA1y+f3jRjKmVKjC1
3kHxtZnGrStt1QMAjcKo3UdCuqPmL7eAVbv1LjeAMVtC2YBJw9pZemEQXtBGMVS0
sn56nJYPeL+m+19U6Vimcbo4QfD4a6pedb2wtZ9PUgfHv4n3onCyg2NnJ9tkD221
DD83KloCID6CU6XiaPVorE/nqMxSdJYWS+Uo+cU4PjQmJN1fn/wg0t4BCeKoZvHd
4q5orQevYbBaZD0kNgpkfPJvS4Poa/OoEEU7djWM0U8xgtNmIrV3jmOfbTZxrSNN
pvS2XqQBFTk+Eu0gUz/ziFoXgBPZSTGRW5M8W9mSaNPXF+IV2Ssgipe/woBV87Ps
P61xPiAaHrB5NZIPQnOul1TPvp8FsNKtQXLhi3g359HC2zxFCrZmlAq75A2fCM5d
jnWQRrtarzOiZx0L2LDs+QhJfzBqfLzsEvDyzc0mkeEpB/AYF7uIc4Map2Nb4VNZ
JLiLd3/ATlq2yKPRG/9mgP5xinmvm2enEfNcJ2jgUM/xM1COEqJ7LL12TEtMUxY6
JDue8pCMh+/YVg/WIeWrQ+cZgTu3BC0xctjbSPhyHslsWBbi8O77SNP8S+UZenGT
DmMZmNQY+VaG1qnC5szidsROzeFy3G5wvZxoX34lg0MUA3oz24ih6ufBwcFqaCPv
as+yQnTSsCOHUEANZgmEvDj18QG0Nrb9jZa7R4hxwCwYudy9slREfVmxA7Gpd/I6
lCrMYa2MkUqK95VT5OmuopWTUKAEZZNBbrWzv+qXv92I42c/2G19Mfn1Sro+d96o
+fYfwu3PKIljPCG4DWWcVpLrJNphoAgbcCNhZWEhiGWwPbxIqLLpnuNY96i3nQmE
mwAmWi4GN5NPQWLC568Un0OmOh0upE+2emAaxItFU4MFVS3HEEukKoybtJhQ8G1R
LDGyZy0uD6u9pBD/arkm0f14dvnQtY1iLic0HWnU/9qXTEjgS/OQmUAwQUSOeZTp
qkPviUxW590EsWN0Vr503CiefOzlHY6B6c1AReyENxyLQWdkBI7oT507NVq7bcFm
qqPGBWSe2L2dTA7WPkM3TfHLsWrlbHAgZckKPowJt6KPFayr76wvx5HnHDM/fP13
3VSc8YldH6pTzdoHbmNtiYjlBPkP6S5wCUsSR/iCQ6OgiRyHw1ecGwmrCr74W2ee
FZvLGlPO/9bPoDBNi3lMUrX/hC39FpXlQbWw/WKhFjRh7SkLhbthXqoSLQfj9U1c
UP0ml8upM+vcrhwr6GQqXpxUvCBtmO9Ydt2HjC0dyAqCRG0ii1lJczC6Uqpt7AJM
MMcxVh2dtI4md8FM6+a11E15rNvYbcpW0NfapA/apGwdoeY/FygCPeKWUaCF3Yh6
RmgNetKhu5jrBLngH4RTaBNNrDVARIT2cJ4+SGOxXT/EEXsDTm1jU+6HhAFsoHY4
/jw9i19h0kxdw/KXPDxJest1sP7nc21XB+miTMfVwI0ICfE3xibg3SIkiZImyje/
qxke2+WXS5WCYD9IsiuQ5K4Ui/UucUrHjCumNdOeaXTUCvHdyU/FYqqCwAzcWm/b
MUlJywIggXF0jUUn1UmPlOktto0mMXQxHHKEZDOORFxdKIuC6Ld+ZqwduL/ZFaGT
ebeEFRD7rhVXC+rPpWcc6XIBuzBuym8g5HirdXrlz/UeqGvmL3Jhvt8AvEcPnteQ
3dWj4uvIjvCOupPJeqU7CBA4SA3enne1zK8Fqh5ckZcRtJ1EeRRFL1IuGm1xzREb
PcEXT6W+MuU62QGxHJLnhMRZIZ9UAJe7Vs0djrBOOPC2CrsaMfjDX4/ZqAwcLcMi
v9EOK2QMsE9y2UNYmDTBXQEtFFUOJl5wV0q/xC99+arjRRB3+Ch3dvnUNZ7Sd5fw
3oAhu+WqDgoyn63ntd/iqPVV3wxu+ro5N0F7CKa13bxNyFej2o9BVoQnz33bLWlz
yIekQj5J+NubQaNpl3xAvCthJBpCPXagKdQ+pxWNZh2Z9yq8WvQSNB7oR1Zf1pJc
Ds7lAANr3n6Zlj/E1vYcuwSl9rOqPxd7WussJkoIEnv7NBm9UQmeK0tEbKeNuklH
L3Xb8XOZ1f9h3d4qCQhKor+wXyVUkMDyFMgrvqNK0PGZHr07sviZ5ni7Xkhun+5N
pgrePIj75njJiNoktUGSHW2V9WPvoC9ipA4a+GDWA/6fE1L3pQk4sZWl8UHjIAd3
e6PwSgeyzM2oH5m51SR4TfxHxi25AbtQwM4NjIX9U+qa4iBT85KwBYTax9wTZ3/4
WrVI1peX09N9CH0WVRWlPZZOEQ5A3OUPHN8JzhoQXaSFCZ7T//GDi8535kAJ7U1Y
42/oWxxjNFlz/J3MvpkHNLdaxpBOwTmrj/b2oytA4oDu8P2MiozoJu6XcST7xVEq
Ma/NT3LREZaOgqk9bkNacRT8E8xqCY++5vDPjZgRISoaxvMIQF6tOUFOwVykOL4K
513ZIif9Wq3WVMqN2A1MJXnVza6jva3RSsOKd+OyXR3JQZ1sy0Tkbo2uxDwIqv+f
`pragma protect end_protected
