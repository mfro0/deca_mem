// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bkrdkb1Uh1JvWxBQt2Wz618sUsrMNvbdKvuqWMspmv6jO57T7NmNIkxNcFsVZIQS
7FPhPVW9A68xhwGyXi50SgWiEC579F4rokddNdkViJi1/XDD3G7SJm/GWA65hbC8
bL5fI9E11k5Uoll/VNKYt3aRXyE443Wh9gtu5ZrUrDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18496)
Lv2PqQN0jAmhU0mk9G/lX51NtMFqyENe8yWX7OHjwnWv8ymQDMxGubzLCcvF08qI
raz+W1AA7bfNwJ1aNHHmix6BE1/69d+pPFBMKOio1lueuOO5JA2mzuPQMVkUC9i4
ODJ289HL4eTiHaoY9KJpr5NHPLxgsJUCsuc5ay2X4Nd56KYu2sOm5H7cfGcJ0DTm
ud2WvqtR0Opnnj7HIKFX5CxwGynsbqtaCCLmggGBn1M28IYRrqFUY//ZlvY6Amyn
pCIym6PiKq66BJW35b3cgYjxgGkMyadRgXujZC2AD1aawH7QYH8a0p4CcZW/1cvL
1Uksykuv3vem/NdpCM2syeRAt2NrCfQ/Ke8servoxdJW7CZzBQCkTTFC1Ty/C1KD
cFPCOiAyjPU2IzdVwu7JwfA5mL51cRScNYjAMPPz/I2Mv9mn9QRylSbj42TXuoyC
i+bRYF+50EkRPGKcWrDe5WwZ5xf6hf2csPqqTBJzdzrCnE4KkKMCT3pculrcxink
Zm7Z9KpFUfXBiZO6u8qcjEiWnt+Cm39bQ1J3icc62wO6PWBu0fXPHz1cnQ/30eHM
iuGEiEIUUSBwnsluSVRPfe9YPUkBXIg0jv7oNC4hF0t04tk4gjxpP78ZEfZbSuKH
bImwmwqgi8YF38+mEyVctqkYFDmB5FI+0jw8n9Ji5lqESwtDXTDHS79q5pxBohMq
K5tqULgC0h6vac6cGprBTWON2CCQwT6FzipEAKpKXBzB5TXnKjAz5tyc+CpXBqWf
GDp+IzTbOy08X3bkX1JBC2aK32w1wpbrHNY2U4rAHUJ+3mgWuOOjw4YM5bzEN0JD
fj+rKp037whdsJ45RHp+asx4AuTO7EasDRyK8DR2qUe8FJU5FN3qtnFcAPeliUxH
Zz/+qHbaRHLheO22NUGFL1naABDdzhyuedFPH2aOPRna6pge1u9bJTicDEyh7PFG
GAkxz0Z/FCo1OfXeX+x11+AoxQv1xqKSpJnS7zdLPalW/yfGMGed+PLW5AiJ8ned
prTBQ+Vf3ye0ZyGDMPSJAjNFgjiF/BXFdw5N/zwDEPDmUiN9RU7QrGje66nMEypS
oUhznJg6EdIoTvh6OjpN/bYMhQ/KNJAmxSdutsPzpW8YbPOmBAz4lLKBAOtFOQJ4
U/AFiZoTj+LFiHQ1XUhZGHsb6EG7OWz/lSTOsFbhk21nj7lzgUVc7Z/NGya0Hqvj
pEiv8hxfdbolpBTh4XpF8CXELXOh1F1/LseyfGKQEf04r3QXRrXGvdW2MZVsIIL6
qCt+UQy5xPIwyZPk5HR5UOZzSyHVyWE9cxrFdiVtZFwGuvCBQ+j2WtoNygxCOpBV
73jrwB4vnJJVJal2tVmNBcw5LPLgnnyKWV9xN7bQ1MRnaVygFvTcUcQ0GeoVDiyV
q28gdHJziPjhuZq1/kUoPFDrNrHNq9H9+mgW16quGy7hrp7OM0vqBEJzInhpCyGx
QvQ6PmnwXm1eDh6OStZ1heNI4651Ojaf0Hr3YU+LFJfs5END86uJJgjlfBMXUuY2
RWq6FtyRP1PgVLxxLfNU7ag97RKJ+fwy1NTEIDP1eOJAn4BmLwOA9qv4tACF1+kK
4JTujYP2QBrKNsbd38yZDIZ4JVXAklPGNoYYpYnR58v3HF8ptDYeS3HAmUK/mQSc
57gArhejLbUxBvGPf770xjN+ARhpPkyWM3FNuVQm1BZGuB5naiV3IQzXkRfpWwQ5
kVxj7tRw4+aM91msD2ETYbLoqnytLIjTwXXPRBv32ZgskWXtujGCSJsc1RFlLv6n
1frFSJH1ZZ+wu63nnVvuonQznjwUnCl2eJW1S5mWn4TPnGO304RlO/3Adw6fi7es
AOUvYmTmqT5dR754RWLM+m612cwcfhTZ5DM7AHikaJ0WIwLuDhxgsUVJgDiLq3v8
ZZjYQafFgIZ11IYogf9lPk+jxS+DBSxaPUpynMk4r3GHBpd460YzOM3k132BGGo/
eoBmjmWSXdyps5oBfmCENHoIjqt/mnGSUY2jzCkU5H/t09OXPXeD8KuUfgid3ThQ
4WWFFwQc7uCctqlB20DK5gG2ewispaToQSDPAE6Kh00jQ8cdIgWLLPi0FMUBm68D
S27Y6FvEb8BSm298a5ooMPuvLwsZWK9MjzfPW07cXEDZSEQPsDQZuFFuO+A8wGqf
jirfgNlri4exmPrmrDX/okPxfmQ4s35SI83cvbG7eb8QA79ixow+kA1NmH7tS1b6
ocaxpIadDRYkMNcNwPV2xz1Jr9hBxlTNQQ/I8ukfRIReIneZG0HO5MxDOsyWPIJY
Ny7Pue1SSOTFw7nRcRHw6roCpLBNX1UX1o+bxsUnFGrfc3kB6Fd5te41ZUNPUVl/
jkW4zhqkShHpMJCz7QzylOn//kKTF+EWwqZO9rZG/V2coYiqEV4zWE+SJAKsLWOD
RAz/9DVgzl6qH/DX9G3J3RjRFm9uwsexCUP7lj23Qvs1pK0J7DDf96Q+E23HImyP
/XjDlOyEyPG2wqUoO4MQi2unVqeepyEN96pDu8C8gPcx/VQcoMQUiouvMKQ6BkSP
LfKSrhjxPTwxpNnmfzwDjoeDG/d4x6aSs5ATKMCWilgIlQvs6z5F5/yNq9dyIhSt
rz3wCkPwuJXSjodVAnUFu8EAzlpfFLOnTyvJNWhZMFKwcpMByGGLYqe4ls9UiUH/
MCiIf8CM0i1lFP/ZAr/x7DEFR8PFudvD129rgQ4aN68VEQUwY/N5ZZ29snue30HA
prVeiVqtR9U+B3TNlD9Nadi/9qSoA4MLZNpC4hjYn3CorjOB+4HReya1UTXOcarg
ZyPAokM1n8SPiDsFb80USkCPd7Ofwtnnbt9e2bxaPpjneTVluPWin4NUZ0agOmp2
WGRkOF8sU3tG1kPNxXAK42ZHIjO/FQXvHXiPKLXDtN12zck7mUlTnP6tRdTqoxTp
cn3J7NmZPbvxtG2/YkKT1/0zbDXY2yqw956k7vfTlXR58C72U8YBeahF85JBzSVH
RzEYTdRQHoRjOIkTlVggUnkbqcmdUnu7BSwv4/fnJ5dvn7zu0GiiDlSaZzvSmMDc
Pr50YV7F/KT6RKSaIiDMnhB9lkHyCVOi6OQ+eX2Sv+b+C3FEUPqffFe9ww82rBBn
6lwrFSW3mHTaZWgXtiYEhEhamWR2Wq5mRVISMX/PpVeocCPeduG0Rn3/H5htkro1
WIp7pNBw7OkDawsJx8e40FL6zVP+VaY7z+5DsWUR5MYXzKFiT6e2aiGHrC+BXm1X
qslKoNMi8Qy05C89rDFsMaP7y++TzSerGSMIIpyZ2Iln4oaLvOEMdR5i7dPAHdwQ
gcLryb0ZMVwSrTo1DVL0mnaXIl70WsIMFjKCtP+eM0BKBdsa8zmcy8lhDe0ljb61
8dOq08ct62vjSk+JtbLHq8gFQs4WcCguX9j29/fm7KRCK++3p44O7diTEn9wKLur
zuWmjN+4bMgDmiTVjXgjwW7cITT5v6JW5zsqfyWR2FOsdANLnwi+3QgynS3iXkOk
5YexQMlR4OV6CB2MleMKK8qtn//XT1U3ki1/tLeyLuHh1d/BvxQUCPuo5SRi5S+y
ipnTS+FfU8Vo1eRmV8KXY8KH91YnMGPZ7w3lEQmgZO9QK6PEUkjm4Bc9YcOQrBEO
D5oshy5cvgMrIv5munQkNu3RgXgI1mA0nHDouYG5sdXdAGLb+1eFQ38OladEZoQl
ehpCog/xgy93UGOzRO6wEWgs1UCCL79GGivvnZ6cpGbdw2NOtfH7tuQCPmUVO9gE
c46Hk4D4bm80iOgXXQ9Ftc+M4ZV2kJePaog4LcIaWBKJw7zi+Q1h9xg0SzJAfDl4
A11tULhOAuNXky7k6qy/hUAOQqPQQ0f5TB62+X18g4UjS9vrA4CUv8s0OgUSHKzd
wbAON1tYD4f3NmcwYvVrSAU6WzYHN2Zh7/yR5sksv9F+h/u/Q7ELJt/2RbOQgEHd
foIL71U1o1zAu53CBiIQhbomjmpSx3Vn7HuQqUc8TOaNMP6u8DJzd6oSYRBTbVm+
B09ZF9OEYXjj4XOmTMguH57EnzX8hlvj3etP9qILHy1Vg7d3S9XacUEE2EZBL5gu
cx9q83jg8vFyXXayCc2Jl426kJ2OrO6dtTQMZHuovZciVHCj6ehuiWw9SmaS7BLS
EV4NYL0Y/8VaX0rw3cJca8gqnZUz8RMeGGmuuugRJEX4FRqQc/CHIs3pQvCwa+U3
QdB7LPz/umF70Den6KPaLNrc+R5jRdBUIvJe+a/UVDVhYuoCplGpB87qrs8ootH0
lUNregPX4/Fd18gyjBFqloeTuGDGSfRV9zOit6yoVOqcVClpYdQIEkADEctdFIRK
VY66giVG8jJr7oQ9dsfG3hEE7++pZ2zvP7rspjdm5Io43nhJ4U9EDhUJIgis4LkY
q1g9Rh+hQRwCpB503TSUot4nZ02qK9ChiNhjjYKRHdg0V3bTTqUNQ8ZcfJ10CkvT
Rh7R2xUHd1200rzyKwSNY20zc577q0CSQGOLefVBIeyXoQLa/nornWQnAzUaeHi2
2Gg7WKBKItu6ajudwnDeOLnP6b2efVJaAchpkPOwMTiEY5ahSwEgZglRqdWN5JC7
J/msqzUeTyUyevDQc1Wpgv51de31GWBu1iBm1D//BFKzfgh4emmlqlotr7aO0dXw
IUsyXN0lfESidotqm2DXByuJEJbgLy/jswZhzeS9Y39NODW0iIUg4wBH6RFH9pSQ
jita+kOAkG9PPLYm9yCzi4mGAU/V1Vye0j7JCK4i2kbxxZHuenz4/wZrWtBb8iiY
ZAskTA3ain0G20mP/Kj0JDcVfT3ajQqlsTQidp1ASWQVTOXFfk6lEtu4tu+U0tFj
I3LKJgIus1AJWs6HSaUaKUZKm6NVWBm+onXuPKOq3A8MGd5GdXohQaOIEf0LVHhf
hkD6kqohpcJ81Y6Nlt4pLzvVD1AIFlybXAiFqwjRck1E2ihxRU9GXKE1DH6UjPuj
qOazymVh+p6zo9ya9fzgHwIHUTomulejKz9BouC5u9cOGqI9LbU6OjuJjblV735T
F9jVxZReA1UXS4N1zk7TzduTbboLspLmKN1hKj3D6P6C4jkDDaOiV4fe65oj1K8f
2EcZCWwm1NqvHEWREhhOuQLQtAV9mMI5hqx2TR7pX/IJY7gOa9zEimnCMBA+30Hj
YwD+4NnEEqjlUZM5ydeoU9I8hMve0U/B9H5RTSITB5ZmkqNVkq3khPVfwD/rGliu
TrD8C2BClmmSSsdympusLQurgDnq4EM8c0IIdP6dMlyY7Xze7KYfkgPxbXFo+R6a
0YYoEGUGz/u8RBgEppQN5hMYx6olotK9nQH2ZG6elLvgf7Xf1Ce6haWqJWQMUWgn
a0y9DvoFe+WLE0LzlXFV0gdG2zXY6dK/ORho0FtvgWKPC8YrrQTTXQFeggecS5Ac
/UGAo0/I+z29/NOSCwWr0uKmgjI+9qSIE3/H9ZqDxHWskJ/7CvowqGAb05uX4zjP
atZfJYH2P02FQafWDwL0CTA8vyCPELFwSWDQJFs+JpjMoy05t4zTD1hjDY1ci+F5
XKbbiPpXS6BBGKDFwm/LHaGanyPTReRRObQcl/xQhQ8oel0W1JSOTppIWfAQ7pN4
l4rjwNAUuOS4ySulQ5tiYJgWIKXDpPwJMgWMpdYUhaRr2QKA0Os7eqa6LCcrXvZ6
aRuS2BOg7iQTPiFMh+VaZqDGqmpleleip4Ui3u+qoY6PwZnyjS2Mayj/BcZR/Ojv
tDFYoH7p3m8qgc+LpenUBaEXu1CPFYQLUkbwJTa9PL7WWxZ+uD48Bg1I9O061crn
HDHq27USjfuF49nYwx0TMAmoQJpr+QUuTAlPmIgL0MMqOY2KkVUpaFDKkTxa3Khd
z0M8UR91LGjy3hQ388C1AufrzmuzXCsu3BqiGhTyjMGLiSVXahveAo+99U701Myf
iroW74bQOM9yLcKxH1CuMBBNtGFkmv4byYGXVu9SrXDO6ATYnFZFJHXxjewIjNxw
LQeD0jq/Odzk/OPwujNli8rkKykWijcbTwzPMWD3sUxXt7C/3NQ9I/KHBizao7dL
Gi/4PG3PcReDAsLmu1d6VG8rYXKNxLluo2fJN/se/mkvkOBdzRGZVW5X3fliFfhx
vdVlbOOyq3vpbOf5qeOAoEGoCvUaP/OL2dvhwdvmHkCxIpVAtJ7Oyecv2YF2qm1M
yTmYKq0uUGpMT4+99R1xItHBVOLmDFjZftvkpgAlNHVDdKBvGM5JV6apkq11IphQ
qG+kQifKwU0zWuQFjdTNduGoOnZziqE+P4L3Cm9gGWeNHaNOvXknB8FoLUANCvMp
wqzG50hSCiHaGBh7dyk1VgQQ4qBGctrnTbq4wqd0+xlfqorWp9n9u8XTw95a5yfF
tzQG/PzpIoUuNu8d+jNbW7jD2rD688hxn5IIyCRM7gIDkvAAtHQ6ftO5wk71Dcjj
C/QVEBRWkARDH9V2dTmvCexcy7k4CMnn2+s/pt/RIHYlqcCiN7Md3+0E3iizFPkX
WIwnFE5cYNPtqwavKuoP7HdvIfGP7qHDW7oNtuDRdTZrIT6DlZkoaWTNw+wW4Bit
1yMDIlpUqpbV5V9iCdCKzWtkG55LI7FLtiNsLKcvoDMRzpa1ssR8NvQTOGmqeoYa
kFIjPywSm2S52ce9ncV4Plih8FuHOR2Bk88y1pXBRRNNhX1tlZme+p+QkQdXvT+2
YRg1tR0CEYz/vCy3pLv8+wl4YaBoYfh8a1lAyB/8+nYHfrQa4SL29KX6qVWvzxyW
6idZFA7gKJD9ZZzN//jn4rte1UfHPGUpL1zPbmlcT2BNyCMJJodDKiyaJhev6riR
WABueYWIUQQ7RO7XyeXRBxbjZtnV4xEv1AtAznEPoFQ3Mf3WjwtKh9lvFH2fXHYd
R5vlLwTRr9d3jk3mLNMWER+rcEGH8h5R8f/nH5n90j0QBLw2RtPfGTf6jtM49XmO
Z3iuf+w4Ll8/uhZTIDJbu6pi2dhDN/jG8q+dMIZXytf/jIyWS/p+s9tgVr2aZPR0
kQWrez0YRzdcxgbqN/+Yh8ISYp+NRQZO8HaizndjnpIv1EYkNR4U4uWbx/xxlEwf
piCe4ZntHbq6CLcJK8+O6aIpYvOSHlhFwbaPnPR8fFSKEYVk4YxlNcDpYuGbcRkV
hY1GJM0OQFuZyxUi8vw7brETwh0fwI6lG2KcFBEAbgCR+U+h1dZiYvYNk3/X6x3d
lzm05g6ABTJvl1wBWot0KpLJq9lOk+UIDV8YHAdIL6UCcD1fSK+XuEHf28RGTsKZ
tVtpAcnjvrxpfgs97lDljKwgQk740IFsJtQ9RlG7q2UTMP0XoL96jfL2fq+yHYHa
Remdnt3gfToKkAgVVGmErd6/VaHO1+TlQQkAcTEeLI9iUsjS8HNLP1pRoSfbGHg3
7kidid+cJ3BO/KVuzkNSBQlM7pT9DN9FLK75K3FNtgQTbPTj6JYO2gDfrk7pYhKh
yoSnft343QGYtkBZNuj7xBq8ZuLfEhCgGkJWUrYBiKu8ijgQyhdfypoC1KzTwANy
5lAaEfquH3UOCMsHqJFQLSNMD+2oeFJycwKvKqy2uHtAkRSsUcJWDwaIZniU87MB
LB7iVM2KURwiGQ0vt9Yi2YG/mSmITWGibRcdUTmgbXnvi+Ryla1IYxbou5frK0tK
/g8zgJa7EETGhgUZLCbeDCxvMe6XQDAY1JrQ/4E1d3ZTEDWghPn4aJbGoF/8Ultd
cr0CCZMGxPLvVq6aSMKgbIlgJ1kDZJh7g4j4DLMBO2OcCrSoNImO9UI2cxwzHjHr
gx2EgjXmEY6tyHVSdJqb6Ljw5OcezJAsPs+gy4oSbcec+7GFVrONiUDV0Z2Lvgh8
V0K/r1cFtlbzK7riQW8cFQxFUNzFpmHObMD87w8QTQ0mhz/uSaeLju1VpyV8OL8f
UugDwpXarVyIDRGo/XSKt+RrGRyetAl+LmHPqovevyozO7enRJU9xgUGYcd7wsqV
Su5hM/NHvAqbYXyx5fIMDlDbDFc1RapPi1IiMy0TstfCl5LZFQdaFm58awZq3YNe
NyG+X/m3YjBX0IAK5xe0aa9UrXUhqpk/zTdO577vFc4EwSXZkgxnjfJP45JRrklp
otImrASCnrIW34tn9QO9t0A9cyGD6+/S73BJcDqWNJ644IlMkYctYU6fW1InagG5
JV0/7BDA7T9UICkE4VK9oT4UDbm18RIv3jEB39jJmXN2YIKOeYe/K0GyLG/MQIg0
pfRgDz5rLGG4R1GRH1f4NpNCfrQvIwh5qPUDI6ahSp6oK79gYqTjANunFvkHj8Jj
56nuVv0cGvwVUuBsT8gEXtMlMu6dWT7+Df7I7joTViY7kVm4wdOoO7iblLeTE9q5
5duFmFq3AkwyCrfcj9rdGin6ERlDldnB1B41Fg5cm6Mk7KXVET0IZ4ioeGMKnWmZ
tt5wEoJ417ypj2VNVH8VyQg5isjw+iHzPruhDj5+lIAIv6L+CNuYeN4Bg7PwyZLO
wfuif4KpcxQkplucjy/+7F4DOz89D7k8PCNBjL6XESDc0tZky+bD6Myl1UlznZ+N
Y4GPXIWd+wJAPaoDvWQqbiFX7vfYw9V3dPDcuocT4an3uRUCeaEGa/F5jIauOVnU
FoONpAKuhIGg6ZrfuaPvMNyX3b4DOfzVZQu/A2j+WIh7Vs1VF9FPT/2YfVwiVcJ+
jwNFmNRkiUxZeh/EkfyawZdEuHMbmYsi5GefZ4dgbwnR4trZWF65vb71c+2Ho96R
JUSZZC7MPHxtctz1Xw8hrFX+uriM+My9C99MKygmRGIFp3hcViGCOhOpSEAFto52
uGPYLJAyKZKDYsijcV8JoGrMfngY/R7n8FtuDvCKT5OsUoup9guMWmTB2ZspYoNr
0mtPCR4/K+lQWv9STFRXLvUqen4Nbry4+oHmHB49Xu4IF04RzrYsc7VBLfvLdqE9
9FSw9qXiHhXtcExQRCuJx7SS2AtAX0YVWUklBGHy4F0CSiJbZDCkIGXQMHksQvn6
Bb9h+fGjv8WOdCBVeGBmWDyCL+3cLiUMjTuYFrhTRhQtTP/e20AuAS3DnrOitVNF
3/rJ2AWnsiIei/rUcjU/RpOdtVJmgt2RZa/OFo5ScYLmP4hqp3dp6eUI+s52+chI
UjvwjCjlFmHS3xJWl6cqW9ycjXKuIF7CZq2meXsxhwGQkJgcWrkQPA2kE6UjNpbB
DiMQ0flyTxz4HYfj5Q4nrQp6CY1QeFfUPjqWlCFljAixUSeNbpY8H73DJ0Or5UgM
f7afIS/5qdP+9fe4HDJv5zHT7f+5xQhmtt9SJEy+O1f5onEAZFM/H5LcRNYgV9M5
cIo957P4U10pyR90FJerVzNGtvIdAOZNGUK3WyS9HLWnHbgkh7wblqIenlaDeJwC
lgRBfV73gk8vae86ww2fL2ozQ7ewx+378vhj/B+uIYsTYoHWJyHLC5amlIHRZRYs
KQzxS3ZUwwV9I4gMk9q8uj0KuoRjEuT255oGApI1SWMe+Z4YUe6RDm+/JHvQI9cM
OWweHNv+S2VDQPv+FHI6X72y3KWRzcwMp1vjD8GroQYqs2kB9Vg1HQNYIp87wj+F
yzy8QVWpU/xySnAs7hUxNnZJqGPZPCrXxtaK+TeRG/NCTXHZj1ssOw+0imfAWvGx
zIu1v2ky+YEsvptatCkkKXH2fJYEu4LK2T9hwq00YfN8h/HNFSoX4j5Nl7c4JgRw
rf7h8wcNo4QbCJ1jLaF2BzM0Vj2B2AMZ3s5Dhevfelr23TB2u2UM3nA8J8QQJ1tm
YH2Y9/3MOLTG+leMhwUNK74qDKLHUosYWN2K86NlggkDVokkD87cVWlRs83w42bM
EHu8Riz0TbqWGnYU8zRnRnyHxBx6z5V8NrMAJVzDd/SP/DllwMqliMCB1xvkOwQR
V3ZcIuZGF2x9odrAHNkjvc9SG2EeYtpL9bnCejgvwBkEYg551yvWmlsJ3jUdoWeZ
swTEuIvHTiF4q6bB+Eb4pcQ085kOohd51pXxNtE9MmXJ4jkI6mjFA7L6c2kXa2LX
AOYN2x0t/hWUQWlrdkHmEL3ceLnVJCWYzYctz1RWp96XpFwaQTxUu2NUamFDKi7C
bIukXXGh+QP4dPBXD4AkkYv/a86CcJrSACSoOV0rFE9MhC0sbps3o6HkhT7X0m/e
t+qSF8Xxq3TioFHkDiP28kYfuU6ZhMxUzl3hR10GEDJkLG82byG2BdK613PtdDIc
nwhNX+YreOqlM6F1v8uovavPyS7tyjFMGNj7tyCqjFRnVky8dB/UusWNf79WpcaD
BETxE4z+oLTcBOSHBwykg3QPmTIOKd6sL7IB8XpqflJIyHexUwHVWEntpalvYjOo
InQOoOjfHpV6cq8igJkojRJBAgGvK67ZZ7YPW+iTwXVLZYM5CgGgxG+FhYqiDnAu
yeJWt9lsdDOXjk7cN7XyckmVOfFb2jc9zojhiagExzD0rhQN6EmRRRD2QlB7kjII
B+ZmiaAPr/iSPRdRzKDPfe4AsjtivZYEezjSOxzaD5nGp/FK8Zh4ZJ3BGSMcVuNx
GIfQZbCuQh4lbu1g8jP3Lq2JF55NbbSSpxnvJ5o6VZBCxmCKSWE3nS54m2MB/ohY
QWABnHYreXDvCKIR9qjDeqOCZZuKtrts0ZhZ6Q784wEm//wr/nI08dD7ZVQpPst1
zxt8N/ELfgz7em/nyRp8R2pEogDfcQUFntz9SK3RylN9ABg9XYHvQjiN06AhLF2I
XgwMrczlNW3el+QG+beWmFBw6YYegHaXwJ71PTGXOH8T5UJP1FzfdW9i8ROSTExz
E9uiIdTRSWtLI3Rrp1xoUy1iO8YIkwZLMD5tp+RrLLrsWve6PobVs9smTn87jF+9
9EyWAhGaZI4F0LXzSqmEnv6UbWdsNayftmEGk9QBZovIHpE73euVZVi7Q+gDAJPL
VRSBJFuTWNeqtyXZId8BHSreU3gMvQzSFhCLmYeWFHu65VaFmet0mZnjbGQsYanR
ZDSbuB54AbSVCFB4+6WcuK/wkxquEPHiJRmCNYpoGqeDp9fFxVomVcR0N6LqduJq
r/0mddsKkzkSjxsFt+s4x7aD/Oy5BYw+4U0OM5DYgMvkajj5ZtVqW3bj2lkS/NVl
L7iqbojzpPtqwf1XvrCv3tMOsvywSMhhJuO5CNoUWCSbreUuT1FbJtcKw+eUqGZG
hVoIDI8QgQapiitDrCmjNwG/RIcqXsJti/zhaLYUUzuQHLSDn+BQd9StDffrGCxk
DRZl+nFVoNUVv1sQcTQzPWC8qyq/Y9WoelPOjnLkrNK6UVDuGKM8epyajsZbBHtd
sNtBkVGCjuetqtUECj80d7ifcuSxw33IXuXZDTQ1Lg4GJtew91SwCh9lXEuRLptC
TTOdLC/jRvSMpFxWW+FZOjQwTpBwBuIFpwcPLJKtzSv8aIeHt63OrHZwwEdDJmyJ
EeaPoaY1tEjDfTvvJyEm6AVaHapPSRf3YTB46IL/lM/dC8TWDR6AAwY58FWQZpTA
zACIEkIOYBoiaJTUfSmuaV+KJLAzniX/e1kZy7HuFI5opFTP2bM3S1RpbawKLT7D
mw83sgYTR0EgqvEtOykWlYNJETcNuCFDfQWDl0UjeX2ehFFHlgptCrF22LELjP7n
sdypHKdSZiH0f7tK20G/cVdfof03618udIzmUDZUar2olcMcQng+ED+57vEWeUey
zk9UgbCoDXszWEGSIwJuXMlePaFsnk8m41/l7pUq78rWj4g1r0NRz17bUka/QgrE
HzOANwXYPNIgzDS7rDgcRHEj97YHPnU7uCRbfbz7jYYfUJeq3YOLBhr3oerdiLtz
VHzmhkvnTDt06k2FjTXv14VC/WCh5kNdQwxBSg7y2DJCl/EUvX4YSKbl0HEEJoma
wuqPCVW91z//cBNPzpH1xbRrc5Ti09fJV/k+RaeCRBKSi0ivu+QE3Bokns151ljR
VhwsqfOohAoOV8fTFZzVv31BBF4sdqbJvXCdsPm7eUmVA2N3vNN7UYSaLQYMKVf2
WETi+pey715Q1TIIN2QrS2hQlBgdmLqc5B7wm4CrxgKHJPRfInbq63Nnyu7Ua8v7
f8L9PZOUJN4Y7oN6lKIAI+z9YbPjSaSPcUBiXWM9FNGLDqpYJ98on/wY7KgpPjwT
+qjq5A776eiwQMF7oVPcfZCgc3RgL5Eau07g8UcJCc+lfmfDTCYdz3pzavb5EtUp
r5yZBNYFspc3JQBb1qhGExt7SBolf6l2ooA4bMKc7taT8UgcqlttR32Qb+KwZfVI
IMj8X5BAfZL4TSlUg1AVHncG6StUwdYfJJTQU5zHWXVecTjNXkupBwRTxn8N7/je
uX676faKXt5pD6KN2A9F/Rojg4+IF8CLlKT/V36JZkk7mKYakGS+FnZsPdQsGTwx
+6snGUBt8Do78ElZ48xsAxeDvF5xZK9ZXKJrtn5hlmzqq6PbD2UrVNLCeU9PbvqW
MAVR2CTQ4fAZB+8/L/rbnaeYIpgd+EWT2MCL1LotnHV9PsgzNG3caAuPJBLU0X7R
6cio+F3v7x02a8lF4HyGwZT3NrVqiF8b86DZY8TQ8HVCp72dAo6Cjg/uuJSqtnKy
6wnwDEKSEtNQP4apkGxAkDSfiBNen2aoXjZeBSpLsSl1OiTuMA5Hd/sJ6CDfoDFK
EVgA5F/cSyYN4B4UN4piMvKD/8YepSxbxgsqyZmxQo64wJs8xR/Udutq59N4XOT3
Eow9GFXgDB1vfxjz3XpeE7qfjTzhRef3NSNgS6XnTRz8u2/6J7nCZE2haxGnfIX6
/Qdqo6DcPoZ+20hKSXLroxVZAUUe8K2uIy07tMKNwnpEAUK+VKcQwZzsflTOgOPR
SKJLLhf+WRW5Vdglo/vU8BDVoUgP46zyGrEYBC/CLKb7ZebEpbYwOWXiSIXWlS8j
m6K/l5IEINTqegcAfsAF6tlU5NTZVOk52WSd4E9DFueDHuYiCwlmF7iKVPbZfjr8
1+Og4yPX423oRh6nOinSVoKme8pQ4BxIPcv8Zqfcea2TceE8+zOjEINrI0aPvOAg
i8V4njVd/w7kucL1iImqYWAob9RVJKrjhKQrPysoD32SYfBcskf9n+c6HB9VXpYN
zTuHV7g+fwTOjDbBylg6ntuPFGTvBLrcuQSLewC3cxUGj+W8glvJjWXgysprB26p
S+kFZ56rfWV1frDZ3ZNe1jkyMAnIP+MHu75YqhcGv3/875cXl8/VpdLMEIbMe97e
gKAKVgEOs1bwHNFub5+PWUnVlJMJRIEY6rKqk4DBDt22069EC40A8cUD4+CQ6gp4
bNJ0SSVxC6iZzrSoMu+lUrKhqCT6OPctdNvsieX715ywBNOhluEg8sxqPHj+zTel
fZNUn9+tYVIKsetVx8R+Kw8rRn4o5r79YJOCfDILEbDaJQGA5gevw43E6ABRY7Oz
9w7Wf1eYv+kX4IHYLyYiJudQ7F3MRSRrE+/BqodIdnDNrOe7fYtPBVpVqfFp4K5g
f0ZDuGyGqcxf3R/LCxL38LK3iUcDJpelZmihkFuFmK1LvWOJu55EWntHjUlp4SLv
TVVeCf9pH/GnGNRomFS6+6QTMI3/2gy1RoXORxg53diS/uwNf4inVnMnYlYH/K7A
Te4XWdyFaPQ3MwxNK5NDAFn7xORKoao+0JXK3/Uwc5jDoLxRE2tStQTxGOLVKWsa
fpWusVQzwjQZ8zIR2TKYg1Zt8Uj2vCEbCuJgomN1NWYIObl00CNiRLVl/QtU8msV
VUAmhwwPLz1fg3iZdXdu4Iahr111/uEpju6BTizfPmBbSa119H1AuU5seehM7Y9X
/3/8/cJ8Qlk/o//bcc5XlA/6a4Mi1UWbqBKjEKFLFgue2E0G3fteJcL6/jyxhyt/
cKpK752GiXHx4F54FU1uRA8PSJCFWa63PvDToQ48TXMmfunj0cSWms70t7L5mPBC
K47XfIonDAsGs0jVvekkHPlV0o2jZ1SkiVydbhqneGgRax8conO75Pfc4IrZ28tJ
c2++IzDN7nAvxOZ++ltPM3ZEnSvd9AkY+0NSdW7QDr1YGuFGYwJEjRnGHSvtX7ld
wZ/pCBxRuZSOAKZcYyNMW9FeVzLVxvgX86gzVPFa9z2iGpqOm+29Y2LyIJ58/6TW
UsDANAxrBXpB24CTLEIBrb9Ie2SenT4N2GTGLvofOdyY6/rha3fqGJ0hqbDQYUzp
ltRm267aTSkvluOMMRSbDrVTMmkA/1nHXvUywUDLU9mezhSgTU6IfiLDJlvPK7RX
JpWjhdWip8+3A42K0gWe/Q9yU3jnam9IxvwyXli6AYMsPK1L9U9x11Lz8b1cArg5
nkMIQX1+t/sJsHi8vPDUrQh7lAR4dObvg2d/a14IkrxG0CxuGlagnGBhdRJxTcup
vbjVqXLyoyL8QCpdRcUkOHKY85/1oBl/TNazl3gFTx/icFKicO/oZV95bjg6OFVL
Q3oBr3gK9m+EAL7a+poDsp0+djcNqhGwo3K81rayP+ah/wuTgnMZXOcr9FQ9FR5P
r8RAXmLE9kszhaNdJsvVHFLL9CZK1JUdci7HQzuAmw7QEwJpYpCjQmVBwk4uSfEt
lJNa4egpbVWyWpCgZ6nbvu68PrxJYyXRXqGfx3bvnxsXJZMy/f3NG/WdNzUpPlkG
ABAPI7/8mtoYA4GCsNac/JWV1WYztQgFBZOQtUPUU87d7fwtSgxDNAW791ErACJw
Cs15XAR6yPSsCEfv21nZ+BVjAFq6kwcZHr+ctXOuTkuUP0FhvaVJrS2mdN62aRJ+
M/79Cbmmpoiqk1MEAEd3BMm1fTOGuYUtShc+vrGXBlJm2Qia82sNk/uDKkS8qx9U
iE1VklwGavLLtGQwQVLWTmqDwVHTc1dzqMwBQy3jUbkvaRwarqb3BXTI5gS9kNaJ
M9rJMdxBU4tJk8ASYguGWhasooosDE3W01d9VXxm/g2fM7ZHNTLMyioRXVDxff9+
4owgfN5Fx9JiXaYVaq4MkrIyFtUbAokCedOfiYiVkClAm3jX9FNJKNuFQxQGVuuT
CNtqMobLMgulXqK6uY1Be7vd+S4Lv+dhxLKSMLhdVnLYW9PrvDj7UiNzDpCwSay/
cYFQeClcOU4y+4WSTlyJq4ok3GoSFiwI6jPntEikXj1iST2ScpuDkh85lAtdp/vb
kWKba/vQF75UypgS7DMDiovUV2gSvy1vRkfmQHiOQvoVh/2GiKIwbzve8GcXUjY9
F8VF68ms+Xh8K5PjqtxIRYBV5Sx/OWaKGiDM9lTEvF6looHLZ+QhsgtPaqOMM2xm
veZdCY4yB0KjCEBdC2n2e+sCI/Om9F+vUXDdyU4Ufb1YkIBUDjshE9rQcy2tIdSs
ti8tPqV9uHXNmN69j3RfCv8WBImTc6+Qnlx9LqvK3/AwgCKLTbI5zWykaefOgXm5
ZDqEeE36CQoyw8aHzb3E94raOG4Mbv8UAaykJ8haZrJvSs5gU4Ns7soSWKoHW1k3
12FHI3XU0Tqx3QMthsn8r3cuEP8irXATB/4+++nu518bM6Yp+4v0LZ3QA0kTEML0
rVWqnpKtjXl1wfcJ5QLLftWEA0gugD1B5yIXm4FhgHuXN92dgmXYtXZPa6OTz75D
cVDU4+iaT8gZNWNcEMt18cpcxivs+WffHMSlcJYq0Ig6pnCNWkJRLUIA7xn3M+rC
GOwhGFSN5hQ76a+n643anqDbvzL3audovQSR1ZEoKBPq7N0pRCZekDanPlfttI5m
BFjrlPuhbOs2gt+i+no/1y21tdpUf6HCN+NOeWPb70G6jBtF5OPGTjG78hQDweo0
EtlzxpjOGkUJkmhc4WTP4x6Yeg6xcwsoj/xuUHiFmQFtsE4O9MGh9RMDGKkEHtVA
MdfvKjM41Nnqu3sDCHfRu84WJY0j8nC1RilBFg9xbmAcq9iMSgajjbZ5eiGzg0SH
I7PmKY/maj3koud9J1UFNAKjPnIqgXe0BIsn9gnQbBNeC6bfHBedM5+qnbcSnU9E
2pBX9wO8qsVvPHxJygt965KRY7jO/PCLD9DPYakA0/qyy9tCM7n046sMAd0tn9Iz
hrBqyEs992SDU7K046C2sboChcG0yzWsm3npQ23ZOC0pOn87xOYvbDP3SU14Cu3G
Q7MYGaNgHbFlkBXfHees+tQoHoKA9djLntAX2NhjNqNaEfLECS6wyGezvaBzGaHr
7Hve5eOaCiXYzrVJXH6gagWqjxitdXn0NX15+z3MquT+/GPD0lXE1G7ghLrRQ3NG
njrdw7S2sUNOPehFLf4PY4/3xMbm7aOCwlkB2Pajib5RW8vDPnPkwerGLchwC+gO
ja2tFkQs/FsRmBGWBakOeC+K3Udz2HRk9HIUUO2EgQCKiXHHlpXTi+G+Z5tJK2Xj
U4NGcc9nx5UfqY1PbZ4xN2glvKgsR3ug++HJ5vHrqnMJGSjEojjhikcPM3ZQeh9a
Ph0ktIARZBZgJNcQaqJ9CLAgL6A1WuWCQpAyXM4s+R6UwgarXYlefUJ1LYRHePom
ikFi1tT6guep4ehObIZfz37LYD2TS3Vd3P9C1vMQZQwrObWfFWSVFSkAlbfmsc/G
6vV+Q20D3Su9qaAPl7FpQFH4zdVErH2a6qiGUkzrjaekCnAM1bVWvB64Q1a8WxlF
a8uzGhheLmexJwla6nL2ZmZ7njjFQqF4vtTUNN34+NiTIAURIwMxAVLVkcu+9+CU
hyORspJX2pU+Mnne/xQqliryn+4v/o0hMeHd4tVgrpTpShJarDiL2aBbj7XmJ/L6
/eNmsrw2uWv1amc1YjLiH3PDozze5kSglH4W8N227aSFzT6IwO/mvi9m+GMRfSwV
YZq/hbwiAsxroRC8coHKNtH0V7YGhOmVtYiT3XdSh7rHzb3yFuwUth3UqwDMj0Wl
Pi2LxHxY+4sNwv5KnYU4f9iKfWxvoV7SYoavlXnCyZx5BLAZlxh8ZgFTVaBNrkjQ
pv9y7sAGyuTTp8SjoWAcEjn3RLqZiCqtA0Y1aCbDZhoBCi+pun3fHH9Hwe2rqAja
sQVboCj6zFxfPWRWT+ntvH4m/k+uw7uYmBIA8HCcxDF5XZGZDEfHS4kWTTBhnY56
pv/RFFw86ibxDf8f4qFE0vSa4q7LCKIOiiJ6OhVOG+VjiHWHfQN6jDGgwY75IvGf
1JNG3wgz1jafo5SiOqV+iev9GhFLg7+Tn9n4O/Shb3Ukvkjz5AvDEcAUf8OlGm3I
uJmoDJQBzrypxsbldNlxA9vZklwmhOEinOiBeA6EVIxtFObHg9apwA6dvvp57PXa
wstU0kiV1Av4jtMg5IG/4k0mITKlKwP+nklMXqCjF/yNaY8xof0y13EpVRZbLo3K
yBgqkFWrVRS0PjxoYU4BcFFr5qX8umiv7pZvk2AaRe/I60KrVQik7JEaW2KOVamm
Nql2edZst4J5HlN7aK/LOMTn9A6Avbd1+IFV0d4j33Pn6Ta8Mb+W3E/nucIScBCn
6LaIKe0vmQh0Wpyr3LPTwnvOZh03xkmXdFTf7hPkpM4jlF6ze7T1mg9WZ8TY2BEe
Ut9N/lXE4jOuZfagdIJCe7LPVcH+2c7D4akMDdeHZwWNwo3xhJzK/Rj2pyItO9NG
+XtlZK23p3+Y0b8mMMSLJJcFWwCbjggj1jT2eg3uzdjLEXgGM6YGYtQZILcff+pa
BIygxtBFlVxX02pxiCEOOLjYaNtzZ+KJHsjDOnb945g/j2AkwFFkVRceEMv3OAWO
Gf9OS51GhyI9nF0hPNvjUJ6EudV3ROd3e1qTbIPdtyKWvTEgSEy5drffsCKQYtS0
Gl0atkhlBDV5OMKuhADV+kYkyXQaQ0njlgadg4ozPigYG5AD6vIiVcRfB+F/SKb+
ZIjOlo4GLcdT9vwpmpP0jmBYYBKckUzVfN7ZQVw5HgFv1nEQZ4QswVR2JJ7vdRKE
Z6rmS649lY/kFKbg0K3j/YlieGtNxgI+wavNrL8iUJpoIBmSR59w2J9uh/yTGLiK
xuvxcoUi7nL1NkiziAFwEn6YM3/BGcK5d+7ChpcHdk1/G3K4Jlywqz5zFSRTPhOl
44GBGN2oHsyJYVPjzudVwmH0jls3N9rwUvr4mL0k7tNIAxRlgipeXnUf/BnBBux0
En8b8rdaNXttneBERQ437+RIS2kB/uru2T4GewJmJl1d0I9y53WpTxyJQF2p4Nhi
6qGPHfmdkS94edkYhwWFwmZKig7mZe3/ubTIG0FQiKhvZn5fin3Jb59RQm/hMoLZ
nEeCUVcvdZRh4enFSkPyHiVxBUTGJHP/hp/Ha9yGAJqze812Xp1IfuucZGukzhTY
fvPqpMkMCwV0b+6mrV8CdKyPVnNb9VDXtVqOzLshaMPUgHS+ppKjnyzS55/qY4pw
weWqhiWzODUuKOt06UDqHNwEw+nf/+E4zmL2XFr5h/io1CD4s/ll73Rzbht/jSh9
zJDy+8tItuWuHMx8S01KRPh6wRXMn9Q2HY8kD6dUUNN/zn08TE+Usa9h+F3orA4K
93Ty8sbl3XSUGlkg3VTvtixmMjg4aI36jbEmwJRYsXs/9J1dvwv0OY9zo0F1aVQY
9SfF/NIpUBw7+xgb0FbJEnGJwKf1EccnSazvXM4Ij1whIRxGZSvNQp1jtQ5YAern
7mWUz2L9RfEQ20YlYFeGsLIjYtnGQ6oZnB4JDwGq0xqRRqMTMo4zk1dOD30twOy5
1euaLhTcPQdvRafPupUe1Etof5JUNw5KVGidCjBCLI4nW7pFBjHqtc07XO3CTrR7
/DikUOCxiAulMZXvJmGkx6C7qvGpNoD4h25hv/zqFDtW2IQhaPqwy5SNbEnmqZgg
zaQgfnrNwQ+zbnsq3sc8OB9GY1nuPdcd1EVtzKsx5ttJ57EbkYiby3u5Q5pjTRas
t/swLnq/TgKgAavV3C3Ol/5bAGA5gfOHa8ZF0ptYEsCE6bf9ycAvELtforrSVtUC
pNBuIu5any1nNRadRaKT0FA4ln4p7Lb5xppa+TZ6rNz66rEdKhNdg9+HGllAsSuY
ZgMpBFor+pbJQ8dXRbQ7qYPmWi9Uiubig4GoxUq3+zclwZ/pmVneHCtd+pEQwn7h
8dVe+mFrMWacQXgOriniPQw7QSpxWB/nPmgwT+eyDSQOANBvKARO068DH98A67sd
pTRydJ+6Nk4SD4Rdc9ivrBh0WNSXjUhH/hU+SqJcBjJD/oV5iEW6eb344iXrRc0S
FefeUiRe0jPT+zfefhu0ScyXfDbDdxw7uxXgrIGCWd7vJZIvxvAvF/jw4Ilfeibu
X678kb1o4tzSdnyA+1ELLPxydN2yKJsKxijzD1Z5ceiTQXkE9GkR54X5p+gzeKO0
Xp3e1D5cLdoIop2FQrVMj+8MzaFT58qWQ0BhPSztroJTbenDURtNzbhpWTFQnvIR
Erl+RKjNhP5Q50DVluuI0m0quGWie6KEUgXTPSPDXg6CJamuRhGVnXQA8G/kDimx
ChaYi3NCDnF045OUTgU2BaqMmCoqXHYhlF3Zmkgm7NgiLvL/jdwMQMmVgORyuN4x
itPs9bpeIhxUholQNE/vtDATFezPLrM83u67qdrE+izamsZLOerBzt6NjPUxOYWV
KBi/H0KxUboL604UeQ8IUi3xnNamqX/WDJcs6FO84ucSEDSH3il6AMGk/oLG495U
0qLV8dydLq/VrUuv/90iU5/xH0FhdxsGxlDxYJPxdQWYVBGJqRzgXJ8h2hMbBAJc
JHYhVeCdMuympHn/qh2A/KgAusjhkSw5F+5w/suSVGKJh9TJKdToUlWLVv7exwc3
owhfc5kUrDAz3gL4I21ZS5Gmw8lq47dUzvljnbR3v4iBvsBhKSOnzzU3lnie+LDh
zTLUzJhAFa9MkyA7MfO7GYL4k7BnzWNknP6O97MFbqaOTwmAlv58RatMoZIe2+C9
8ZkdD1uOOGj7fte7jEcNSC4TJTdlJ0WfILMJyYRUhwqASJPtOSxgo7d6ubMtUfZF
B75n8Rh6KHfZKdnLeqyvgLSB6EaFnOKLcZAKNZ3HYnw92KReB2LZ90G22ffq6KEt
wlzEJlaVLRXVzcTsLALkFaNPkJ5iW1nZzCk2gIyE0lmMhBZMvjcTZ5o8K7m7q8EH
opeOB1Bao3XCFXQkf8HTqBsNXn7WfD6ql5a4toIbtC7eltsWyJCpjGBJmYM8Zv51
zBnsLi6Uc7QyUpshZa1GA97Z7LgCB7jlt2i1tQ61rzzCzBll5Bm0qhGFDde0Y9hP
d2uk6qV5DHWkvZ3RCJ59QqU9Rddjdy2dfRXaml0CbN/jioujJ5V/E1mcni46UrPs
x+dyr3cQ+aQpIqBkx+LaTGh6oGhHzitB4rym/8uiPdAf8I6ZURQVCWNMC+jpRwf+
UTv8WyKeTWzWt/LFVr/oKdkGY+I4JCS5RhR6ZDJ5GXqlJzOlvhRikrCCaneVCKvx
hUlAC7DQcTL7eRh7G41/YWwwzquxTFQI1sMpKG2FVGF4RltYWDCVlVH3qfP4AbMS
fB4TNddV9MOUAgtrbGAKI3NrrG8tYzSX7lCNQOWtMUdcF+3wwpaw3HuY0vAQtKfD
+saUmeg/Rylyi4iEeMHy0XuoB0wZTjao8Lu97/hD+tNZO3g+uANH6E1qbgdT4/TL
egFoYvO/jzaODpcfL5jsD18P597vcy94XSBCaeACJQOlkWThZFPKQU2Qd6SPNmAe
fmC9lABSxqHQeW7LizArLS96YshkRXVvhUY6lf+vpx1o7A9arb1pY1wyG1meMVdO
lfWa4YP0552YH3NBJY6q1n+74/7jTpCv369axnHrSBEyRZKHzIUCyZ6AbhR7MTWm
lLXWI627gj22ju1H/lRY91ey1f7tmhJ9AOQb5pNrBMJ9i4kaGkptseQ+ji224g7h
XBXuJubFYhBQ58kjP3oWTpJCrUgj2jaUaNy9TFLYV9DV2MqD8KWmL09FuSNUEFnE
5ApnxKFEOUDUDSBHEGXwvgvwUjNuLSfqlhlPzJpfWO3dG/CwHXpU/S6UroTrMjwc
ZRzD5dHQFYriJgjhvy4z4Lr2Uxs4XrA614wlQnz8VcioVzSlYJ5GveRGehdQ/U5D
cmQKf6QTAvog0ZvWocuEceiwkT8BKOeltZT2JkMxt2DIQMFd0hq+5c364sQj2fsX
sKneMFo67mXh7pxZ7BR3Wnz3o1tpToYLVdY3LkNCrJHzQyJLVA/0UbQMotQ9fgPe
EqFF6lH6i1C3iV2Td2C/iya9nEG7y3sKFluf2cUUYKez0SKOU7MQisKWulyMbA1h
4VKRJ/gs/lzWr3CpD3KHG6zWi+m3vOBneOJ17aMsRlFRJUrt4YmDqueb4qA730FI
Lg+WuymfxZnNH6ixRiTUFmida0ewBPk94QmOOJrE5ne9CAVxEcODbX+/Aw7LOJFw
53NgWI6Uj/jybAq8tNKuMixTA2kJPNxtXTX5eMjDOt7U18vWcvjjNDghUhGOt3j+
FS2D9IJ7tA462XKOAFjsFGAt1stTAzmvVGYSzC1ZRd40tBOLGjgyjd/8elr3+38H
6/oeQurR6fCJPXrMPvkUidtfNfbLOb5xixO+s6VNyS+kxvBRlIQhRLSKCjQ9D1yz
tftGWzqNkJpB+3SrIHyLQ8u47IZcbdnu1GD7Oi8laFsAX/JnLVQlPyAkl0JbVQCU
3f0lX3+KJKH60F2MHM6daqHZR9stO1SP9N7t6KE5QCrPxPmL+MbOLoCvNpXqev0u
f9qes3auBPVnxfFuL3NL3yY7uFRoZfJv4+lcruwmpwX5v8TNrHhoNOqLPFEA9ztA
3amw57Qil/ss/RoPuLYn4Py/ByyCrgo4UVwrofOYVGe7zVhrYb1q7eA8MF6haMoL
sqc99sKZ7w0GU1mjfYcEkOiLoZXDDEpaKoFxkXk+8NNp1d2Ma164bCbJI2ly2cQZ
DlZNz+0XFdCVbK8WVEt/Voag3eNUAOuiIzEaU+HCwP5HlQRAyQB5+zsWx45RRXwQ
ysY+qwsC3Ll5OAEymIe5kgw6SocHbEwxWbutw1xpWmwzLz9VZs5Ttm6JLGWPKmzy
Y6fwVzYKq9sCzZfR6edHb0OWYsjIkwgRXVeWbhaK/9EOqKQJw1E30oO0O7PL0ZOs
l90lRLUJw1uxkYN6+Q+gcSka/dD4mdtrdMHGJQldICE94Y8wAMpZwIjgx+fkogpj
DcWP28qWSKrl9qBjEBeu9eQG8tUKtNe2guUEyBv8NgLcj/VulXg2x7aaB8ncf9HM
QQZiuYU2nk8APweXImqN7tiUcLYDMc4FkEaJSq/izU6h9IIOYAbj6VdIjEPiSo9g
4uSV8N3uTq7CR+FjNkOeSPSCZR7iQp59h+tpqMNu82iytRdR1Lq2JCuGwCS9roXR
5KURyYNxZFgTmur3ZbdS/Kb5QTY4uWN66UT2CjtJfuuuzkwNsXc660vpFzKQgLp2
JAF1gC30kqfNow3Ks6AUoiXOsNiXg+gB/m2a2ekZgTgb+i2yIK4Ta1C4t1zM5v5V
dlAOdAXHokqcQx2jqweXsl/ZxaMwM2Zpw7cL6fNJfvNXl0o/hvoLgGa5CnWLNLWH
baDmrM3S733qdTTnIZ/4B4F0FQxLGajvXXjpRVuSO4xHY81Z3DbgFBkLfyTD3Fep
uXh3eM+ZsF33l0tjwgIrL1EYHs/87aiTo4NL/UYqUAoBk7EeWtM3lVoZs+mqdrPy
pYTwdOHKx/JKhJ6RSQovYLCMLF0b9eCPKsbraR9vboELmDy7jSQaUvOO1fP5iLCK
/RmU+AFjq7b0A97GZ1jmWhsdbeQAqQ54DUMu0eq45pYRUJGf6fuxInbWWiNRo9kG
fofNj3r/0VKbRVh0EXNKZDB+9IeSzS4kqGXmOl6IrFwcDrjZ4MQAy8VKm6xyctrN
0YUuE91oOut8YukY4VhDPxkdqPBBSGXmLo+wY20fijlCgOxWNVdUH2uxLayj61G4
Ll5iJFMX083OZlBIEKDtA5h3AssDF1Qlb3BUHETwB+UccmyWJWHk1Pes8i8QMEeR
kn2EczLVIe9jBdVRvELVfKXVOtJIigiXxUV0rDVEM1Y8/QEHFzAOtw+ZJF5a/+c/
9LK7AwW1Xa/X0apHTS6EQ7N9ERFPgP+MBj5caDBnJTrHEnzVTHX2s/DTE7xta6Da
ZYreZvh/bPn7Jm8v2VjOjyW2BMqPBB6v8Yp7izMXJLAsRaKr4nW286RvRJGdrSTZ
8FLbeqb9ISJnX4cSIoQ/i2tQfVrStXB2F+vVO2a+AjVcGn/R7Fi1B+CgcVLT06nL
COIRK7pCF7QMhPETmojaIln0jNbWPPrzv0cI4aUtEUlM9JuDphocIG0HpdfXG1qL
o6zCDNzuKELdzIpp4EJtiwaR8Vs1TE518oMdNIN+KTX+arZZ/7q8H7P4V88EgfQF
oDsPWO16j2lnu8EzOQxwm12W5TgCxdoGEJ0e1sOAot4M51RhcRs6Srm7pL3V8Zql
i133ithApIbQ9l7/8vrzwKOsm+58JfoMWB6mJzbYBY20SOLW3ohTjvWOhHTkzvmF
fy9frUtOAt3ndOHYNBlH1gv+h8HSXAaloCJW3D+r88eXpeAhMGE7uaq2vhh4ZIeA
0i81VZqcvoWHQC8MdyORAiXN0S6SI6WUmcf7QeiHYaXfWZ5u2akDeOV5rVslZ7N2
FgejWpNbwBNNe9V61ij2XwN4BckwmGUA36Iod43CFY4VqQ1RL+6np3ljT7EJymSa
3laz2e1IkATVQl2Ski3Mox4T1SvQnFGtFMu4XvQOW52ksApwWZ1zF3ttmmXZOyKp
6C75lxhkgejBlruoaf8jNY7Hs7ZCgulwtaxoF2mvyNajXNGdC1hgHuhjuaA/Y1Wj
BvbSvhu0HpSHN4IjZF6AtA5n7dSsTdvQBNEu/FjTQoGWDhixqpQgLd6TyunCCb8/
7+rHVldiNBKfhkWnXUZW8nDDUTnqXGXyRBT2VHoS5p7LrlhXsjx87TqZN8nigETq
1KHpmoByy4n/dmM3s6y4wY8jvapHByOqso5yzT1Fk0bPYqo5HrQbRU2cfPRoCwS4
0ddQor7AfD3SSDG9v/GpmgNDqbFrjlIo8bBN/ifHuOLlDXVnFUlaGyJrbxUAhht8
s+v4PyGBEeVEZDYhZjisbd1P+Vnvu0mDCND8pQed2S/I7Tzz5U3o95ye8G69CVSA
WpvO6B7iHdAlPhu3kD5rWJH2V9v1BYpmXuho7DKHNvHtr/lqWV4FETSy9E+OAJfh
hzIhFA+IYrPs8ao56xNI2gnkY6oU3ItjPNcrDgDWzwkEKy58X3BqorUdC4ZCDiyK
n0BqPMhXRbDVvewT7EtD7jwtZt3qVlKqw1BJquxOaSt5ionuW8n4sjEk8duKRoAX
6CJkS2s8mlgG9JYGWrV1lo2a7pwnnaZ5DKD7yRIRmiNgqNhmhjqT0brtLo88MMDX
RIQKQvjecaGYhjbZ6LWeEfFH593S4tYmkgAK8/ZAEYldE2xW26t+ryRPrxYpaknq
blooCr/EMfcCIAmav57iOUmfh3gNscgwa9krHUYV1ZiqY/p3JwZTmOBSdlj7J30M
oL9mZbgb1kweW+ppz+9dLGJl4BhShQLNXgG0MG4BW06znNJ1UzKr3phKrRrZ85+E
AngaBhxFlBrE3oZnz/G0UBwRfMAaIpNo9KaZk9w2i5E+ABIkDt/6e7AOCTmHiDu3
RoQm5z8xOrXMNpQWEgNfUQ==
`pragma protect end_protected
