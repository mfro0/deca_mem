// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:50 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lD879SVBWIm+cxwyaUzOVplax70l4zpypsSqrnaGrZKW4EG9glKLfv+vYGV8B/gc
d298d50Vyz1H9QINtyMLRcTJmdDwd8En88VVRzw9TvKY8hCKma6fdXtME9Y7Xf8a
m2dmDdlQYmNhEOdzMJJki+fRSVAlQ+tUfLsfQozdFq8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19408)
T/miA9whCeKQ0CkA+xkHIXlqcwwlsyE/LOqNuY8Zk/F2BQkpiJeOVUbm+yygC1ws
uNoeCsrIHnrNj9f2UfEaHxHhNbayHVlKidIkAUvXzlVv/ezpAqL2usB4k3gmrp2V
lZh2jyeE+dmU3msAT23IlZipAHFPSv0/1PtexO632t9HEYrtz7ztbBrUIFRS5zqv
PY88sliXo//7ZMNnRJbCbZZxc0F6L8kVZ+b5XnwWsr3jLq+n+ZZ2ClTcjg/5uLHX
xkCyXI/+wlT0kYQznhQBe2UYuxTAoRUotcoNc+O2slrhgUzD7QyuxSh5vJpPHaTa
PPD5RFdnRYJLmiqjG8BuzO6jPjzp5BDJwC5n6C4dGjVBaB2puV/g85AUqt0JzwFe
mpbx64/uVfixi63x4sTQjgKQaqNqURbPDO46GQdvbFBuPLL425kctbMcXP5PCFBW
7BD4mJTAcXNw5/eqKqgiWtgHFfZf62OK+oNpRx0s4mWpctuaFkl3fDej6DknBehF
QCXwcc4TjwjIiWDK8F8WtTyx+AuaRvxldC8OIToVIMkz74DXhNig+0czkRp1mZQr
kQ1JZNtV7jcK/ZT6nOYRLK+yfiSBUkK4rV40N/8IITJQPdHYBEp/gLaIzJgzcERz
ylQOANlBuNZ8wz7f9tz1Zj2Uw6RR4bqhgq+Jr78iI3J7/oyvrnPVV3UcCaGcVRKr
acgt881Ff2n7J71lZKm8NMyryDydW3AcayfZcK2B+tuQTSy4gF7FBeKAhh/PxNz+
VtI+qhhYoLt5sszQ4Q1GZG65KQfxKyc6fsLIciq1ScPtJYRDhzD/KnlBwt1Hvsxw
sjR3/900vNLjBH1+uhb2CqTuoJxzJA2Rr7s+xJ8B4ZtRz44a+jS0ekH58VeMts0m
rVqF8TRqzPiSIwuyARUGbnq/SvRQDMH8UaKf4M5f1+eU3yPC1sDSO1+Hz0fYqfg4
RuJB64x1NHZ1gJngFrhVQ1UzAH6dXgw+FD+8Vlnk7jQx6uGL+NP5xrKWxbkZJorF
dl9QStLp1x5TfIrLi3/cxilhhSt3RXSKAVIjslEOAgeYpksSJTTuR9o6YAQIctsz
Mwdqp7GpS+qJ2fFGX9I1A9SFbnVo6nuft8Wm3Uz22D5MzgiYZ0cvC89tS0OuUh2j
GWfgJJW3iHvJ78+WXr8fAhbn60bstFxJ2QXN3p3zM5+ANMilgun4lpyIvoTtg/Yj
H6VSNUBfGl2PDPd/f345v61VULuHDSCwyaQYNWKp0EokOwAe2htH2uyQu7smcO3O
POCO/9ymZcBmomDJ+vDqgyLP+GQSv/lwU+fTW5CYoVieZX3CTuG2VlHSswxx7VwP
WwYI/fXN8RktOugiT7uKbMlr/UBHPornbsUvj1bJtKxuWTlt/4RjXz4dyG0WtjrM
NVuwcr5CFe9gG+tDaNP41eFtjjx7gMKbxh2C4ZYwQFKrpPOLONjZvgHnm6RMzUKo
PZ3iCq6zhmI5yIm3WK3NmytJ39cRqKxB7DLmE0VKQ87M/W0uLeyl0Lf+OKBrzAMO
jG/GJVErcYSi8yvq+scTZPc8nMl2xxGwvVgZxGQzw32hz6ohahhre4XSu2bO6R/s
3euo2T5RAB1kC83YCx95csCBJGvHZZ/WdEaOZ8KYL/trGysQsCPMMSoipw8wHIcL
JwBKqYiOU4hS645I3LmtHhx8M4axj9vRjxhsdX04r+3YG/9ON4gQeuslxjww7rgr
rHz3pABld5l05qQkBXqoeh4/5AkUqUc3z+ZMCt3WD2ftuLW803magT3b6La6Md7G
2ktOpKHg71vO7x/BcJ984NcCJ+vuUG9QXL+7qDHaXfi8e3qfDlEdwhTQqqBcrt1f
ZLumB2SC7p35vZwOj4dTbFAcfnLEd1eI+57NV1ZEx/evNUwF/wlKB2wLM2MzgrND
kQuilSVKtSFufEQIbE8MBHzj724BwTDrzHYZpn/KtDjg3PczaftAvXbeDlUAZgux
/N3uwhl+NTiKbKbV1PfDXdOYuX44MjzAk1FxMbuooK1gVlzW3IE5uF/cEKvdzHDU
Mj7h+1Xx05JkKL4VlcOn+ojqz9NQBiI8ywyCDDwp6YfOmYHJRX1vfO/UlVbRqyzZ
s3kTlbVlkg3aEYZSLj+iLuGluNLriJTvnzFmIpPkj/dfDXpl9GLHYNIRpcw8lQKA
SoRkVGTqgYPBN8g2M6jpAbR8s92cjJXnbA0k7+q93kdz7FvWH/hTHgJbuoyzVdtg
J6jNCPLvc2wQjBPdrsPK6qTXlxxF0sKGeOdsmfy6e2plofFaNcnTxV5wLR8m/OHH
vVhMZGUa+wC4kG+5cGqR9Fw6Pp45Sz7Vh8XKT7brPbuezpXlqERXhOgGMvgtgtMu
9VwWuoKfM29RBVDnDyqGzD6sWBDqR7C9V1duHhLNIrB5AB1QGY+VHc3raPyOjV1R
wv8hjh9EYgWxET+MZDB2NAfiGUowNSTxVIaOPdCDXV1E+kkgDAr73yD0ZO4zBC2l
Hn3sbdjLcCqq+h1ZTzXgIsLguBci9GsNFNPdUGmC8ccrs4Jg21cBYWc1pr5BIq9B
ij49pzEsmUtgwbhoHeIdB7y9mzWvsqI/RjhMg0eFCzO5quSgRCh+Am+2Jru6hKij
V/wbDT1s/0FsJBx6OZnusYKcxAs4AWuIWLrCAlXxfQ0kTRq7KRh8xnpsp7j6MqkK
ImZugsGvh9abIt4tij5XMXGjNgVjarz5HGfoeF2X5Ac7Y7jpQiYIBHmqjUpl8G+f
Gkx+J81CZhYgL4lk4wkU8SNRl1UJeQLnlxzuHluoh+jJ5VW3CG4KExlG/0r7Xc0z
ErVgeTiL2XQVBwSP83bCR9zyrcV6NJq1hCyS4wTjF8gWfFosQ08VRpEFoUpwS/gE
MBjQWUtiITzvzqZ93EZk1Msw9VkuNtGTzpPDUyxYZbkXmHdX87bGQ64XEP36eH0R
0yXbmJS/ySa3hKZTYTM63EuJ+DMIbr0G3bqMc0QDJO0OEKfllKbLo1o/RTdUocG4
+qQ3faKVEu1IQMffVVDigI9aZIuAd3GHOBv8KZ6lcVJlby1xwLtYnkS8zMiOlLHB
F+KDec/NdpQqz3I2mZqqOxADt0Cx4K+pl4lO62ylqs2rreIAsBJGYiubzXNVBpIS
9I6PMKyWkSU7KQSrpV7Whn19kUWcp217/SjD8EW6qKwQ3YhHltIzepgsYXm8q790
oN4QRAjRSvw7g1mUl38uDoulmy3WStsxmwlJrYqE+nyDdVNBnrRRFmWpni8zd4E1
Ho9dUZEKE5/srGmAbvhfDQ1EXgT8nwC7vI7/jnG2u8V0GDG+0FqEj1OYzHePa2KL
IJZZ/hlksTSX1nJ8xAv8JoFyhYLnQn3zNhJZ8A5RVSeDr9Max9ZUT3hcH16i9UVs
iqG17B7vYCiBsoDebWhbUqWH0Z9wFVvwdVbrdHGMvrJBL0yIvwZkEJC+EQtD/sev
9qWHv+OSHFVeXmYWJQ65nC2L9ePqzphdI/GO/BqC0jlqdgN5mk1GWN2/ETODBXad
usU7iwVQi8Ttl3/u42NjOBzdJqsd2Zns6RuIyZ4fNQ3fDKOR6RZ9yQr9aVyJeXf6
pV5/hwQ64kQoEgEXkGTg4BkKT3x35PUofjH1iT+D9aZmcNj9ZE8SfOPQGUEODYuS
GIaV2Xi6OaIUxh3XHiOMLaIjHYHCnZThk1GjDb/h1nG3SBCxA6DROGPf4UmspPP6
bmEgwBjcjGEjHqdR+LXCa620lkuCC40KceTsBFB/jKgdcEE++kKoPWsLr/9K2ya8
CSprRSAo1p/QmZ4mMx4DLszkOymYOWowvgRqaaR50lEy5GCLH5cUCob0GE3UCrds
G/A0CCuPjclTibDzRfK8TO5TEC/7iQZKjMLbS+c/Tt3FOqW+/HRLGLZP9Zqg2pn4
TckBnlWJ8UFtZOWr+x8T56E9DR3lZPyFyagYf+DBOXrp+BLdgy5yfeDEaaACiTjk
WNA16iDzqzTXvF5uZd8gXSjII2p5zdJL7jbDfCq8osafrckrMqCLnspFRk8+6ILo
Uby06qyeMeB32xhotSWus2etkAigNOnDpGOX35og6hGexpaXkU/qNNKYZ4ZJBArD
vtdKKMuVhY8F6AbqgVre7ZTlXedv20pd8Y+OjROk8Auc+lBcddTrqbCUJ/92XeMF
Uo7cuiqlal31RMijGQJ248cqf5RHvpTmhHMto8M6/Mbl7+Vw1552k4vVGgGKh7E9
LB0fbZAjMBsyozsF78dqeeFKp7qn9geVCWCX/WX5vZXq8HQJQ7rOcNPP4n/0hpRl
DoPWkney+72wEfWf/MZ7mcK9LJgQ0A27ZhOyBE9VjeY3roVZD2GiM72Bb2yIKfv9
h58bYsANbkuZg1Vvlwj6RQjYIyS85hh5qpSMSggBRzpDD2x0S7+x5yTxmcHYWxbo
Jwi4bx49PqTXqYt5kCQaFNhjKb6LPaevwLRjtltHgbFTWOck5Rdm4vm8njTP5G9m
l0R3+ogKNLBCFJK5TV1HCVjPiztxN7PvfEKzGdxW7JFGjmj34KgTidZ6Rkz7G66J
bjT4Mq2ctIg+rW5BYm1hkG5T6MKLED34eVoVw/mNrl5P1gYVQ+u33a3ZwrDnkoKK
ZtV/pZObKG+6YS+rKaR8cHjTOQk4A8ddshoJkWk5UGWnaPGiXa5AdLKborHizxbZ
axdflrxxyLKhgKADbhrDn7urPtheuTrMvdWn4XIs3kDlkLlQDMaFW5prCOdaJ3EK
n4jmJv/G1keYqGt23YTanyctmS/OWxZCe3IMnlbvQR99ZTfBhYzCfAo826qm9Hm1
pKNskSMxcWv3SafBcfY5RVHbOT/Jrd1gNBKebKAb9rTN2FvDZQTlCU0s9Ln7RKSo
u/WBcvrGNMC+6au+7xx1iD7GBp9oJOdm0CCdm5ai9guy+avq7LWoDZSZolOBTuSA
kms0mRkwMeYS2c/67puQK7pe3WHNSn3wjig0mXs80fB9iah2kPlbh4dnL9ckVNpC
MF7WLLZcb1uUBbkkBGZFJ0a2sEqFK2XmhJLfklR5Sa6wUG4M+q/jnv7lxc1RfYoN
Ym4PkKldAp1DJ0/z79hpCnZG387YST+1QQpwLZU00qKx5AvY8iJkOMyTXT04LLCB
7lUSNJtvPwh0tb6g8im9Jl0djE7Z0+NOHxWsOe+ahTGZLJhUJet3LexlLdlKWM5y
HmDHUe1UpP4cH4HJL1xsm4a4FR/rBCWg+pgWCTkhBxAFPwaCxE3HqgQULMaBcovf
CxXL62DtEcFu/Nm+Sn4OrSK+uFULlBSnwAb36RtOFpjir6b33GxAbgQhu7nhjbFH
gckn5xPaWNxHTK0iJ7CoMbj/TJCvp49sfzd3oES84TYNqKWvdCyTipWWVmjCfeOj
kqcMOmIGovp0QrHVe6FLho3ivmwWck3a5Iw8w/ljZ2WKXNMUoyef06UpNBB3RXQi
6Ere8+QK1SRo8SIA3uGhlsX0h8lJb+KYWDQYR6MJGNCWZHtZoVwk2YCyra8hnk+u
7iHF/EitiAYfFQfe/82rwYyg6N177c2lHF2jwXoe4zlrJvpLa7BKUuFmFJXdyGc/
EL/2L9wJ08T53k5ofwRFwPrtGMqsBjTGTejBWJo9G+4dmizfcPS5hgJyYGrf4src
PSJRq8MgAwNt8l/fH3oe/8jRXBW32pAMoeZGt+2qNeE5zeHq0CeB127tzsOii+xj
xgCJTg1C4ToXas//b/gFZ8foGtCrBYo3uZUTm2lAe8c0LgcMyoou7N4fl4Efbwyb
WtNkztsYf6dvGxEhHUk/eGzbbyP0IDpWEY2meBupsZ/1BmVGmGa2YvfKSkLpS9jT
LecyvPaFQmy8xr2yJoARe1nM4UfLs3lQ7u2HN4ogDahNP6Gd0IFUlAmL9V6tvSsR
7ocd/uT9s1AnllznF+8fK03EqHTfFFZCCH77wveuOPaw6J7PrXYN9Eu+EzvzqIRe
m9SkqRQi75pJemmdz1asqm2A+9jVDie2NORfWfCbDJkFhWS66cvNLZoDG8p23jp9
0aSEAUuxvvHRpt80YqYVhFnEOHVLEftB8mGDtdfa+8TF5ePtARQ8qKftANPy1Ujw
EOSjn+sGfXWnfQLegqKmhyACsxRGHPtgWLRONdgibPlvFPK37PziaNQOhDcNHqp6
YlscAxCySZFyOzeO04+b3jAnI96JOS5DsmQkDi4L3f9cut0/P/ip8AMA21RkFZs5
BFipBioT6rTe9g0/niinyAXUHFRCZFvdz8ZSvLWsuMLSV7XCKvn/TCkHUMVVwWPO
oWEeVc5IoSlAPSxhNIpsvq5Ov3YTpSPUtcYhZ1iFHdju3A0QhikSUyjYcBPu2AFh
aMrzomgbSso/Z3UXqVi7OBA3b8zXWDgiUZ5bndWWQbFx67eRFDiIZYycIdSfRzHh
GW5oDqsEkqrX0ihMqQZnvkQUUIlXBzw+DC3RACpvxpoJUFENHt573Y4wcweGPzm3
cykUwzfBqYdmOTsGdMpexqsvlhl/hr/fHDq3q/xgBiAilri5xdCM35qA47Z+gPw5
4ds6/rLccfl+G5u6c6VHq1EIg6XYbWO5U9jLbMgBBP4fWVBEmPuKUVtZRBgqEjHl
JXmeyYNseCW4Pr2sog67xcjHAOpbEwuKzB6RALqmJxFfq19bsF7ZowkS+gRfWFb9
2T3f67O6eG6lxXg8xhkRwE9uz5BQlnEbYvr40tvMSlACFY380bV0BYZ+O0lWXcdy
OghR6Qj16V+cajqYL/Gm5aON3xxyQWEEMEwoHonXLhDb6+mHdb3rLkFklm7TR6Sb
s17ySeg5vR/E85RoXY/3m/vbVtPiiPmrQdrfa2BS2tlLqpK1+XG0TPiPevIvR5aC
bpZ65n6IaIfeArWT69X2NX3oo8MDgoEzEcx3mwB0tndNTti0SwkzdvQKbQdKi8Uw
OyWW3WtGkRLSKW3l24ugugzQ3kcNv6gvBULSxiHpBHvl4DcHaXswFNZ1dkWiGP/m
ERDpgzJmjuKpX+VLv9r10Ujc8cyfVzTiZhz5dQU4VwxKAU8Ui++D517WaYT5XMf9
M6IQLgvki2BbduHI5NNDNy7Jm2g9vZVLMV8UVsUXS9glUi0e2vXloQlfJgin0STk
XdROkfnbQ4h3rzJ5aXZO7ajPEzdNe8RT5nNnak0BqRKy+MGxj5pTfGfk7+OvAY4o
eID4A4uvfCijqjbaxKSv9QLqs2KH7WvRW/I+q0YS/f7G7LxlckqGG4OYFJzFZGq4
PNenHgdfG+AGe7B5wpNGvgwp2Jy/DYH8aqfTkAUzbM5kt5GOjiVqWNwisfsv9RN3
5DqE+V1sh4Ua6lItpXLLO/CDVkfQ2VRDqg/R1DMljkgWRSv3B7043Ua7qmdYt2sP
7nuqQRuftfg5NWUFKbPOB3y89u8hnoSdOnoapxBsxUu/7qznB9lQ7j0D4qXj4ez5
lwTGUMtCVYxNziHb0mXV8sA0O+Vp61OUBCThCiKGM9AyEMeR4iZ10C7/FyTJxsq+
o2PU/e+cmmfahzjVRYH/Ua7Ohp+GfuxHLZKX6et49eLogkQaHFKpW1hOsPV+rwny
Vdv3BvdCJjc2Yk3I0Gwl9NzE8i9eHu1RaOi+tiaACsUJDE3rFpW1DAS1t+nsGJRb
dTfBfGrKCM8Gais7c4tL57ev3MO21WoJN/Wu09n6wSAUEInUha9j1xcqbIERtJX5
NrwefyhuxKL9cGxBGS7+EROOq8J2vbsN/fug6BZxSy/200zQhHVxXvqc5rpQdyrd
I19DBOpm8sL7raQFQO8LKa1hB0hXUdcSdRQVX1jXAr9PN1F84kKmHjSEwo4tMQTY
wV2o7jhrTYMab5UxYSiRG1LjRJajnSWb0+9Vof15zGjYFGGpYTdb5t63b+ji1od0
ZQ+ikc8YjGfIuTR6vUShzMhvgcd7cWkjxBkdtzLKrHsfLeeXWqRmAJhJee2f5+ir
KGsGRP0Z93nppscJcC9Pn8OWfrAC1fU+p+zKOJtde6DrOqZahLirYyMe02QgYaM4
woPWeTi1abVbqtgiJzooHfRi3FuwTtvY6X6cMVv932URUwQ8+WIx9YSaHkPUiIDp
KxahjqsygYVyK4xf/IxtVAenRJGhAPJJ9uD7ITSwEBlN1zqIMkgGqN352FomspjZ
BrUpmso4YWIV30vV74B9HJnEe36vk6j7dOSdv0sNozikhE+HfjCSztF5uGXRgMGj
eW5NEQg41lFgLz8xQODuXitW5thlSiiIPaWgUpQ8C+ir3VXfpEGUSe6vgb0t7ApS
1x8y6XDLeHqHi2FOezc5clMzcljhzuOL6f3T2qOvQGRWHHZ6+zzRyX9Yvd+FhnMA
AhccbYIbOL0+GnLh+OB8ojw89uPvJYdbnc2F0aWL2mIGv8Fu/nLZoMLDdu1Ygy/C
xeFM7Qi5d4XDf0U/ku7fWz9RKOWMcpQzCVtpdSGsV5m2N8lH6NnqrHzTKTjibE3D
FKX2fLvEVJb7BmEZtIJuicKvy0ZatmgZEKpQHY8/dVSHpb65a9EW379EBpd2Q1CG
w7zex2nND25BTCUrn9CoQBPHCtT4xOxI1FTtSnqu98tlBiiXCHK4ofvkgZ+PTZJV
cYkMXcFeFMj+BO5tt4cgUi3Wh1sUZ5tTTTMo78C6XXimpCm10J4Z4lKCSR9ldDca
+UDxuESdzLTS2aAB/Ibn+soJrTB+58zW5OoYqcjq3jg5mcfgyGF50DrDL2GE9ITG
tbN6MPOcsS8JSKbcatbK72A+7alXD31T7dluzATLfWOjzIq/ROP26QelRo4zXdKs
hnJCIkjPckBESzwp/Hj+8B6BicbpeZWWXOcFAqd4ZhhmFROytWs4w84dxqQYnNs2
mD5pk/e5rsOHjiLXQ9nA9J3jqH1NqWFCCqCWjrE4AZlaW5N83MV+KfWvT8mSbJ6T
rAWQK0luLX5RAGrWUz31T4Nl7IeZRRQ7k+en+fOV1zK7sCmTW8Ds5bkm0lTmV2P+
RYQiTMP4G0KpnrOmMiZS82V3XDZzrmQvdXF1YXfwY+pXsfICk/UAG919Ew8I4IKk
AKg38Xq3vTBRopj26iXtwnAWNjJgZ8Av77Ys962nJc6sklT/xlRnAv1v61yQGttI
BblTktPuijloXDBWPxseRKY3CWSqqEBxHgswtkxEuCc+ipPbqaMucClWxQG3MZtf
O6x+FA2oQhgYnpAQl3XoD2zyywl8P1imA2XktMMWWhVU+bJbTWFdh9szOi1hNktv
dlKlbfMYHSFqE+UCPeofqKZWfH4rQtCIpMZQN7AC5WLvJPpEKBqnR45M32p3XwVh
Y+pqNvx7dO7CMm2li6btqsYyHK7g/wQvwH96ZEMaTo4Vq9wKTM67AaMJZmIIcDfs
2Ex2taxlUyHCQvVJmPW2zKNJ4PtpG6kGvJmyvscb1cwg6ZzVv6uyDvOktlrvl1+w
1Of1sxthJGSjBPIHN8YT+tdwuJ03yFfTeUzpcYGS3zl6AKrWzh2YTG6rPeNQzBvi
QOf6eEMZ27fhMutFEsxDgGMNafayNd6sxTWngOPbRWbTrPNTcoSIW/Sff5ZOI05r
eJdBoJwTofTqC7/c9qG4WgfM2yBcqNESoGU39R9uNd0/6ui6Tq8Z/UlnEbhaDb6n
2BjSHbOezmGo7XqcrjWeAn6VHRmQJPVOltOrmEb4rw6AAsLQhC39xSlNbhALpml9
jyf0qDYCJZAzLRQD9GpQHKZrCn1qoK9n/LEUU0qcELRxSGbroXY7rEth56n8uSfE
CbrF/k8LHlOJLfwaW5ddtFqy5lsl51j0KYb0dutZFyKHMmZczqawOyKcc9kZ+yCn
jSYkfU+xddVaPcVAF0stAsEhdb+DHbGMXhHfWA9+RLBEmnBsakikIjK5Y83l9GQc
Hjviwoaym1/dNmb78rZUI5zW7LJ7y6OCuJUHEDHZSd8V7qadO9GYMVxjwUbavUUJ
b4MyFvhSPS1zqErlCdwI4xo+2nbc4zSf9/5F7UgkNilMXoftxZY9xQXlCPrU/F6T
zdxMRsc/nTIS+aIN7m628Zr0PCv3Pj3ERDIjSoPl04wI3p8K6G+pXL5ickiV9nMS
iUfZv9xoddd2RdXId1DT93g2oVvLiMgaxL8svwjyNwmJ66glqnEuKauf9v/NMvn+
LH66rVcF3V69jmNhU4yH0HZakYRQfcjhfp66lRucY1GM2Ui3n7/zXAjK72StNImC
ndhLIcxRkJpMj9MqoAQbjAhH8VLRIBKRYg8QuMkfLLu/YUF5FTbgXPy3BZVxdnn8
lZyFVBPtD9gmxhUFB2eXVqM6UMlb5/I9AeCIj2s1hefaR8DoeayKnAVvUulKFEBG
/5Q5PSqv4Ixl5EBqUuelbvLoB/9e5/rk5jYKy+PJt9rG+EIolfROLMti8LisCUe6
+Non9m3EEgScKJ3UaDSNmGTJCcNsKDyV9+f4tcX7dyUfRh2EmXQGlyz90fg1C4gR
a+Cmp6ihjPJHDoaKRFZldB3ITOrEl9ZpmvO3jf7BKNu5cP+EoEgGAR3muyEB2iFs
oDxzuxNmcmALTrJZUtEIpic+tjP2op3h2+bX20tzYAR49LhhSKH+0QvbkwnYx2Lg
aePkSeJokU0w9uUc+miRrnxp5+gJmJoud/dTNYPWO6+aYtyIdbhsugzoh6QlvEqb
S2zFb30Pev+GcsfwIO5B4/LiDfT0nbWc+mDzvRGyr0qiei1FYfBEd+Qt4JPCa8ym
eZrFBNzq3CR+80WJRQ2B6v0Azugw9E28mt9fKfcm1DZYgvO0aoEKlEfa0+Kra3Od
xKXzxvkK50l1fBPCqhxQaY1/l3VA+sBTJrNkjyM5F7UcAFVRsik/PtaMTxchR23N
BdYRZGsBN1PmlT/JLvQyrFin+oCeogoQcJHpV16FyjB4Kx7lmMfqlwAYfX7/l5Z7
u6D/xdWBCPlzePmnkLVZGACkkJGeqGluwp/istoY9m6IUrMiiGBt9ABUxXjtZsVh
y963RBdCAnRrrUJi0/A1SOVRKe72vhCxpXslYMdfOQZg8RbTsVsh6jAnwqPxZWsq
7xmwCerxZgosySbMw7UsPUhM/1sCiGes7F3jqNwbhLE7Sxj4mqmSeF/s5gnIe7Jy
1u+5fouS+/lzYmYo1ia/cUt6KYrA6nkiosXY9QNlnyWAzrGdcEsWNDxAdEybSa1q
2TXqDdetx/wXwYFx0zPEP6yfTPcjNMVgVpnsalFP3EQBWNt+uEjt2oKLmEYrCVV7
GLxW9MEXfPlCV5SmzWN9yRC9TuCLYd82TqjEppfimQx1idLLPsn8Fu4aAcD7O5CH
NuUfmjA7eyCRZrgNK/3Z1fM1ZY5xJlg+NkXDg4wsxS8ZKr6Mq4RfLyfLj0QttmN9
UXTVn0QhxKAML4if3LB5YcGiMY5eqlZ/F9D9ju6ZN6eZkFCoGRBTSzcXiHsn9qPq
7dxnAQi8o95ibZPbaBVLz4j5hVTmdvskpMyEtc+CMl41ttE+YwNOZjaYp2nkI53s
tEvtLkyY+CmWGcXm49lSyB4hmEvC8qXtTiPO8BciA9X1Q4KKBvqaIcWyiUD187Vu
JNbnlHopHjVmfoi7TzTNCa13r9njhkQ/lwTMoxOdBVlBQPQuTq3U4sWMlnzOdkck
yA4yZcXJAxSij4D7kZNUcq9gdVIah27cW0EyG14Ldw7kMhusmjmz98dpFf8Gk3fi
cyb/vc6QDgswo/XzGAnQPf+mvReDhiBp2I0pS7VRjeO1QEMMmQ2HvgZgIw+jUCy3
fy4RtblAAdgFevO5V0F4OUf5aTp+brd+65VDPMC3oln7s8+7LBnzSWC/BWAMvtdI
c33WFO8SWgdYxGU9sP81Q2rq9VbYeJpRZSdyWoQxiwpQcBkWDY9gmAZM2QUEVsfd
jFNv1PiLFsY+9WuGHDiD0VPih2LCbsliWnimfJnbPOqjgIxcvOQKmozhS7j7RkfL
QjHdG6QSCZ2HlkH5SnRrPwaqD1/uba0rTS67yt73yqzY2iGfW4niixBNYrc2H6xX
dPfMNI7ZyGp/gY/GLAmG/6yQV3CTo3tWX5ZFM9avfNXNiHNm1airHP28POUtvI/s
X2PCC9xXMlMHBjiwc/1yKNNku8qr5ZgvJ3G78yYRhsOhH5KbkJ/wFl5e7Ls52q3/
Tu/WF0nU6ou3rAswBy0OdT/zS5XWm4/fP7D1ICdTYNeux9cnoTpqMvvK7Y8gpd3Q
XnfdCnEsEl4nFDMNg+1/KFY0yLALgpdwbnWb4Uhqiu2J0an8ruIue2no0FZf2p7A
SoHDhiUROQgnGIpJvNC/ycjTozSvQwpyJId+CdfLYcjqKC/g61NwjgdJRCJtB1jz
BefrcC3K7n3swYTyQpPB1NalGTGjLV7zun0AWDC/k4DNTGgbM9AfZktwj8ULtTAT
gwf4bkSe9PttUJVZoGi89w3qonqV8LZPbIuzU2BwIxxBNH9dDtZTXe5CFV1ELpkq
5+bEwkuJIgn1dmjS3asX5AcY/Irh4R0ar04CKHlmUmIFdtRkMXLszTBIVghbInj7
0B+z7rek6JJFrSoAyrF6Lao7cJUvYw0MtIH0gj/wkcaRIsls0Zkdl5DjbgCzGUto
MWq/yy2M1KFXArkKG/HaKEh6mKV7Uzf0ucBiAOj9bCsdpuq7k3M+okWhRk3ai+xM
E+ZvmCYlEfeFj8aD//ZtAoAVlVybUpBDNT10KEcMZ4wDHoK1h99bw7yQ+97R94ig
IkQzcmrUgxPyz17o5R4cF4JfNJvW9FyrJQodPvA0nDpxJJpkvtHCdwbIwTARiqHR
fEdRS6MEXKJHQ2C/U5o3PH0JDBX+jTcEVvuGcgQt8V0EDVPwX3/KHLXm3XV6JZSv
mpVhhQc42EZwT3m6Mu0WwraPR/Zfvfb5uf8VGhku3bj5PgxsBFAmpKtJFXax9Esb
s2hbyhPWljn8bFM4KjjPo2oREk2SmHKzrs/QL3OYrwV7v63O6B0s52+DhP0iqjfb
N0ro+dPO1cbFvDZhSpj6Xzn6YWTR59strwjpVS0j6yh6B9a6nvRs7kXTw4O3zek1
UJnW8S1XgOTxvPe5zq2aC8QRlQ7cRWjQc57QJr+7K4NH+f9m9e9ENm+LikQQBs2L
vnnjmLrUyc743SWHW6sZUmS24VI+ht8Hbv24rlVS4NCm2ntM9CeS1rNiWHvlBCcR
OgaBpuHgpRlqwLYFKQt9OaLaDcP/rJUe5gJpV6lXJgBDDYbXUac7gtJZC/s19kmC
MhbycJgkYJ+n4O30HjptkGf40IIx/fM4H/LzKt4iZNAwrJdcWTs5ITuTESKL/iUw
hwrRsrUf9tneXfWwOyJ6N34XKRgJeO7lLmqy37izaOlpa3OSGqf1Ay1/56UKRfRw
DMX+nx1xr29nlplfKBKQxJufRtLEsamSzZCAKj9tfscM0M8w1JkZIvD2qRUzcToH
cnckAFK36LL7bcbC/8zmCdGRd5j09fzFFguV/XiOBKTLyJUcr3MDmTMcs7v7n6o9
ppWJzN4jF66d9l1/MpIL2ElgKpcmceoS0oZLxK/iILIoYgfRAzxmk+LKnAG4DPoL
RcJuWtRAkgIBrM4t8ccCxiNBDy5ybuh5RsV3UzB/Y2NUo6lapOvJY2VLGlWFK82e
I7HX1y+Go3vc8fsOGR8JBQ2cQWkuxlcfOHn8bkVaI78iSgeNPUTAI6l2oFJ8cAuk
iuN5aWc9JlI2LWWq/wX96bzSU92jCobjGJP9yF2jHOtldG1krbOHiebsyY2Jdk5h
oKUPF8krWuhi0kCJGyPW9mnACDhwR4kQTflN/ylFcr8+PZ06R/Pb+XUXe1WFah1a
TsU4YS39rX6b4omkACP7JvwCMr9P9kxz0UzcVyDW89+2Cy6a7j5Qc8XbTSfWkRPd
Pxp76m4pcgN4uK8e1pgUXp70vpoUkAfAFmWsFqUkgYjokIg9QznMC8dkxhY9/sp/
hmbtka1pXFqRA60ENu3KPAWNH6Zy38VDOVVXsvQQ/bZTyJw1SySvGI2TOj675DXq
qqv0woEJEfYXc3jehZ3uwz9PNoI39OdLvYXvrElfYRIxHdYpnNVEZKfd4p0wKMnC
xYX1bZ7WvQ3RPHcZzbnsZQSWGelJoV9/le3uBbukqtD/o3rjDxL1BIymcOwMDp5s
fquJCRTTyb14WwaWp0zWAGsgjXcZhdjEmwQvr8e1m2Q+W0VWEvbT16X88MzMq1V8
wS06ixwzYdo2Od/J6AuzChoxZWZAyFBqz1UpXFbpuvQUtcuLbBUtFiYTHtooRfoZ
APiJBdRR7f9oH6JSA33XLMrjaNb/dkJbBFvyX9rMTK3gA3wdthE+bGzNeDaJyE5Z
/vrSY34dvAyfxSyj76EeepdHSKe9PIKRdyckU0YKyPKNL7z54/nAT//G0+7rtXwG
nb5pVAbehap9Z0PcQh/0kqepLkd3+Nx+Sve9Z7GPxBZvFos72/C+fG8CpPfQ/pv+
UyAyESRQ3mTdTc+j8Avt2w6JRqdps9jNUsK8Q/1KjUOYLsa4YqOk5yoMeeAK+mnj
Tjb1kVNxPrwZKo3w/M67SFTLC5NyIbtM7aJv/r5pU5OaUvSbYiUGqnvGF2UWsbJV
TokX7DJk+cvNcrYPdTb8BPHkU6CbGN1a2pFGPBDwm+wFQOC58K1Uxwble7iyQX4v
T5TZPkDV2uMoys3QsoI5vS/kzkAfa1/F8Z0ypF5cnwsUk1ToyqPmfVPPct3q2wTs
81+0vIgTvclllZGVmsoAsSYC8ScnEVp+EN5lQC+auVftaANS6/n4IDS9Egwky5NK
ZMXCO+uNdscvM/JhqaJG/QBai55LhsM1pr/Bv3luSCNnwTZwOpMoMt7XeiLnOFtl
7bAyeZgP3v7SCrFNYCOpCeyLQpzsoKB0k75yeBHAe0QJp37L1FoGnfRUnryLZKEL
njBkHWBrubsMzLi1dazaEWEE4RqVuCOU9dmFE0OI7AnfwMW9hd02l0epDUNC3BkS
HCkM2g4MFt1Tgv90C40JoxjMRgWRWuy8yfWeGfSznvUESfP0Saka0qOF/rd0T+Iw
SdKV782tADoJv37vIekVCsJValzz2WupHXMzZcXkH/cuQ6yY+PC1YpKatka7MLCO
pyPm6PQ8vCrE9n/SmijqLkkYc+tbuGkI4ywyycwXBdxB/oOf5s08ah9oP0F9/JcN
eTAQY4Ndcf+tL8dUX8Sk03uHoVxXchrllWbvyYaYNcnqNUZ/9B+jDLHaK8+abHoa
Iw7zDnBUNayq3RY/k/IAG2CnXuSkA1OSXPqPPMMJmXb3XmfgNnYbS8vKwXdRrUsb
SAU1m18XBGGIeo0pDeQdmHk5D5FTNzCdqEsQBfpGoUfGmp+pt0RYHmaQh8CBOCcs
gkQHodv4GDb/Y/CUWIqWRmZXZrWDrfIPpT4qkDFa7P5ulQ99IKX6gHDZNRQRpLOM
jJXkCLjAwR2EqarzemUmdbC/iXvdOwKlP7DOAhg4qaoKME8xP9mKLB1cXWtOr30s
Opxa6lHySdbelbAmDEKsUCJNxTKqzHZrB5CwdIgsqT13I2epR/4XyrukXEjgxVIC
B9EBTNK8BZz0ywCIzWlAtBZta93QqhJPBlkYtx29cJ06rRzEo4RgrpyWpnXrRZJU
g2bSOn0FR1b8blD6aZVNZbdZHAq1E1q6SMurYuPXcs95E7lIRxm6F4Vo3axJ8Uia
U8He2QKePWg/T3xtW1VlbYGRBUKy4OI0wQ/v7uFCeUNmOhARExu3pMslp6YK8w9W
sYfEwsA/aG//ykfQ/u/LOHGUm4k4Gwc9Yv2sEOdcgBad9JAlMVFT2UUM+E0Vqe5I
ry9C8A9tsf7TVCIPgRud8FLwCwTDC+MawJ78eNWyfC0IZczVMg3fcWnJhVDneWo0
ns59ljNfXHH946KtnWWXqlNiuWkVGcztWfOhxwO2+QJ9ydGO3/Dy/VXMpLEl6R0R
vF235dGTpK7ybL/A6RVVNsEw2safHboEIAzH+GBdSMJ6QJc0zJBbgrVv9cDy/BMz
4wRmIhvThTO4aJbjLNTFsulIPxknz61ferZ4AuOIS13vrVYujI4mTVPfSdzVOOAu
k2c59FGEA80jVBmrWHxTwYRtFyP9cvZGGxuzK4GPA3+8/L8G0KgBwAatcp5WyA9r
XnrTTHvnFv7Pds7VZUU77IUH48kuls7DcDqwl/WlouYLjQGQAIxm8aJWw0bLp0Ew
gcpTVaGLHtOErEu2w5aHFPFoR3zRyiprpO9dQKteBUDsUbuWYys0Kwu05cubtozf
5WHOcbeejt70xwnzw3rIishUb2WUVlchmTBY+zWCJFlS7rG3Ol32inQTJDDG+ZjA
5jZU7cZyWGZ4VlF+Eb6hrpc9jiAee2YE9P/k11KAa+qGWactNiS/iBL72x6bUu25
Qpcp9Hw25sVWI8PKWX4aJUkWGl9KjZqJ1catqh6KIEY9OsFtAJnjnLtXRn06JTy/
EeJ8xuSzIaMx4E7SVOhjpDsdMoOte3TPH8KksxI12nnudGi7rCIGDdR4rkyTILrT
bx7WaysORKQRn/xr3DXPVZc8i0RcNRenUiEpYIGr8oBc32POK/AxioMGbtmW5FLj
jFLVuO4EBhG+iZVdpSTemGoRzry5xF8D10YPP+PE6XcFaCg4GHjhIBdodi32rwt3
ucLPIev3W6chGxA7BMKhx1o8+d8CnTCECePtHdHPNLDSaVPZUHfDpPXlR7RQ5C6r
6kRp2UT0Sl5ty568yF3Jwmrj7QPIH0kA5VnXK9XrxnrEfA5p3BeslMqvrDqCfxBZ
nzpRjBDoHk0DO/oD/1ybJ2kJ0GBLGFktNi2lsabt4/fbRL67hN/DkAr4zz589nOK
w7/jf0pl3q6ubyIeRhuLZyOyX+5YWt4PM8iMIMvSeYTHzhw5/uybb6LU/d08KsCZ
mxGtN1au0z0LRyuguX6pC5zR/dLj/QlNFr7p9bMbUklLPPNAnk+nDODAk4nCnOjk
9gRiilUlAcZElzmKizDg6ni5Rv6h0Iymf4Qetrotk3+S4pxBd8Y2xL4yXE2mPv0h
Yz6ZPMjArbIAZbQtXKVb+G9osiJn1Q59dAFl97ZJ9M5vJ0mEeSllEaVlqplfPGhB
kDCwj4O3vmOV3sEu9IpWvu6vXQ8kqm2hVv5X05HbXy9E9t+uPK01/SDbKadES8PO
vzlXzZb1YMIgMG/6KolX3Fy5erGW6a7asVrSF82A34DYaDl+dEMVGk8E1ar/MYVL
XMxFwvfbV4XdvjTVQdr/Ua0gzcSHca7QoA+yocT1EC5IsVQf5F/HpMWNdMOi+NwZ
H3mRNTIF6sif1Cjb6Gob/oRCO3AvYFdQ5BPGRpAB76zIYMYpGFMcvg2Rqu8Schx+
zSFI2CK0N4yUJdZjbPnLxH85N0skPIHFDT8G5tq4Dk9hJxQtyvWGoYFi5rStAri6
rRKiHyMouAm7G1tD06qMoxw4yXttFI5MiSqjIaubmYIq5El8Ah4C0EChD7DHPwTo
IYOb5UTJFacH33DMG6BzWF0JFUwhWCWEbCq57QNCdWslr5xWWvo6sVN5dkdW5bkx
lLi1B5q73Jfg56K+1DKyrk7kpN1C9lzLlJ2NDPwhIaCnVkXCdoPQkxWbh5YT1zaY
ZB7MoYxSCrsCDkB/MvrK9gnGagPl9sqzsf7TKO28p9Ysvm3jPtAdf8XpB7uNaY6C
Av0nKN7Zc5VqniRb/xSo1VDTt5DjQjgZmOzuVOpy9Q30qtdwnkieS7W1u12sKIeF
/Amgl20B3yB0V7yFPu7wmHwzgB2TvbgXtRFZ5enEBF3LGgO6dH24760ZOiXB0LHb
cy5ANhjkqN1L+jWtBkzqdGqGaUQVejLfygBmhJH0jTej89UpfxszRxRX/iQs1IvR
uddMpTfHN9cgzXHhq+Xa6g5LCrAlDiqDfAvye8ca3b7YpFc5drEWa//GdVE24QTb
GXA3Wo551+r/sJm3hTsBWHZy8VogavXO16es81bfpxx8vxa8XZZct2ZjCPgzHgjd
J/i4+QiQHQtijTNWrD7MHPoCoG4L7Dl8yzk3g4mQI5e/rBYhoHIP9cAmTVyw6EKZ
1BJGxdWeykM2IhWdGRLoECI5rEfzGbIFLZpZk9Ch3i7Dz0Jn26qJVD7Ih5yQbI5T
93CIKmN19CcN7m03OYQ7DUaHnaIyEtTEos0T/h5/uTnEAlx3Akamc3JLrAb4lp33
xQet7/lLHvbBtvNUOd3bOVHZaSJgdtmn2WaHKGF5MgBgxRbS7hIsLQMg0dyAWvWC
hklWviEQcir5TUTcma4OuHV68uRgE5sxQhZrbr5qIGALn0cLpyuDG/QU3dV3s9fv
mgXnxIlc5gnecib3rE9mo+MfxV9gjcjLlpL71MjquE6UCeIRPrJQuw3T/CKUMtzM
C4Q/RS+qGLDO3cJN3wiAK8HGZb6hONc9LZDQnYTMSJn7anGYJ+xK704YzLJYKmwD
LkOUgAsdD5iPttjjh5m1hkFNUEJGczMReofdkVLoGZflb1WfsMwjFYVObYVIByzz
S7SJgUEjkPzDyWeOeci7s1e/Six08g/xnC5DlEyUQVwPylxaqr/S5Q6kgnL8UoAf
PURymVnRrhblG4DfWYeZ/oHfvksqYe7+EKKvxhLLgDwkHRXGe2FyDHqqVj/VapDj
jz2p1E3jMrwTJC4DDqWMqyBSLbrpgvTc7RAbt8BvLjrCsRjzwzLpKsOdiLu/E0Fp
sNwOekWo/LWqfbdnYXeK080dsxhdBd4uLt+ZolI16JwpJIyen0F/k7Sk1B6v7x1E
x7/mx73CPV1V3k3IKVorR3igWDKhCfo4bSteWXeMh5fAzQ/wbIOH33efPaT3EDlw
maP1WgWsJJ/bd3bccdTEzNiyrt6w/XMxZKlIAyyV1BZBjLvyXrgYDsUkFbj1IBjW
4cC2BRTZthGDgLHHG5DrDrM+u/CaUtoepDbQbOguGYc9psyHObCxc3WAIBFp4mzK
cBoZXBSXANuWVgllWWsLgkz9qk5bgvDa0Czp+mGCwBvcbjX7QHYxsSYM7EqPV5c9
1OKBmOYjUx6OmFnWgs6WniWCufPuihd8V63xDPWd/Z0C6jnUh68lflmCTWVKJ6nZ
jJYBBfDWJLE3qdy8KrO5Hi7WV+Ewnfe2IDHiqiMsmaaSrA4wCl+JO7IemLJSJbGf
e41pXm6Fn9ShuR5chiKZFjZ1lZC5HnMtDPxKf1jL1kBciPnCkegFp1tQSAkEZvAR
deOUgXdLjrleEoCpHjb3Kv6QnvB6Hz9NzWwYS3d2stnX2VgWG/hfK3Vr9WIsOMa0
GTcbrhlntsoPVCCnfI1fkfjPR0L1bB/ksoqhNRl8wjGAGc16rhtF18D/nNdx6H5V
2tGDRUDg2bUKLjIfWZ5EWEdM+cfHgAYwTi3uokC+Dnsc3NH3YUIAryuKLS2RmjZF
q3OuT9K3AeSHT976xjTFtUzB2E02GF6TNMNG0SrHRjgqY6Cl8PmETAmMaKuI4nSh
0nMu226Dvi3NxRYFymcnoiUv1hDMtvUMYRRuUh7bdM9DHBsuOREJBDpKrJgGOL48
IRM+XOXXrNF5b5oTLPJUR5mJQfonFl+evLs/gfohRbKrgZidmNgDiJBa6ba8JhfL
ToIzLV9Rk4Y4muzev2eSIyYN7CenToSkDCLrXZzJSa1XAcuiDIJdDeEcFepKYBMv
zhvbxB1xdOtY9RhVBlnukXPuqvo2ybOd5Yp6YaZ5FlRQh29A0t/2WBcIgJjDq90b
erHCP+7VpvTkv5Rz+zyzODDiwUgDQrWttD22fMe0KlzsxgCvCIcJGh2EHkrbV/+m
tJGOthmgBD1AVAJV2/CPkbOLoPTFHTGT9zLdHQqtVhfNqt/tw2YQj9zcZ+Su4lZb
uCrNo/brG6U96eoX8s1OylIZA/ouhTMjrosYbEARWaqf1nW1+yTyu9ULQHPc2fKR
g8QF25rkFkO42+Y/6RYfhw7RmFl4NNtRllDjOX17qKpH32d1JZzl7zmxyEoyNl5O
MTjLFC+NAwfNbduUv6PYXijqSRLzAQ72pDGe2BlDgAxsJM0DyCzkZgr2u98BYzPr
jGvWdtF6wQSOQPSmuFKIQq8ty/yQB/buoTKpZiraiiFMucZhamZLg4zkaZN6YYVt
BZZ8wKmsOTVRJ292yY+Fwa5ATotO6rYv4bu5shKNQdGRgEevcbHhgLnhDPpjItoW
64Gaw9z4EFUdHw1K1mV/hi4QkSK3w1Sy+4jQ7yitrPLsSqeSmprJgTObhpYPxfvv
iEx1F7vuJvEgJy6JGvVHVlAW6xPPwFpKlC19b/uF48XzpWzgdwYEgz2WPIHDeV/l
aHALocIQCPJeJ4hjBIzoArFVblSYUY+LLeV684a2/oyxNX0gzsVJCKS2II8w5tZ4
codMkoaPBz0OpETtMziNJj91XTOkNwEMcra3BdeyCmYxJdS9yPcHmSiTBlnNzxmN
aO7Rqtp9du4QrxgDy1gWWsvSMizWOuRq0xJtwAZsnam8jgimUDdPaH2RtJHGxr5K
fDLr2CKYKDdmM0r83Z+Zww8kRPRZ4+83eAXRnF/yAZamwi3Wjsk6iQxpwfLuBwyR
mvkn7C6YesVMV8TIDOFoo7sZdgEcUf32Wh3Sjjh9969ROxgtk2ZenQ9fDYObEo/Z
4ZSsEorOOgmuCwwJJfz85IOtsI7RxUIz1gqfbYZ69pmHdulzaJANWyVdr2QCWIT5
WDbyR/AgAzAHtjNv48CWtTZOQfNcXG5WebX7yXl1admGbM2mj2GTRtvvqoOt4gOm
214JPs5tLXKGc92iwQwwknDkSBc2g/L+3Fl/rKcTwdg+2lkUhEQqJnJURLtZyK0H
T5gBCOlmCCTNQT7hZ05lcseFrlXNrJcDtsPVbIorfrH+kgN78Mqokh1kCPx5jzY+
I9uhuE8TUMWEiMcKAbiQGTrXX3lUDmMfmHSqTGWujovCB3dljbmQ0ep4sLaUpt9N
Y4rdibOdrmLAqC4hFbsqyYSTzHwLsuSy2z4KjmAKFbmtxuZu5utnBrZ3CZ15Atg6
t9mvq6If2oQucx3CsGJP6Gg2vNaBkIp8fBcuHQ8MZwSND/lru8QlbBLLEddFyqyj
/vvWt6J7/dAzGSVO59LSA/MTvI7BkYTT6TeyRlofac6c/ZCcRB5DFal559dSLaiH
q4o0CDg0wz0D1JHI0fldW5oiLUKsvc1WIR0NVlXKIfyqITIZnF3Md1KYlIuKJxTd
D81h8aYxKAl6WvNYsFFV+9lBikbeDgsz8mV/Nb1ivQw4u4Zlg9XzL+k4Y9pGEhv0
3otDMC5CWPZAWiaFevh7b9cg+W8jftX/dus4qyV3VFz3Rbcqm534dwCTGamOPuCY
VvrO0x+Lp/LG65x2T0v5iyKEMRFonEQHI+CaX5ibhwFTvgfprG74D7c9BmS1iYmX
FKiGGvVVccujdI+nw98TWcQXkQB58+vxUrdlFf1+KCd+fRomYhx+GAEJpIWM2Sh9
uS/mOhwgptr75kwzUbXZJdH/IIAOlx1xGfXtzoDNwmUrdO8Bo9w3mZ8wxfz5run5
9fSbhbQsFwODbCISusPqQGkZX0yfejLvwBVbtrzaiEDVsdy8mr1v8XeHNNsHypks
lcocKJyP7wNVFGeMEoDpBw8KGIOGkqK3skTqubB9o1wdszfCDxUBSTvTjaZGr0Hw
q8gdjVJ7LYxoItGSAiQXuQm0/dQ6eyBXCEZPZfxJHnFkqIBycHQiIWTkOL/ytyhP
VrYqMdZuK6yVXJKqjmnGe0cWeAo8YAqLFc5cn3Zed7pLAg+hkqC9786rxu0JQzhX
4yDYq4eGEU6OQwN84cylBVpcpKYNTznCJ7ajNbMk4EKBEy4lUYxr3blwpS9MX3RP
jqxD8Xmu4HQMwHrBQLAEpTuLGXq0CQE1AfGADql9YuKke9Hd4Q6CTxkz/hrLkPkP
mO2KT4akW3vEguRT3y49V3YN9CyVzOUsSHphcoOq1FTfBTZguyG1FLTTsxJZvmrE
uUShjJ06KF0CfHo8SgJRHskMeUO+Y3feMgd/a1223Uv3EC87a+rnI3RKgzOYHXzn
vi/ROfPjJuacuXiaVAuWlpAg5aYOuWWsyza2gtkyYJ2j5Wmf9kGP5zFbjNRcE7hK
PbX7JAZLaVCEDhzdm6wjbjmKK7Fe5QSkeQZ5KubtEx0DwxLTH48yzesAsx57bE2l
3HD5tzWoR+Y12DUqzHbrl7e2mg2ePwxzgcGSUOZwAqy4DU3aBOqHubI3Io3tOV+K
+/gi+u6R/TUJUoUaLdm793BUBY6eopOQ5fLLWkCGSIVG17ZAnpkq5CiLZ1wU5Tue
yG3vm2ne/VzJZQExMg8Umn/yzWiG5TS2hYifvUdSnqlzL48DHaERGMAeGZOpJ+eM
UDN1Pa7iRgOZ+rS4ElXy5SLTTIuyah7PGEWjQ7LoRIO1ePNs0eun/nNQYA2cTV9x
p0d4jU2lk8NHAn6QSuXqHeMHTNpoqBhWOS9eiJQz6186l0it63Q4v/jgWqflxJak
Ksj6H9E9jMeaq7vfoWiyvZil8QNtIKyHobdpijvbqzBXwNlo5psk4cCQv8melTEy
jh1VUjsuXLk23HW44AD3Q711AujJJnTMLJFkp0/deFJgTVnkV5srQAiEm3veeW+m
RDp5OwG/+OhZgD5IMscY03oB8nXLRsfBXJUMN8ioXaNKPVfufPrZlgWxwbRCncMF
u4tuvDDXS0Qua7pja0Ls0HF/rqIx7Z5TjO3tS16I0z/z9qK+rLzikTJ8kb3aBF8r
e2J2AYiNWrA3o6x0iSn7ZDz6kBb908TCd2nqicFLG1ISGUkllf92HtYSgQ3drdrb
jknsueClf8+WRQpAymNG+WDN/XkZAWt+Ov8YM8rudmm7uYLb0GkW2Wg/URXqJqvC
8SC0YwBSwjgJP66fLOrehKNQ2wbReGp26AztaT2Y4JxYcZ9uRvVktPZrf6SUp8Im
Zg5tyU7CJyuItHiU50AUGkYy3x6ejb9gxHoOGR53eyEw1o/8/a8/6Ab1omqG47ep
2sDyqXHvphmRHrsZwX/TAoIIbVoaO9gxjEGBw/aVpxfAX9fBLxT/+1tI92iB/c+e
DuaulkoviDX9s6MfLa8laeKUcrJ469CMRW6lDBMBvJJXAt+2885wlVuwvAyRt/Kv
ToKEuHnUR8efHe1Z2xevNHrsukTA8R2PsGOfCuFCKGos3DP/4YnH5rnD3MDTVdVX
gWzM5lX/91wz2t4SW0DF3YI7MfMYh7HCKgI8dnuXkR+Bz1MVoxRpMJlxPE7Pi7DH
3T6TBwVTsOzGUwh9UVzs5hkEGZhn+zGE2CkrKMF3TzpvMfaDKqUJAfUgeQ+5njhT
bTxoS+pC8KH15ijuo73NkwpQb42jdHIkSPugVyQthMQh33EqLotBKkxUMqOV1BI6
TEv7aa8Yu2gI8NZjyumZrPQgR5PteGzHWPWKBBYTGQTPY95D+zo+fSNIWMbvJ7q2
9Nlwl9F8/8boeMfwhKlUHBPmsyJriZ4NknSHP0QsP138Mrh7PcVXcXIx694xOJlD
r3cH7rh3rGp/ndvJ9rDQB9kMPNO4LcguNJ1rf7c9CAqTC6XPjcgUpSZgMdPISbIr
5p9TV5jG6qBKQ61oTXaF7uHZL0qVdlRzGg6tLwsyQhh9dxvOourveNwwOnNOohed
KDTRcBzxEv5+Iz3JYhWo/gxe4zxMq4vxYxWUdwnpjXKVuCdNIplFmJ/xVjNNWx7I
nvH5ShyurW6hRcgvmnJhwcrXu1CAeTz7AVn1/dN4LZTBQ1jt6h/b1meyiniiFcs+
HLOAdSYomCzUWE/T74JFuM2jzVnjC5HW7A7Fa/6qziA5EwsKC/Dzfer4VfKLsptr
JiA+Zf+5NEvH/3LkiVeABML3xoykS29op7WOWjoG9qDLaU0boWtkGH1KCHb9+Fwf
xddtz393P4mWFj5+LWArzc4O1o1ehyMx9EsEP1iaoHDFD9F0JkWYB9qt47CTD3N4
L0MO6AQUNRx0vSdvZegIECxDkkPT88yXj/cmvzoYCZFfdDiD1G+8Nh4TMxfctKC2
faAVvpKyaoROyvmjLiHMXU8jwcP/xaEX2UvGlePuSy1x1nRXQgJvM6W2SH83H6e0
Hz8S1D+z3iXZIIuNimOFcGjozXAQ1o4InfARjfElwuPHSn+yOK8AKZhWkMHaNBAU
nYr2zVgosAWlg0Z9oBhMGose8HEeGq6A11t1CvlujDdmUidmFiDx8HK3SON7fsvf
Gr94TjQUmYOYcetWGF94+KgxT9TlgpwO3VwyYLdQ/Alvp1ChQLTaD/CgPeIiT+tQ
ZaSX8zJZu7Umf2SwwE7qut6m/UxNOuMYPxThj0wKEmP/0OuensirRtil2gP1XvrB
WLUDqtOE1rZSoXKsZ9EolkdOjMbCaMC5tPV2UbYbX/gr9wrl2j8pIQHrFWT8nqXU
LZDpOSWfMgsUGEq6pvmr3pwpOCWHeFwoJqOyXPMpnC/10no7/wJGo7DjcAB9cgyQ
lCzDnxWuDHAo8XZVITeklciJI0ui0q/OE71kZOaYhNrglKTNtqmfX5XiWeSW2cfQ
nQEdwLhNUcCR05ZY3D33inIG5sNO8VEqu/a4TDMxJKe+JUm2BTnjKydNbPPB4Q/3
n5OVoCuP96tRBAPsDCVmG+oZwSgfVUXLYpW6CG1CsTgm07OBZBCPdOhI/KJE60fK
ha2YkF0XWIv8LoCesa3UDKpeUbnPYjbiIhY5ANst+0o+FrL6JsJ6vOraKEt0+fPX
Wg8Z2PHFhLuuZ1bA0lq1rOGCoQWc0AayEbFqP9XCWDxKnEWS6dz8rCQypeztZjwt
sgm64GBlPqtAurXn3kb4MaOlmfufWyr+dBxm9niyHPdYhsN0BoRd21LGlfm+wg3M
jCCeNh1MHHDOFHhzFkqmB941uOvq+Pn3Gva9cext+VQ0Cyi8SGTsYVG/LEHLsFBT
bnCkuc9FJOc4UhjU0oO5H+To9dopuWp8JqujfVjztKM2rLAbYw9wTXeqijWDLY92
wZR3UZQqDDQlRzQAP0DQNB88LVxIydccom2y7C2Xl595fRP/i6nfKYavmZ0m04G1
MOFmgbfgfPkz2vgGxzHzM7FlXwcZFe4uwPoNKm9tch9s3h2rl7cfClE6HcYKogaQ
xOA1qAIOoWu8IvQx2X2OlCTL4F0lBl7aj3u63+vOeylt0WJ6TcM3zVdAgiZhVUwh
E9Vl1KPM7/07Z/nwH0VkdNlne347qGjLRViNUy3Qm1ZRElng3GhJn9h8Ou8Es3ET
nVqP/2JjHsTWlWDTQUMuy1RlZpfpqdFb+QFv1Uv0loUcWLMDI1LFr92w6gvaN/bZ
5+ko0R12lJxuyq5Nnw0TqDdtQrJrjMGV72IvvVsfLpRbUFGcP4AvcB8SLo9z90mY
ccmUxB6Tre7C/Ghbvnpdl0g8kbTmFXAVtg3iMUocoA+mLBd0Do4AHTCYyfi4fhEq
cfalBhzZCJCTEpBCm3gnWJupZBlbJrWeQq16m8CYJNmGB/V1iITGZVuMpcJrcd0K
hxm+r8PZWM6cdQco7HWBAZdB5r8AbjF5ak0ok8b+1YkyH4/SmX08Cn9vv3kRMZNj
drEPqRI/zcM8qZjmtMsn2TKBEDBG26yIP9r/iHbZ4EgjzJQESdjylHbcNw20jhrY
6nvetAgTPC2sQKUqIhP0+vTk76FNGzPj01siO/8ZlMZbxxiuE/fuZ2ZMX6LTiTnU
QogkO9+8MBBGCZJuU6ltjT3LEyHRxNgzzGyesh2VDsLoD2lnbFpqRcdzEp9v2I8Q
Xl98UhAKGcGrO8zlH42k+jF8In7lQPMvg2glDVBRgZhUsinJtRv1KsMG+KU+AbEl
7b6F1JVvZb1t+jHa1ktJR/VA/LUME7xZihjpZe0cWmk+fNM4G9s25NSXAfZpT5vR
U1StkNjMF+HG4AtuklEQeKXCaS/1SMOCEgCLDgQqnTx79K4e4jlQe9l3RtTNedt3
U1v8YRrgwPTnn217yM0ItQ==
`pragma protect end_protected
