// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2ZlX/flhQk0MUcPdy+eN8Xh5gHUuLYSNfOzINjzEK2Ppe03xNxaXFNaqmGb412ny
mD9FHUyPw/1NW1vRSEN4lXIVcj/CeSuZFpJ7Js/fp/AlirPy/67DHb+Z2t0FgRmN
GUMYbuJdGdUOe7ErE8dBVLUoy/C2JGQ0imCNDPhgVL9nmM/yKyWjqQ==
//pragma protect end_key_block
//pragma protect digest_block
Yfbgna2pBPf1+mBOJj9qLP9vfj0=
//pragma protect end_digest_block
//pragma protect data_block
JYg/aSVUOUnvskoHbEzsdJ31IilNu+c7/fL72ml/ioQir1xBpk82KOlyTVaAlh3J
K7SgrLUO+wm19FgxTU6r4U2l1gqUtRzk+l6x2UV9Vehqv8t/E8zyyQU4wB0ZJ0FN
chsGOcJDWh3AvQMWdukwLJTD12G+OY7OhiZ/BJpfdEH9KqhdUqE171COr7DHDbHq
y6OrHBAkuGGcryChoGfdBlctJLU5W3xN5UVkMTXok3cv/DqV6jG9wm4eCB8C/hcQ
qB1MRq8civsZh0aXCxTiQJ/89MlG15K/nfXgYDduUgvc11nmCpADnMejIdCULJ9B
lSwygIFfecuw0HAfPUeKiApLBzYU+k+isbZh5511kLpTTA5+cF5abJaU/atvehOT
A9OXtb9BDOcyzL/MWG42eG3PlkIm9fUkfQFgT7lMplshPvBqHFgRgbQvolvUx5fD
2TXiOY28uC9+FOs98tPNLgknBZ4Mo9TbHVTiW9TjC8XMZgv26WncTHOX0h5eSJu0
RIKlSxnDMmdaoVKbdS0ipUZeLmUdTl5gQPDTDWgz3KIXxQJkN6fiuqp8MBBYEUQd
YXj+8/ZjcgTCtDBLLF6bv875TsoszUlAOXWbibm54+UK8khubOk31f3TdDYFFwXI
hjoxrv/4RVCzKbZUZxtOs9TaTHAL+NR9cG0RCy1oMeveZHxaza3MxE8bGRuyzZof
ZDlWHX6d0eqez0dwtVfnxbawDKTyTDbqRXS93qAmLNvPzmrDxcPr/pAbNLXVmI+r
k9jbK81URqnBoJ542PjeBJndH80fFS2rx/kr3GhjJPuZomuLXCowITnvWpUCyiwS
0UlE/uY7ItlI/A4PAlGLXyWu1TnvfEkjV6RRXvmV9gN+KBgIJP2hnkyf8q5dk8Fr
xJDLknXG/R89doHsp9rnPWU+jJYpjoh3gEZsADGJyl46BS823ZppBQLwpU65p2Um
NmXP1+2HObEEnTqr90QsgmTBnCOaymeiX1le0MQ6WOSrbMR8XELF2hai5dYu0RVQ
2t28O6MZ34KI4/1gYDVldCQyBjp+0aRUh/4P4z2J3mQISE6HN2rypflFXmohayiC
xbVojbR6dbompeZ7En8dR+2fXEiiH+LhbSXNxM+3WXgqQgtJuIYatmvetrF2ZAWa
IXmVuQP9zgKj8RR2PKb0C1kd9uS1OW4+Kwxrbseg1KhigayE/oZ9u/GY13INoJ0+
VBSsF7cj17xKYAWdpsMgy8SAHNAkJxp5yxi20dlok97uORu8AlJ1ksHP1vbdcg4Z
7OJZovitB9AKCudd0RIasRz1wjdFhzd25yQPFVTmR3blxwN44d4+flRKh1uugwPg
YK8WyhUy6VAgjA8FMvaqK10fPNhjmOl996V7jkUBq6vNJuO5Mnz29rYJkBSLLuvY
NjNwJRt8/53vkBWWpAOp+qcVVtLBfiHsXbQuaFIWitsJUmxTvFEAcxIO6NWqRO7v
tKfhHb5pxihYYzQn4v+RDTkB0rLuVTXv3NXqs2ZESqqv2o1D8EDueWg4etlp3ymd
A3A9MCqz5TOuLwHwyQZIznVmWIEGEHky/CCREyMAQMrHl/18wxVDZkt40aK9ywF6
Mc1xTG6wFoi4kIEgyIGo2uCM3HxsLQ6+NonDEWiCDa6gvMABjFMjj5diaGJ1Lex7
iPlbn2dcvFTqGGNRCKtGtrz4GF2Hs8FOEtKKVlej3U/7mYOptD0apocSSNF8Yy5w
lboJAHuSMCDpzI03i4Ts8/GiFXLybEUv262ziThDO1rmw/Yq8daQzJ7vVyLnJkAd
AEf8B0cGpYESC/LFy6sm5Hbp3NLnS7CXYdn1IDgk9mPYcE2rkRm74M+PxuhVJp8y
80J3kxPgMRyZF8hJdiijwhC0tTqxGXNYZDZ9Saqa5jwY4n783IsBgVnhRSVQ49Gg
+WVyvdNTmRb1mHqQnwGz6Yg7uT1c/zIFGP8GCWvuHPbuS3rGRXfUtlH0qC7XYiox
CPU2520kAvaHBXyJPBYm+DknkEje4KLP6PLHfYtdOVDrBJwQqx4U/YvosFUYVr6v
CUL+g2/IXw2fscFeiThp0YWG3rkQWud5ds5S8Zw5Tx3HH15jqsismRcICkv18Db8
jaqBZnmAvfLQF3TqiDTcC1ih91rRtsQ7MMmpiOJiynhmu6wRVuWeNggHRbDDO8fQ
BRUI5D1lAitnYAyF2uM+mDzF8dFJfKQovMNT0Ff2zk0mLxsvJv9Qhlz8aA9+RmNp
DB5WNVG8iBMcv20ho4ewZI5IN3uziJo0286LaSbHwYH29hCwXUmBRiSonGYch2sA
uWQEUDFEIDglmZT2DOnioUexXuT4oHq3vxgI5ghZAom3hAsm/Ky7H+LC2Tn8Hpa1
rDOgzhaDi+QsioIHwLmM3vTWJjG/Ho/I3tRqvbUIKHNg5MEmSKtY3kAcPFmpaOQq
WPFqGraV9pVYzL6Usp/oVxM9ehwLz828nGfZIjjh0SrDri/7mHnQJWUbKEKkofO9
i2ScSaJ9bRIOkabEpMPc0VpSvPJ9pZxQBSJbvVqUuda9M/2yO7syq2xYNwMneOL+
H9Xzj4LJ8MAf/Nuhfu8mo6ZHZbTygiR7bJB15U5vpKvqEoYMZnOIZZE0nXZeGCPw
IcrQp1nWjm6hffWv6LpD5WyzgGzLGJ3s+S/sgBGO8qVYyjrWuALWNKdJ2Y5Lq1fc
6Pu0CxZj7khgrGzP3ydmcc+SlOtXz/rxPG7w811rZUQInoBUtOQbXW0U051i1k0c
vrxoDw72GTmLocsRUVFAhvns9AbrZ7s5EPplDXGqr+OOlcXRliLSyzln7MKBuBUr
TQwYxeDK14uuM2M/Dv3XrjOqw7//UOBRAc7CONzRNS1FspvF1ZWOYwPvA2HBAKeO
mxJI7vGd87Z/GEtZx8601E8q5a1kG+1xzH5/MKTqjZ7JYa9VIcm7seIBWKPMUs0c
eyPXdLak5ZwABJZUdeVkDJzCP6o9y0tb30O6aYzTPIY23Y+13pdOIhHXup7uXKKP
mxmU++tMFu1VaRRi7ck3w831N07YKE/G5nqyZLRIB8IaJWX3TZ9xHxl2xQ5Dsco1
Fligcz+5CS863a+LbjOLwX4kKXTuc6QWStiw3N+TG7C1GUQ4zWNsstLL6EuAIPBp
YHKUs9vtTWl5DmpuJ0+P1pZ9IzCOHEKdFBGrftGKbm1bk3DrzgpWvWezHVEg9n2J
AaRrqof2kuYSwqkisW8w5QLxWz1pLv6rjR29aFWSPbp98Tb+8UrPLlbJ1nhoNeIv
K54qzEyrCLeelIjE3gV0XV8M7rFqZTo0Vv7wbYWPofXmGVmngnRbV2qUb7FMeAKL
QVGLtYJawUHfXnwftpCnNqyzlUSeEJXw+wOe6Tuv2DW27mU2C9RPK7ZgQ9sNM0Su
HtqaGRXRtmIDw3XuhFlBUbznpBT5AnUeSybhlyab0fu/VcIUQNRDBEqIjV/54/lI
UrQtJYKA8AIhFEYMBBF0OupQnGMCOXBPSINX4NKkCzpE7mliFhdFweeCVK6LbsKv
+JzvllrSC/rQpkBxaIPUlTnq1Y/XQVYAwxBdXc5kioTgXXnMOcQD3NQHq7lZVaBG
oTgFjUfTg3KAgtypcx6+Yg10TyX9fQ1xrZVIvp2i/MsF7kSgo0NKiuH07Jyy8nx8
PnNh60ICrM3s7v7rJrtHkQ2+IHMz8Fryv0pUxR21ufSrVgQmJ7VKgSLKHeP0nprO
qtO3rzPo1WZ/UNk/deuc4lY8pt6ctyIQNpWXu0PYoGPIdXA0lskOpKYqsMmUWY0o
e8ZsF2o7LnTx5Sw0gm/g6/19NWNGMX9aNuq3HcnhQMPenc57X/cre9NfsUgcgIMi
9eerJkThpUVY9tW62ixgRFvg3CFD79yTmz/Ntad0zI+ijkbkFoGn459qiVN/k1TZ
S1ofi5wX7tK4feO5aBBzdDzTCdl+mPWi8LYjeJ3KORlIC+qDBi+1mT4UqJKAp2+A
NyFXMF/nSD70l53keKH6dkbbsHO9MWdxVcW/s7DomQpLcKD1eIzX41r0uuMaXfFa
z1O/H3EggeRQACo8K5s2LWSMPMfCYv0mA+wSFhzyifWzPCc2Qked3VNU6XqoY20+
OgbQ+48p043oZSUyyCDhwCBdzKGqzjrS/PKYZjLbTP3zAc7dxTrCeytDsDQ/D2V/
Six0Hu6iYwOUAf+ccJH0WdqGHnF14C+ci+mK1Z+l90JonlKBi/rK5QIrtP2fPfhe
sEgDG+bfLpTT2bYQcg7OnkpGBky3HusW/6d1M3TuD7YdE+tHEmsAF0zwG9uIrjWc
ofCU++npWjum4TV+VATVmwpWwjQEFa7g4ZiXJFpLhCtCF7RMFltWittzmoajGJCb
7MO3802VVRJub1MRwM1lb0VCahrGCrMT8i5ulqyF3PBQ+3FXBc694duA/qBIoroN
3SLnG/SY+t5PyF7iOVmR6xd3LmrFgK+Fgh6zMWlt10Uu7qIZGc+yGBjeG64fRhqK
ZJ6Zi7wjO3t8pnp7vxpTV+Tgmsj1zDXfP6VN5DbuA7jUeVNIZaEYBTzfoPAphCrj
C+EJS3tOESHV/3ra8+PQZviBDrhe9Ps3ub3+C6gpeebllEKnUiLFFhRDTIaHsYPs
sa1axID2UfNs2irFa7IM8yiz8LJq0s2osc70l/1BgU/qdueIJbsz/Q+7WDXzIKHZ
zLJRb5msK/F1YbPn+snDcD3jvtZ44IhKpQszAJg44IdOcx/LLSYRS+BqYkttl8dk
ahJvPRKUu9IZtaZVZJRi/RLareOtFg+lNkKHri/tigMmEF1ceRQZ2uA//T3LZ2PH
oPq9u5OvEN9WE2Bp5IGVTWwrBcoCi0Uvpp/nSRQFtqGNS5lEVLFAZ0pHJZIfL5MQ
s9pfIJn7AT3AmbcgVOgJnZlc5tMuDvbTfN7iLcVkMFr46hVFHFsr+I/gRwiVjttK
OY2sF81ulBljpxDFPIPfyWtdbLKnyQyTT5z6hftPCFBbY/sp/c8WvIjV8P0Qw9wX
29pIxHO9L+l5AbxouJ+W6rwyYTZkOS0acq9tW70NaY39cJrae6BTvotwht2/RcCE
kKBl1rC3+J+xD2f4WBaQrNBuAP8Mm8w9f2ikGEoh9kr2hDwyUfEpPjmsNvIldKL8
tdgMsKLB6vNmJAcTMotmNXhV40nuosuK/Npw9GGovClToRsAeTbNhPH+D39EZA+S
f2/H4VMhnyQ5mf3/tUVTyQqNnsD5Y8sOMPtuZC2iRwam4VlUR1OceBxtgvRpdXkA
Yqdbi6e4CPNdNzqDXE9QvdiOP2F/yF40Evb9OIZnHfuf6u4JnA0T+3B+p3O8ngFp
sTOXuaTXgENfD6cZE5mHPTcmUI8h2nltYW/DuKjDanZu9b80cWndBvWo0vO71a8z
SfFihgUIeuvlKQC5dQMztGzL13/+5dpJrZQTkMabcL29uUsrRFSxaobTqMwYCIE9
F0vQUeTlbY0E3sOHwZ25CP4j9fumB+x6YjlYCo6eNbjdq2Lq1R5NvcMX250z+cxe
UdjcjSk2kmv+2Zo+6MEhldxMCb7BFCHyha4IQEr7xXxy/qEfUuIy9kyjD3cYXKGX
yG16zuLasPojJqsKU/ptFYJund45ziQp8ow4XnOiFQRjiXQZ0nP5VqUohW01B11D
Rc+TVs4vA/0KhKNEvUQK3DyaIQ4vvioc+yAgYTUa9ETAjs3eBHItJxUpblghG6LH
JgSmqgdnBGOl3jwqQQ+CTDIeNFelTDvrzM33lJ2dDxq8SFdIXX15eAstnUZ2Ty73
iPf8TAyZWFCAdrsEuRlXCOjyUeeEZDpToRAdyi9q7hlE2AXUltQyW9J2pG1WEF5G
ldm48a9obnIKR8ZUCewA00Ccp8usU87t5hYWK0KTwlT5vOfHn5MnNszUopoL6Gi5
Bohkw+Q2cDfyMBuO0kb1JgsnDnuUTTPTLLXonAkOIWDMYANaE4TthaV8hFoHkL++
sGB1uuD1vb4FYs3G2WF693nGMwzTLRCRIlkvq6UrDWSftVlFaMwbZR5pxc4ydhCS
lP3DG6W5yYBUy9SMOPm+KX/1R4abq/+wrJb4cy4fVsiEFQyjl36RYuSE8F0BMa4a
hWhR9S+O7aSaa3DomRtSuw8WOS8App+vXxQNVXaBP7UnWF06xrgqGp/yeqJUu22k
wTYgv243Cb9KehsVVSLZvfF7Brqlpj7xu3jUduzsvzAhNZPp0JFD/Wc7a4GhIj3/
qBsDkX61Fey+m1LKSvFW5BoPLC+4BiDQ/9e8yKk1Dyus8kp19MnXs2XeqaT1hR6t
EQUx6/2FF4p5q5QjkeTTnx+XXXx88eBBBbL9M3z4lkOASku8oPp96EFkcUkwhC1v
5+k+b00WXJvaim+Nnh63VOX1SXgmA8zYHlBRzbXjFVueU5AuOxyXhvtxjandyXoj
h/RbPiyuU0PQpolgFHc96VHxF+sjA4dNispM+7Ibi0W1r7RzvWYnnD2EmrWNJSgC
QZtmWFBM9AO0wCeT/NxEs0NduCC8gMMRLj3kqIWJv9h9B7Cc/Loo9sVAJcg76AUq
9sue51h8pBUSN9ELW7T3C/eQ25m3S3rKw8teMk+V4LqDQui8TFymcXiPc4GEY/cB
7Zbp6VbtRUnrMiatda5zwZ8x6D/v/Bt4bFuhnTAyI0Ppi+8sXqu6jEOrDUNb5qJZ
NEYZ503asLKBaXhVnKIsR4/zdZDd6XtHXD7ubHBBQfSYnqHPmYi68jBkfslo4KW2
AV1DfQQYdW3JKNL0nN+cT1/0g5wAdHd7USefcHF0gJ6G+fUYUUNwWU/mL0k5Ho0q
nzI3iFBAh7hwR1+QCsXMRcMqqDdK9FcyKdAznqdXFg3G/B2ums5SUrdQ5/hKTM/9
FY92hdjwGMBPTaoGjCSgXWOVTrOXZo3EmreT0dzHQ0NpEfvrbq0zpyrobFKUMWEU
gzC+5u4gsXbMDVCggLO9gAGcsjwstIjAutd+b5/MZOG5h2SPPOfqyQFE65x/+J+S
1XH8PO1QcOgfzVAB+asLy4mGOxVEzzGcv2xrJQ76wqjmVEtGUe9z9phXuuDrvO3s
lOOUNNmVlMJmFGOoZ67KEMglWYhse1H0qaRih3qLqCDuQA9SCihoWdYFAxkurNFu
jlcmGM2nMFNLFEp5DZy+FtWEdZRscYcQD+Mkm7e9+71OeX8B4ktSjDmH3pIOhfMF
desb5+zNMxZqg4kdTVL2CUIhv9UASvBb3M2QrRdoMviMn+i1ul0dWjjMpcgheHG5
VGqXVbN7HFUHLA+7NO+Y8ZuQ9Sc9aqFSsan6J5BUmzTVAPGGWJm4Nhm1d3o2gvsg
xlvWHr5YSfk1bkzVVBInGXMlqNFc4HTtC4e4xVTISaedWsSoXFo5EaQUcdh5W903
USPJpJGwbg/rtJV8guc1TvNqbzP3uC1UP86mPQMpsrRngMhumvzVZIEmeQPX8clD
Avyhhzet/YTB2RduyypdvPWR2ec/IhqKXZYONojjV9a9Kq1ZirtManAr3UgfMA6q
irG5I8nYnd1tLBkVj0U1+F0htTtHZR0ZNuhvjTArIYMELw3oaj3mVK6Z3Na0yRnC
L4hmqihrhXZb39RAh0BTQ62vDNR/CkvUzu9g0LEAzOq38kgj+EPh6ayU/duc3U/N
V9mRL74e9J0yVjFLd35UgOUmNw92aelT10OXgvuDJ4uie0a0+W/tZLS1a8OomjIN
v+P723M6grqNBuF392jODivjGjiY1uGLoy0sGBiZdGLv/9hmhhBMLOTcYe+9SdD9
YgwUghPJvFYA0BiTtNaMAFxR97jqndVC05Au7wM1iTA+FJfiSpGgWaoETZQmZmL7
YRIzncmMdCyWH+E3ZHFwZAwz3oc1MgcNNPdrJLHt8QwzItUeFrU5DVBNakQ0hwWc
Twrd5m61PNeQ9uyfSxR7Ujl/LpqOnsLgslPXeJUKTy96lpk1gXoGqQmPEU+f3j1S
u2l+ckmaoW5wETNU0UxXxIE2VSsXu7QrX3DoVVGOdYcGQevq7TjSW+3dSsRTT+Kp
VW6uJxpoIADtqQDk+OQiYH1zfvkmANnKqZM+XC2v7t50fycoIhc9dklOUabxLkVH
YExCcEqoAPJUxlefFVNBcTjZdCb0t1e1/k5ZHcvNesllgr4kb+ft+lEhzXsDwyB1
uecWcV+KZlo62Jq11Xb45JT0EazCn5Kaf405WlVW8oXswl/S9IGo9t9lgATnOtSK
3hu0+MLN5dt69UwTZzOkwei+HMm5uPYoE9sWMgZw/2A+FHvqnYOS4xSuZg3j12xc
XJhxANfb90vWTMslQ9WN0oU/j6/JoRbrmL/0FGazcnBWN5iBNz8uwPLPEmnq2iE9
ufU1vRYxQtFE+LnC3BsdrdKIugFnkuNSp7rCxpTFS7bTMd87L+d/n+WJMtVgymDw
ZBmJCIu6nEwfGYg8PDdaaeq8DWsgjmvwBXI3/mbHZTG5KbDCr4l16UxTmL9aMY/u
3BbFUXYc/8Ywdw8kH2a0sBqqu+wmNoFVOZvo0rAWPq0tW/ucSburoqo4M8Sl8UV3
TyeR2HZSAGAxtT+4mlhuTg+J5YspqJuNxISy+sacR+xxUY5mBh1AO+W8X+lPUtKc
Iitsm6yVdwUhG4nDv5+X47hCD0e0PaJWkBxNFCkCB15XTC8uF2y1tHabm/T6HSC/
WEpYiu/17Qhg9HjGkRHpH75JTLgwByE38aIDUF8fX9u66NcMoimFmaxlXEe8bJim
OcARMEXzKws9kxiEKdBL27baLHo1f6Wfx/rqj2XCx2x0wt7H1m6kDWRv1c95r7Iq
Oi5xBvfVzWDsv0O8D1bnNmAkYB1xNX12SJYoOzXCsSVYob6/96aF6fOVFfxOHClm
iOO5Bh1HvVveQYhdLoOYEs4A4usWngfk+oTQCotipFT00d/bHL8YWseToWLQxVP4
q102pDXmqVlIFstjo3mXisWvP+/KJ4QPb4uRA6qNCZBD+cZQO8Z7QC6IsVvFp+Am
s20stjFCOzL74kZ2Nesu2w7sebh0Tlic5xxl3TPzoTIQtnWWU1pVLKSJ1zj9UUN7
wZqoB51XEjVNS9rwgMtIooQfhdyhLL3rDmr/JKOhpy/1ZAOPRlCRNoZKxdF6mCna
9MECxMV7tk0wrm0hkaziAUogwuBTJEZgiOMwfsKFA9aHh+bJ4KwBh2f/r4WUtEuh
+2Q8IJvadScSOt6TG7A4GfuENtX+X9aEMAG6UWhPGIsWZPcDFzgQjx77losvF7y4
CR3D7T9E1/30YJJUbSWOGxee2N90PxLbjF24L9WypQncdEAYGT7mRt9cb5mGN4Nr
j8I1MYKUW8Gj40paPnM/Uev9eFLZorFaycS5IRqrYkLnaQh8R+pVIPqp++emZ1Yn
ddCewT551DolIQcjmyTjVDkRCGbpNC/Zahs2ExjoStx8kHEfxyFjmjoyuiBec7So
GPFtfmnZri2hfsPISRpoZMGNpAtrwtVHywXe4bh4NyKQ4zCNnOMkzlbVPeJZnurq
uLodTc3rA3+JMpT7RRoDy6WRYAR6LIkmT+6flzRY98b/3pECdEFiHtQZztgxLjC8
6CnznskUGyzbfjc+oCtTKJcOaCEeuuNF/L0IXu2u4yvQ+eycd43SyER47fXjOqIU
68E47qI0kVML7NeonmJIcZ88FFgmoUh6xbSqG7bOoMcXalBDu75HEAUaPQgpGJrt
EYTJKmSPKGK9ixJoizmzCuMN5tocTC3vxmuF5utKsivGlzeP+XVlyrxFdvnBQEl4
gB+zDxckQNN88aCZbe7v9bbRMn7hCdATph5KvyYJwrOgrEQWAducBHAG4PcbOhGx
Qbc1X/dHwcreTrIffskaj8CgRdbjOxhmgrz11bV9C2TTmxWGdx1kLQokKWL8zJ1a
7hWiG9HBxND27MLdnKQHH9zYLVakLzH2N/c5b+W5Q+DwH6HyF9VcDYxJqS/FAOJG
Ork4/Kj0nXllpbNlWe1bQo2dYXAtFpEGgl69qaI9CyzO28mV/dT3X5P7tbR/HkJq
QD7olKz4rsyTFm4l6UNTj9PK5y/OpY4mm1h0VlgHysg/IGlGFe5vX1o0dwZ3oJYK
0KthLxNpK+SsxXdAflwbV9jOG8xaua9lDTle9+5jeD35EVU8AcnnmjTz5LVetFzm
pEdjFXsH+5aiK6AQHKF8SDK0vmcCsTJmExCzOTjm5ronKpZUcAJPdp5swLGpOlzL
TUV7MKzC4yhuTi3apLV+6F3ZCycKbai0YXm0pydbeZFhLWbkCMI8KuqlNzZ6r/5/
9/jdAEu1jM8sSFlx8fGH8S94GtEK6MShA++20YeGtkq0Wr/QG7dzxneHAHrtwTQW
NJKUv2C/v97F69D4lGRA9gULWF/vDdiRFFT0a0yQ+A+Thh7wjIwSMGlCwtIg8b6I
sGwzAilUIXpo++AeNYsNY+Y+SXvXxeZOVquxj9EWMJY76vTSKBJcnMHBw5qvy1Ze
bOZmN/FCJGSEiaxNxPkd1RkGy8MdtRfv7JiJdFxUO93GqMu/22+Oez4ib75aFIMj
tjhGXVlcKEDRiLkXP/MDtbtb3k/zIcu2hF+OtNmnegrx5CP3VBg5QPjvqOhxSWIj
kowFt+PQUZWYay7Ivj16LthXNQhV8A8kLtk0UljOswWj/4zNScd2SWstZe3umhQS
9aOZ/gzh5pJ3X3MGLJK41QzbpQp0LW+n5CShpVapVAY9FC482gKYDSQqKN0xMWKZ
sY3tfbGvZnfQ5OtR/wAM7PizoeSnI9HPhPhJNVYwxIl1xU77isPK/A1vnY8t/ldh
GsMV15P/894PH/yE5CdPAHfPvTellrCYe5+JlFP6QHF7TAGawQ0PMyoft/AJGQ3K
IwOrm399RR3Ni1fPm2cenp5sNmACfVRtR2BEmEvWRJ+NF1tkrXsm2zCEumHy+2BK
OIS7zbwN43Asg+UQ+/CQrN97/tOHFPn1t7O2vsmi2gQcJH3vTkcr9G38sV58BFSE
MkRePqocTK9YSNCxPPJg8LWUe4Lahfyg4n/ifgwN6adSSgWz0AV+pgbY9G6wMzKY
gMgYmVX2Tph77cUeNH/yijtYMEPfbBHHC52AiF7S0Hwqdm+iqraxj0YRyyBYiMPh
VSb0JRlIyPxoVHQ69d/9tLgl3XdkCIKhfbDWZOhi1BW7TL5SfiytN1UbBwf4ZhT3
f/rPpBsRg9YZv4ZLjA60bDOR8bEIU+Bvw1mXS41XR2hRRXa6PKmP8xV7ij6DkijN
QwJhnXkb2tVXVbOi0T5DESDwX2/8GmofR/mb6RHtsDiPPXhpTV8ImnBISR6T20F1
UAYhjrbJMk3MXIWvpDg3uTbb3549hs58PvbF52wE3WW9axkylAkrJg+8/Sw5ijjm
eLbwOr6ECI9sohN/OEUSQl+SQNMgew25R6c/gcuAdzLEnf8fR1+hixoolXX/XnxA
9GGYvHJ5ne8s1x3cnM2n9u3UCiFpTOx0j+HwXfcJxqHLdORp3vdPkhNEz6A2dM+Y
0YX9MmHMLocc3UngOIqktkPnoNLQzDz43tkGwdTlcR7zlG3UcjelWV3vRoxoNp7y
BGfztKgfF6bw9MstDUg7A/Djolf0XlBMrFNlYhwMhru4HPt4MWT4jJpm7ihQJJUW
3Xc4GgTHcRx8BwQL5he18rFT1hn4SnY8BFYV8xHygd7/poCeagLcCk/G24YV/7uA
cCEhgpKzZTwXjO0C+RkpPOBu7gJLflerQYRIWaHe0DU6saXPs8W+1qZu54vrL6mu
TzUj/IJJ6Fwq1miqUR5KWjf33Fckdx7WRvfRpYdAE4E2ZuPdw5JTv9o7crTtdVNa
cIyp06EhFUJPDotN3in+YdE6Ffzs/O9d/xryhN0Yz26Tz4PwpxL7fGAYtkH3zjTu
KQWFq2NcJIvNw4/vGrGxnOiXh9OmyvIZ+PyuyZDlQWki2T0HXPCW1N2h2dixBGdV
I2WfR72DLhRpnZAGYlCerio10BYNn/j+SrAOAcJoaSBrKwjVJmwUsKAkibMpRcKY
FMzz35ZxQUYa/1Lj+K1soViYAuHI9ezENNu3Q1+7U18uN8qExe02IMfQDf6UspKa
sGrA7AtLAuoLqZeqrwY/fGJKHG/tLG0A8iC7uyLH4tpGI/VN45Ib+etkqXVXVTqR
7FsBsUEamh2nQcBq0D/Q46bLxyw7ZAi7vYAir4rrESbCbH2ZVmjqkGvRqY4pZ2CH
0gLT9yqJrSGCHNJNedbiK9pynZrjawhYxwpGUCwftjBmY1d9Uv9Kmub1qCjA7snG
w15UTKeY9kRnfvkcvbNqsjGHtMKWwIMRxF1zQhCNbSfuQkyo9LVjwGMb5dfZ3ehf
SBRPq0amJC7uB35b1XT+K+Tz0hSisZ0MgpsVDA+q1uANxVG7vYXJyfFyBzJs2gm7
T6F1zy4DI//ydnf2b8vw1WNcGHs36ItYcsrSwzb9Z79TUsCbiKTVgJRlO9I+sBQr
vShiuu7J6vQRKyPEm6vjcy+wHu6CewgOyXi/uFHbdGsCNr7WJVlal2y2GS7x+FpC
DflnQCLcR1HrMDpvnpHvgIIGdsSAdmiKpkwKMaduL1DUCD65pryzGHCJEGPs0a2W
xpJ0L4a2a9n5/lK/6KTsdgm7Dz0ObD8AvW3PKwqCZAgtzC5xPDm8uqDY4xPUy2Kr
jhnT1vab94vQ04SbA091hp28oqm9PAW5ClbywGXh2cw3mRgYain5ZzGQgnzAlhPT
HRnKRpXfp5/sR3BNZVc96djlt5c4Yded/nHBUazza2vcWu/GKWePt9gM3/S6L/wa
lEoO/6aBcqDPu5RgpXCgIbxBiovqGXpHNFYKbIHrE3tpKimZjlSPjHKt6zGXgYJ1
JenzMOceRXkSnCGEIPAwtEqd6Ava9DpEdKB6YtnF0ktTYISJOqePw2FU5LGhnxeL
rsMdnRjge+i7LDV3MBgYFq2FDUcxe6jNIP0xvwNd/fqN7dvWaE4zdggu+2zucYNL
ZA1HtGY7SH8BuAgfOAIbeWIYrpFT19ncWOF2WBxy0OHyMlYHctFyZns9GZwCMT1Q
vRuzZHj85AWVbXLFOKWaB3zh28IVIcsm85T2zL9+CZ2O4ENt01WnkGS1eW3vCTaB
NvFJh7zTH17LqEtpt3vcQwjE9ksrKSYfJqN2M5uKfjf3ujO3mMXAEnkk/4ypQ7SC
Fho5sRmJ9613M9opt/vklOzZVrFrwyP0l1MmsO+QzyzQd6iglYMIxJiY3oBuKzoz
6+jueUKU3YzQHAHFSucnj0zjyi7xrFV546Z6SdKMrzQq81XVr9+ydj73qOQXoCeo
FHyUhB/bsYCfw/QDp63nxK2Y2yhFDiy5OsrG4WR5aO0IiTFs+twdgzTsSGJvD95N
AvEpW8nmI+R8j2ohjaCtpWC3Q0193UA2T0OOg2Dqwi7+tFnVxkxeZBEhwQNtUV54
4My248Vmy8Cvh6y9oqo/Q+gGuKhYhWVYfi5PPwUsj/RJJtwZ9lgl9WTJxaUid09J
/zr3fwplCGXoPI3ezZfKqHUHIeqtDiBRRqidkJzHcbUOpBGEMLguK2Gdab/1tqqI
9fmnD4L44wdehkUixCurU4eeHoPPja0Hz0wkRTSKlE4BuLLujzxMPz1dqWpMYAWA
nrdkz8vztICG1O7RtauPOqODGQfQoAATKW4WYeH2fTMOGYQFXxEXKBuiogRAZ2Xz
KyRbU6hZH4GHUScVphlOyEah//lgKOjJqQlSpCO4YiRA0KaYyE7cgwJU13ROmVZ1
tSl00zBiOAHYaelbosDJMzTUbly6C8pEk38y5iUDCatzdgQ51rcFn8zkeP900kJm
NiT3jLZo7HwOy5z6IIaOVGJYStCYRs3tw6AlWf5GnQJjmdqMH4mk9Rl6XgbKrRyA
OfsDmbr50eTKMPQo/6oTQdamHzrezuUI3o8Jh/lJKnUEEUKhwhDzQKC8RMSeNyjM
qHQBot/S7slY6vzo1Tk5j051SXb05YqIy49xwXzxWa1RaH2s8Bbj2riiv9DGwHeo
jDXO9GbRyH66rHCDI1ktSy+XUBiBBdL9k4JFkgSHXK3p3y4cwJqT0XKcfCoHsyAr
hxZyMtoKdXqy1UAIwGKPuoveYgM6285hFb1Xp0hebCTIAsNBo7kR1mZ3YUKq24ct
ntqJaipypEx5CXEs8Fklu1/5jHaisI7J7uRnD6Vy/3jCGeRQrpTz3BPkDdq8wD2d
N211IxEXRxbXNXfYacfV2vZuhHmbQyPKoY3GDHHfNDReiPjhvwEt+AZaomyAfp+R
/wuhjOGvstuieTvtJXhC2lDSYQwxzfjYii+GQY1fC29M0wLclXAxFWjK0iADLI1a
xOyn0DqdKr2Jncv5yhH8WxoRXJyMmOHGZghP3FSLd45PL+QTSpTMmUpcVtI4vrY+
aSw8+/nW08XBatVC7mTWa7YIKmVZie1LOVHZKSL9FGRB/TuohQfo22f5zwpxtlW2
yvgBp+nG0XmC+hqX8A4UhVTuz7uBBMwTy3UmjFZkmwf5ijbKVbgKzbcPBnFCjSA9
ay0UWsqT18zXD8BL5OOe+KoKOAmt4aRmWGgnOSzOVjAeh7p+BOmez/BDi9kZiZjo
AlqbW3CgPYlNwbrbCrRoc0NIV9DcqPwByOiDRZcBJkbmHAj62b3prp7BXqQnTfVn
Rsss6UPQyPrf7IexoAC42TT1Xht4w2RfPx2MLJ05zF8PooerVoh9Gbf1WtILZVDi
bIsmD5/EdJx0WNxGv89CYt1mk18NAhoCa2u46l/mg631ihS+dlMK+x4jPNjNUbgf
3SyIbBCqpXMBwbn+R1JEhAHxtPqeKacZx/D46ua/hztONu/fZQJN565JwdB04zKQ
KAu7bkWA0dIrgNBUYqEUy13LeI7qwM4LgP3++2TjXtAEL0OOLepRdZt9emDQ1k4q
gtcFoAri8GWqpWg938xXvZH7pbmmymjJBl5h0NIDeSEOmpT+v2D+DorvioEpd0Xy
m6BUGV8UM0+ZzwI+ogd8mNbdoN+HRzjtUIBWHpW5H10IxzF0whsojUKQ0qXjwjgT
CPuSsG4D0Uv/IAVBpiNyBBt6eLEKEgNBQvn3zyW2z1wu4fZ9TvrNP3k9bANOCdd6
Rm1jL6o9gA5i/+uIABKjWICciHGHHEGFk9Tqj9+ef6u0Lvn7rIchnc3QqHEB6DZD
PhkgE4xFVrmbhpINgNBWdecynRAf7100OZ7B+d2POz8I1d91QIhbP2FBuC9H9q5n
TzEZQquQ9RUzW1y6mkx1sCXFAv0Zkr6EaTQFVYiJyUJxr4etAVIZ1jsNRhQrED6j
8Clai4ZkkX2UPZDuXEpvf7kJcO5Kdas8mo0VbX2QOB/pS16EK0jmG/soGiznzBYt
MxevYfy/CZa8aoATBh/NSrzoxYTZiK278+l731Db08a3J1k8p8gySIdUYD6TKq1E
YNX0E6kYupuTlXOgUQYKV2wAPFs4Css3wUpXeWhb7h1I8BACPxwn0R86HwveMq5P
zbLThm9Ei5gARJISyTUsjVUew3Rz8xeMCmU65QQEP2VrvOV1/KdaLLpNOL5U2Hbf
gvSz1uSoPN5BlNPOdtBYEZ5mAKiAGtf35Fssr4gOvYkxy7kubLKrFY9gHNwtyZAD
qcdbAiEpPk9BOlVn8NKMIiDBftmQ2b9ozAzVLtAL6Z99pn5Ph9fqzGpTGDKyg9BF
J5gOuD7yvoN6bhv4v/DTSH2V/xuJ8nuX5ZbDTT79Hda0FcjHHm6wzewLPYMG9T9t
7Bgj71X4DxkwUYW7Sa/EBTBmW1yQcNl6/NX6rOkIGhWy8zbif75GOEtPvcewVdLa
BmvsttVAdp8yerdsAEFGgqCtUsrPstY2tPr3ZvrY6JRuXUBjFxIze4Qp43pXgakr
ce5ZDBt4wQO/I/g7MLo/rqDVzwsj+TVxVEqt2N/wrexgsZdFO7uIKhyVUQG+J6Mc
DW9umitLjGQ4AdavgZdMCwQfXDWzB4LNfdCUTMb+n6zVo4glROSd+oZ4XQZk7f5C
7EejsDP6K8FPDecdx/khWLT/Z/eKuUOvrGO1D6QXSkdAkVfQjgKVgorH+tPVGwuf
y0Ckv56Rtih9t56D3yijbpoKQF4yx14Wkzx13OQnPQYKDWH69T3nnVTVHKo2uJoZ
lrTxz5XqRvX6D+8PgYPqFXdO+3qfc4MDftbM+m12jf5mEAsaVUTDXZo+4r3TWFrR
4p9I9uNibjQk4VQPJZ815ttVVhOTROv9uhSXC5lmwwIO9hE4ctz/9jTGiuAUAAnC
5rpeXXFY/eb9cjI+myc8Y9wwlWmZbElVhMT6ubH1ur+gxxsTKD5lwuEgqKdYNn0R
Rl3D6T/HoRJrB7seaAyec2Zaxq2jIwVH3+15ILPtleRZF5H0zxiKdAshShrc0Oy9
bFRhHaRi58wOBAc/ryPVuhX7CZHcWNi3TP8brWhNtHnAxcs5Hx7DNq/1RJ7L0Nti
wByQlmBYF2y8MRmk/kjL5Jpl76uBNyDc5blR43i84envjvynr9KvtSUjUpvkSkio
skufWaXsVRZ98Xg2toglobxTgeZd6/PywEbcjEp7v2vMXQWRMVKNBa98tWgt6ZBq
EExmQJfotXiHvmnSzeM78rhVcp7q1cASWqArzJWGGqyrSlgLaPxJnUiyTCp1utSL
oEeXpXy30qsyIO838zAnxnhRyWJ/nyLS2zF7KzN7nTFb9N+vZr0SIYBpAbCrcDNk
0hkA+e5m95GDg1grkV0u7Ce4sJmWXkT+k6CsKCxGEfsxcO7CcF6vF/QCNsi2r4Oy
lmOf4jru6PGTuajYkxtC0v/Hnndycg/pzTa3nLSFTmDnPp2cAw+5qMdXOtANZEpU
Rm5jFt8LdSnX7poxr8esD3mH63vMmPmK6QWEQmnv4cd7QdQn8FuQ8+3hMZYNJ8t9
kkhJ8hUpoHhR7Ig302ME3Q6AQuRe4g/zvd+V4FW2Li2AcG1Ei8TUeSEfpNO19TfF
li97Iwg+lwRKvjEIznRNBG0NeMg6HcEChWbZ/4slJcjKOqSxCA8eJ0iwTWy+zivx
E4UT2JkhYwd/D8YZ9RPat4iGXBOERtx/oRHAGr2QdlOas4HHbgVDZ0+KzIiQl33i
a1ArL+NyMRXkT5Oht0UnKiLnjbNIs56SAy7LhqvHigvy58BSSujFgxyN8IYSCTRl
kHYkY8Y7+hNpLh/rNLBypdCqChK8eRt93pQet/7LhREqJvcL+5TcjG9x1eS56ZnW
ZYy/skuuGduETCSclV9Q3lwAeWPtVaVO23AvyYVIpUrH2ZV7Jw63xqtEk9Mzw/l/
0lxtLWXdMWJVDjUMKVZH100PP1l/IgfPsCzrVyYaLUJPCQ2mJolbwF//l2HIUfsd
qb0Kol6798y6GQ4j+zeFi11SsxpG9uCBVmzKe5bJWLtPWaNEga5NZKnGojeuSJhs
tGQwZjd+8x5s3AD+Sc1nXQzAImDafR5e0tNALRqDvz4+rW5XGiBhP//k6tki8orG
gbKqlNMlrnbA5sAaHvPQ+QjeS4ENKt4/rk9GtYuJ2LfAc/k1ZapjaCXaPLgkfJqm
0ZZY5zxc+uH/xoMgdwnfng1C4GRVb6XHSd+kmx3B/54uGcFMfIANxTQfHkn1YOLF
hf5WTLMJ7wJad0cQsGI7SUdFNsZceKc8qxbCPYVkqoNRmZo8vWnQY781b22DsrTL
+Ey3bRb/InoWwPkPFujI3wWW8E5obfeuQhNZtkYVP7Q17+NvR76hNY4UrqPycO03
u/vOrqsxv0Zmt6e3ARQT3z4Ay/XSdV12BWUtBh3cWaM/DWH3P+B6fgufObDjw8sL
zwUmL7shiNUv27biuuvb2xVALoZ2xBDFuBuqZCow8LebY20OWoBXxgwoLo+7Z7/J
FcKIqIwYKxNLX6lCWa405RENe4Q8FYP0I78Fc6NZlsEdnZd9P1UfIACLucK+I1f7
50zskVQQZ0AHCodCkfiCO6yBrrwdDe20yJtNpD29CUOyTyxAdpOi6ZReBAK9IgOj
g0NtGiXTNMvQhNFB7w5xTuwVxspmLN50PheqHXqE+YiviFfZvtwePOzhdSasDt3t
MXEIfLavM0rQJ0XJX6iQRdQyHuUVIHa3p0CVdzaannZTgdPMFkr/dGZUhwo+eRWc
rA42UkYctroFng9/j+R+ZijoE7f2d/qqsq3Y4YNZBEZ/qj+5EVV9hlnEJ2fcSK9b
DXkdVslBH774tzzvESqvxE/wXhkNGIbyY4PLmOaR2vEy+sRfpzlOoEzcgpPelZkn
NdvGQ5Y0OQHxWS5u/jPw97kvKsKp6HROAXBu1lQSSu8OvZjmDAyWwRayxzdYQP7d
ZHsJiHmmr7Opp6L/mJyKlXEwO/2/kliOnjSufEaXJHe9pxeXcpIWQfWE9PMZLEtJ
E4BJQNq9IJ1UGTUq+EpwqyqHcfrX32RHoxoQDufa7UHkeq/SPZS9uxqrk9aNkAgt
ydOssBJWW1GXU0jQObjM8Gy8CmQ8R5TxyrM/X8CWQ+8GKkjHkO5MU7ifw8OT9AYI
VmwbMYLOt7SKfR8BiBhntrUc+BT9Y8YflfK4syOvPnzVSK5NUh6wCHyNvc8fsl2Q
Vy06iA1sWnp1zbdai7YYp61yzj3LKRbQHirvFZTv7lCoTv5QQgTlrM8YYyVwljw5
afMhrsOTVec/bKWEF9wk+zZzHcDmGjPRsOQgOUGHkNV9cHW255lwbpG7PAjtL/pu
MMnUP3dXgTHylJPAJasfU+qPAiAvybGLR2yyBqHc4z6tsu5JcioujiXlCIeFtP2k
z6EEbxxv4cweBoOJFXWFGJHmHGf5ov1LlwUIMWOuGMwAHeuPp12CSers8wRJ0yQc
ufKEenDfW7TYWCigYh1xeVXPsK+/iwX4OvRYAkdQ8pllmo1nr/ZSJHx3xpq6Ei6b
84ok6omZbzR1+6JFW+/WUzoSEWilW2RwBLi76oGxVikVnnTBL1GaxGJh4vzOf0m8
p1jXuf7EVxYcQb2mWw2qd/zDcduMTvizT4IGOEoPw6HiwDry/5VIdSd35wB/95af
/EbKh/K9EQu0tckLjYNLLWMQV6+bZXNL86vb2FWsNTtHa18tIGYhK1LEs4K2BHyV
ap5g8zYvhjZEeLOB+X1moffN0vRX05kpFyyU24JdHBBP3/99uSSibQBg2wp/kUuY
yzqVtaeCbgNofeOEkuRXAsZ0AqFddtgWMFvpOQ1Jv6iB8LakD1nzfVpy2gIFIcpi
I2sN8pIJIej53S+DlchfMrKNexl029e0dtQ2pc7uNdmfzMEPvcNoJSi4vpoKR7GV
3JMedmNgaSWUrnSHckGbanBPN5XmJLeIKXU9Omt2+3+B/oYzUe2i5wAFWjxLEru2
6FfeIi3nBnM4J8CxeOl5qLI/c/yfibKYQ7gPNmih9V2xsMH9N2paB5jnvOOl4//u
5xRxLv7b5G6BplXjXP6Mrcwwsl9ca18BXECWMnPKpRRWTSEaEWQG1dUC9wmtj4fn
JoOpVx9mNB+71fyJQuqw+KG1l6ypyMOAIbPSL7trOghDaASVyybuAqqUgFV81Cbf
X8xnWLykGV9NLs5Nq1q9V9P84w5ulyStMYSGsljJDBrKrHD+oFE6XYhlHs7OUD/4
J37EI/CP5G4l+rfXSfts3KrqusyvEJK1RrkuPqvTApFNKgbL5AjidZ76qlryPCgA
dSRdOdrcbdqLoK4Of23A+lxbrsHGVp7eWn8kKTaVI0E7wSB9dr0OkHBYGeoQozfp
ScK3ALJzVNk1Lv/dVDLBMnQurHnxri2ZKoyhYHXtYMsTPup10NhmHo+U+JJXUlal
Sq5mNW2otC6HsdvpwZRtC7t9WOcVJz5aylE7P0wzw1u7yxvpvpmdH3693rYPZ24M
1Wj2rYpwM0bLuAvO/vXyesAw/FyQVSwgwJrIi56mYYVKYgadqBxGLBl18OZfMlBg
ZDNJrTu2agbDspCK43xT49SjiIgokVwCUJsLRWiFtVaYB7ursjgpjqMIiZcYTOr4
+AeF8wJ4zS6dkh9q0waoeKrU68J8fE55DqP4n0uvxYWWAMM2qmWZAIRHxWwzJ1Cl
ZDy1QrrzB5jqlEOY2YNdILsxDylW0Ijyvtl5PIWFSyb2bT+JsimXXRg6jC7vMlxU
GQCXteXn0GCAeSfCqaCrEgXs7nWC+KHyztmfkWrFeFzDfrK5HxklCDv1CHn2S5IO
OctTm/nmhs5L3WnEU5n3z+NVumgdKdqEQ8hIw0fkKjCVMF2876ZIwuM4IJqH6IR8
B0pySrBuZuxp7gQYLHFauTH+I/gfh9FQlgkMH+0OPIMoyYc9/OvF+mW7aRp4w+y2
F34DI40V/MwUD68f2Wj5payJJz5cnKXGve2YDv1KEl5VguqO8PSqnfm0hAmKAw2A
m4ek1XTNvDXL9GqSSyGFudtvctAdv4VlhdNG+4EDZ5OLwKdi+TIRy2Gy+Hsyu35p
hh2ibK+Vq4GRazstE5g5ycOnoN5p5iFQG0xJQke6KZ4+L6anBa8Tq7VvBp+eFLdG
5fatQqES0ZXgUqeHvDAJ5DUu+lsCLeNkqBi3HXVN4XTGy7gVs/PT0ncmErr3AC1a
auQCF45+iGzV69qM7XOkRLZlK1JcCWND1/8lTRwjWdrZ4kjLJf84DW4HDiE/D6hO
dzz/llbYUR1U9nI6tJwgTUgF59lnaagIridT6br5t4QIUHlkv5Pg3BKf3KJ71s0P
fjpHp7mEdm+RgdgZrrmUMA79z2dVPNv3VXLiNjqPyvOCj2a0GAdTFiXL0Hsf2w4W
KvdyL0jHe6ZC2FnIKzZ+6+xsLDU/B/hCFYcpiziRHEaAIKsvOOvu8G/MOQWEKT7C
Qd5RXt7PC1f7ct/RXxIgAa5cR0z+7YPcAX5NTubESE429+3LIW8Mcgv64nIzxWl/
0Tcr+dT9hVogemSOVuDekYH/pCVz4noBxPQCj/tHL+xsIR5diGoR3QzwpXttGfEs
+1krCESjrW2vgY9vB8yjR0aLoHfCtceb77TH2Tt2aHhteIxk4OvoGrM4AZBkX7Ii
UoL3dK1KsQIsJMFsIlvrtSWaDQVG3VP3TFmpVTM8nTloHiCFZJL4xdCaNGQBr/1N
Q4xgF8l/v0WZ+GEX4YKVteXh5gsdFzIfGrYl8WhZkO4gvz66yTXuFLtLs9Eqv6cz
sPIWQrK3qKur/8eVUQgISJZ27zbZRbb2Ga6+VdUs/FpDUPD+R6+2gWJ3aLdxHscN
hAAErCE1E7bqAbd57xoC8N7FHQ/qddV1ePWNxhmrmW8vMM+tXQfh+6kWL0jIZ8n/
sLnOhI7qPVKao/cWup3dKBwKmEoCvwPDgFY2/+M7ftfvmwQv3Gpv0Aa94YDdBOD0
vUnlji3it8QVK/yjBJkTFRpr7ut4CjpeRZzBz6u+RInis46y6J9m6fH4+fxmuVcb
XfkcYfop4do1KzzUz8Q3uHYbq30mppTvJZMXzYKT+ynjfnFWW0jg/THofa4gNb8K
rmZorvb68SxOTjU2dGDo3+ydPXyQM9nHXZsucPn2ep2acGG5PZsNatOB3veYhzrJ
9un4C19dtqTaJ8mGcGhbdCI9NNJvIC1InP6Nr/QI3QTjCCNnMjPwflq1VnoYpLeU
z3ux3uTBXCYJLHAuTsz74vyfr/pttwV1bQkES9Ggattyo1cwN43FwZeSs+lOK32m
oARAI+VTLlguvR2AQDxJ0zZ9t0YfQAOI1TS6WLyR34c2BaFq6kb60z9rKDqaGLlb
RDIFju56viMjQsEhisxRD3Hu1pdYFBFe7914xTzetSs/JHWEiTGirCgLNre/SJE0
YGZUs5Ovbm0gKD1N3H1V4pW/rd4XrGt+l5i106iVfKB1Bs1deKSyEY1y4PQ+koeS
K6+Gl5OiFYcaHb7OYwBIFPeYWFkF9FrBSwD+W3WIx97X9JMud2LWJeWc7JkELgGO
n0YE8zdkNJ8CniKhVWJhIkfdOYhIR46ajpSfteV4rg68YcSTE2pN4FRarxDUczOx
XdiDeaIC1F1yNH9x/XWM6gnDSTyJqphLVgYEjbpIAVV2gjg/LUgo10wU3F2UQ0PA
H7XJA3orS4wIb5gxNmXKsAnbasjP3fekit9DW4MNOuL8OODkXypmrimC8TWZm1Gw
oR/nM0vNpvJoCCo6Nqg2nUDo9BRw1RSnHeSSscADnJKcMw8nlbsevNcJETopma0j
Uo+9RTn/Pz1E1zLFQ4iU3uzjyAlVeDx0pRldXefFYyS708e+c+B7chaNUF12zSdG
whb2bdcb28NVJJrSEPxHr57BkjFD4UlU8nHcW3Ua7JvZg8zmRPI0FnMxyUhwpWkC
rP3EXn1BVaaQe73axcQ5ken2WxvFq7awyn/R2lIOChFhBApNWhB/Mo1fdeHMCPov
Qkfb8Tp8aswN1rZSyJ0zZVoAUrxoO+L2h7//xJsGNfnoBsW6V0/U6sWZ+vjQlBFG
D4xNwIcPi6NXQMGNek4swA4RJnhHBCKrpM8Enp6p+bWm8SUqHE3D1U4tYKZ8Assn
hQNAhseWPe9sgnsJbAR8zNwoHRQMhoptKLfEC24ptuptoWHBXFdZTG0sOp+NtQYy
PNGwXUJMtY1KyzAOPRjeD7DsgHbEb+wgbjKxJUH87Y1CbVmFkGcZleBFuFesMeMR
9bqZRy/THUXvlArOuTyxyRki6w6kzqZQQ+KFxcZa3zcd5rDKJXXgBhiZkFI3xm7p
2Rm35g1mgl3C3Y0DX+vftNA/+jhy8iY0w1V+HAarE63jVxcESq176sAbcFM1e8ra
JiLYa3Vdl6qs0ko7E5Mm/j6ABU7QRHUob9wwPFa8lxY4JsdUB1Hpb7UFgxVBnmPZ
tZvFFQNyZewYXPr/9QtxmKVrsrAOJZevvNQFDU584p8nkaf0Bc5BDzbR1k47vShd
Q/Yw/4orybMosTgUZ9IU53HD9Cwn+o8gQLS0/Jukj9NQyu7Miah/5jOhUKuS+180
iIFOjtXon/UQRHZQhIslBqWLt87jlI5P0bdW2uRNjOJF4Ugl+jMX1FePVsqguzYi
SZ2QruZOf4aSobeHb7iqZyZhDDYHOvKGQih+JT9HsXpEOfiI4ki90NKY1FF7QLnb
c823OZ5e/2+645XouGp1aT7lV1UHGU5iSCnFg+Kv4VgSWklmN7Zp0Iews+WjFrEa
1B1FwNuLXwNSJ8NcjLSe7gK72G889Wa22e0OPIrVvJc1N78V80M4L0oQ+jn/DLxL
yG3dBAngMYWz1CO2b0gasJTJUZ32LzlEpgGYC4tjwa2QFciIzYalJTXTA03XtfCC
BIXRf1xlZpeiooHmRtB7HbuCJAlRQZR6mXj2s+m7y+B49zu76HpKNO64y4ztOoSi
99foWvXHzJFjQhPJzOE1EcN+WtqojsiWt4c8Gko/nPIri9jNUVj2mKl8frHgiMdb
e7fA3Bzu2TnaqwOUxUJfWALM6bJ/wTSslcV3/9Z3AGKZY+KGWKwl7khmEHAV9aof
50DnzAh4IyIyBYxwRZphCK93OO42FKGwQViW8rmqr2TSGMFRw+QsEV1wydvNDzA8
s9Y1VNUkAqAE7SUayZPH5NcoS6zqNzgYVzSHRcfoe8OoEMZEQYI6zvVZ50gjPQ/s
bt7/eOGEgQH70YTc26BwIXiGk1Cvv/z4nlWFjssNv65pOT5raUXG+I/wUVLNmyMj
26qtf7lwcuyrnKpUEM/mPtJiVyAR0SfslWa1A/SeQus0A0MJQZtGY/0gPjfQp6LA
2s/3ikTse6uGcUgilE2MtHWiC0iDQzKLfEv2C96BdmPfU06hqNiNh8C/5Cg3+oru
gAouWbVdakb/RXyGl903BSKzOb8cxS72XInS+8ziTnGr+BEEzFGJdFc38tPscsna
4JUnqSreNi/8f3GaaaYvM1SrtonyPhufIbY1rpwJWZAWPK6IK0k87ixL1WEk6LmY
0Jf+VU8n4K+yy3WOTq7mutbz5JO1f93WN1e0JjfUH1Jn0A1JQrJWHPTRYxpMlxbH
jul28JPOLlRVhCMgDT2zUR2l3gJcSR0zfGCqvukakAJsXxJ5lmzGl5P0z3dxXQad
uOTq+1fTcIxIXeAve059tnuDuxoXgz2PUWgyy4zMC0WHSEschBEUIuMZdPDE7Vmc
IDCtz7ClZposnCgimOYKcMQ2oE6ZiFuEGP1ouAENRJXh30JR7ESc3ymFntK3vHRM
hSudNOW8sXG3EsdGXQM6mLUS+Cj6ZMq03CuVrbLjJrF604eGo1KXtOu09J3LwnAs
rxW03PzyCdwSw0MZaqJfynSBvqXl10GVKkqqZCcdD1btdr3s/YrPRFsmIOw4KEcq
K8/34gYe0BLkAAfR9SO5/fkqsiZynSCktw59jccq4o1rP8XN2BcN72SV3OON8YbT
XhegQBLAHmVV48gsfEHocIp/reN3tpnJIVsd79td/In1ipdwpVc2FIBvnOVB8Yu/
q950Wlh1UXKEigSJDffHobC+D/7/URBaK1hOALMlEyaN+8fkYSQNc/CXQsJKiSFO
9OqRa28+EDvzJa1UADbIYWgxWhqmZNmQHQDa4ugrMnsNPhjK+vWTlx9H8klU+/BM
b3Wc42nigT/k1GaLPh9vSJUJITP5NhgG15ignrqbROAF8k2srIqTkwDO5ymDDZbW
SS33VJ8tDyNGgn2FBFOe997RepD5JKMSZYYiyJULg117mTnQPyRfAaUgeZfIef6F
2aTXwH0/QBRt5gnQJ3sBZR5KgikYQ22s/CAKXectuFWu/bnqV9IMUVp7AtGlFuIO
S1S6FPCAlx7kbmduEwW9Qp1PoHq7o8JxfXRedTrfJAbhPd0in1q1tMptRXfFJiZy
OdAWooexfk6e8g7s4g91bTZGJ2rxUVZKz8J5pTUfGHcC3RlKbZEcLbPXkT93ULYQ
Xmlo6aUNPdotgsK1JbtBMGWLf7ZkgAELLrn5aflFo9E3lRxKOBHXHsDKfXfcCNp4
gVKOYl90Ii0uwdMVO5UiiVQoPkqCEDyAlngPD5VfZUNejR91CKdJ2WEY8BSHweij
m7CkOnLajvaXcPMos4E8PUdzzc8jizhUPreNXuMepI46M8kc88LnAD4X+xkbUc57
sc8oyDuQEWEP4XOszITzcVtMkc9bZ3VYyqran748yaBUe+KseQgcI69Do1bd30Fj
2gVmZJp0UELs9beRcBq+Rqz3tyEmvmXUFyUllmHNVLTkbcFWEicGS5+STDUUdOZ5
ly7PyMrjDVodgqL240b1fT2ybxiftTZKycKjG7YLRm/7+7ZdZu14gfqDMPi1YR/0
WklI+iW3eFBy2puCqnouBvnDB6vyzNHZA5mVZkVb4DetNV5xC+lXh0vJwqn2dnxJ
L5xi8RCCIn+b/5rIyCCpJmRGrwT5o8OWLJZzVWdK0gIxzpIyTDc2o/jyz9Xnh9ek
3Feba7XfkA4xHFG1ari9TzQ3j5mHDg4S+F1MPcRqVaxVTwHP9MGqnUYeerKO5xq3
JvEAO8hNoUokTcdyb7oIeA44A61jVWUgX3xvdMga9IYOWJZ3/kMriBIxa6CphNWi
d/FiVZeCqCUSica6Qszd+Dx3f6uf1kTpfp1e0R0y5se7oqh9xOlKxcpSBMlwc4xV
FUy/gbNyEeJlwb+wxEH3fO9hTYIRem9rofojKWdNslHbKHzjiOOvDNSoG97ion4v
OuE0jcZs2rXFlwM7xOUkiutbXTKA2abOTAk+QIjiFaY/kktZdiBCFOp/QsrH5Ymw
ktqLBTop9GCmzDJXexshn7K91lbQ7zibE54fYFoLCaceHnOMgxZK+8y9VNKhWgLB
W+0eqzSU5DnfrcDVxKG/UU6w/6XGq6v7ycBDBmJFludKJPltdus9ms9rqdl/px7z
j1lTWkshnFOQ/Kf7fW5zabjTtFslo49F7qCzEn/zNZlfsIyvVd6b5Kl0BG+P8HPB
NuMcLOAxlfD1t2jnx1S2lKZAhUrfE0d1x5icKY7K3g6Wdmh7byNOBwc1+A+kMwOR
MxsqDfM2TXQHmxlmkKBgI2bfRbe3ujqagOratA/098Yu+KcoB7HHDQms/l0Jubv/
fdMji3boQ69yCt81UreK3IJsPvMBxQkCg/GFRVJXJq6WOmHMWCkGjOuaeThHYxyq
OFFh0nv5ynzRhyszynZX4aNd0+RZfNvFGb5ACGTh26otg9zMVsV2llJFmZ4m1jLa
gl6QXYzwE+gi3gU9gn1FQdrv/RS8r1B+5mR/iHd4pBr8nMVX3ltL2AR03Mhp51Jf
4edQqHY/osgsyUoq+By9MRvEaAujSz0BhrAT53j+s+0+VlKyrntopxx5YkqDyXpH
aqsD53qiZcEszEXGbaX/gI2OL4F3VBqXu+XCn6/S4P06E461X/USmBkmNYIHi8K5
vrxKEfonl2khR4T5vpuZMceMn2rKyj/YogOlvdQrGB7dA679kG/IW00C2Tt0qBP7
37JAuZzwrBRgdq4Uqm3Btp3QURMqm6By8Yudc9DIZZ4r5zFf1/Rhk3v10ZARm9CM
TUIVkohuGf9GndD+ic+ZWp4qeaZJqk6esXR0gb+mFdcnmMaWTzF1n9eX/zaIWqCk
utKQDM5DGj5tdQtsbi3FE7EHXrBm29EruMKkH85YYun8V5WThckucRny9NII2KWK
w9ctfmTulLqu8VnN3FEYjMnojIKzkhUbYv2fCtHPx39d4h+fyRhQff5rQ4B/WqeX
WWANrHbp5h0ZN469DiGW6l1sng1gQmX18ahA+W1joCuXgywE2rfR4uWthhwtjuYE
9MRD5OOOdNPdciMagJ55/oZ1zfiFZWjzYNJmThKlKZA2jiNkl9YD2bAGZwsVO4DH
nEd5J0/z3LYdSbwxEqrJGGJfflptT8ehz+DPOw1T0EmC5dxeCtDZDYKnaB17MErt
vA60cELinuRNnrhNVGz0c7k3ghEDvxofBwxFv3La5u1V3C8GedRSwdfYXKgcsGHa
lbzymcPU01ru8PBt3ditZUqk6yCirvPMXVGtmUDQk/QpnqeQmM9Wp2cJWxkg2xZp
qppvmq5zrTwEb/ibFVQaWoxEYryIDlKxtqhrbYJ7o9i3dUNY89VC9+PB3+7Y/S50
ZWYPl52U8f+T+vVgS3cR7SNhVwAh40ZGRxRTR/rH1WFynKPev4aKe8bDs1xGQf/P
f8MP2hkVhcqmW0ww7+3ZuGwdXal4cxjoP1x3rAmOhvfiibw5cT8zuTVtiwlaqh1/
skLKYfLOyhtfetN/8Ox+dX8a74j8OWDqcbBb481wVwnw3hveuIrp5NB5FVtDcF80
mMXPOy3vM6q511gVkyg+Ojo6P+9+mNPuJb7O2SyV07j3lMSETVPMXIcR0DnnaqHf
uRxry6LfO7aFDjKcyRYyfdiH1ENxuNJ8GuQFo8PWXkxurxL/Vb0yUdWvcRtX7xY+
n0hMsKDrD+twql+JYV8NUQM+rYAwlpWA3wcdTgO0Lt2BqG0UjIO94LDbtuPqoAV3
+7jrpPTdP7f1ZtOnFEO/FORaGqgwTQTxvCSMdwZcx9tyB6fTl1FY1NijIMnuBov3
4gtVc0zr1GkabnzutLs6pB2uZN47/lwoHU+SxyQuzTirDxH4nueAhxpBSeVPNyHI
gD7o1PYDCIj2CQVmAnWy036jjDc2WkTPk+j2VO9kzglRqjPcjRMs7GMXinCwanhC
CwkJ/A5qw2Xcjc2Yi/jvzZ6oMELD1IlQpMMBKIOkThrlUbZQ/RUHRY+cdyiEgSYN
JP9xHiY6sOQhQw1E8NGFfv/VO2LiPYDTMlt0qKd1au2osy9MJkhyWtlkz8OCwIJ9
9r+A1eu8duzVdbYQ4PdSziqU+wi1jQo6pRB0mIqsIRa7lSj4YtaUsjhW+se+l/OO
jwMOEtf2dBOXmMpkXuCHNHGwc/7kpwbaQCeNFwmFJKrykc4PMST3UFeEdEDKop4v
xQZjewyoZLPzes17Fxucl+PUCZQu0AZos0agZfzJZ4OkO8WG9UWNh1nipuCcGx+g
HBulaAohDOZm5cvhWTPoIl6rBoVydUZMSGBWL2SHb+GZ6owtLunPbizbj7RYxMKQ
BklLz2eKmX4f903Mv0+L+UgrqEjYf2aOQ1mzJh1WWb7fc9U1gS0BnHB8CC7HlplD
wL4P6JRA5FaGtoxk6m2P+Bj1ZOSk3klmO+vhZeL/Ah+rxNEPk2vF3e6UfhidZZek
z5BvkSFQOtbHDlaVS+TkT/M5382zf25bPzzMOVPR/c+ME+1HndeT0ZLRikENzN74
Inh7tr/3vqH9OKi/OWwzT1mGlfYdUNA3h8JjHB6q4/QImIRMRXby6X6FBrn+UKSR
JFrnzoq5V3AEDxCkTZxBDNHi0NWhTfTk5xUi35n5fFKMiBz2gq0tojya1LQeaOGU
TSCX64NMOL48rhKZvxsi6SMYTph0TlxlOTgbQhgLOwaiN0s9PsHJyz45sf7OaFsl
o6DNzBbrUDzF6Lu/k0PsMlv8foPqWNznq6LjTsZceE3g9Mjj3P0cvTbK/T7HYjpT
esrDou6Zug3z5xN8OFmBSV9FmQzgHp2vKx/81HXpQCO2VFwtf54Y05ZiJrl6PV1v
Aguo9qBQpfekOE2u/3ZJm+XBd/rhtWMr45ayTi2tM9PONw2GqY4tTMhBw0AIkD5w
mTbvLCbSuauO6K1U2T/f9cTbAvTBytf5BGRAbEa9NFMxiDJBOIwEy9mPQv5UiiNt
pv+UNcWD0AmpuCnMLrDwnnpCWDr/Cs3L1IeWv4ez22VWg+xvL9FprthgK95z4+B5
xTVybx6YW+XcIkjpiZXm1uXndAltAPaaM16nJyAZji5Pc98UZLbYz4194pQLYOHn
AXfOHtHrDxPJmWLn2GUQUOXNIoHcDBe++5T88Y3oSliVxZHdUmyM1n0EVhnKiRIy
8bvENk18we4Q7FomRBpeSaOi+8MvPv9y+ZHbAbU4WEUOKOpzwYCWLmHKWPPZb5gh
JPzopngAHMJgB+ii/bTc/krwCFqHeIeSjDnOGc6HrU57g9c5pq1kwGR+vvl+80aH
7CrrTIqBmHTYvqI6m3k2bGzmU5rsm+gfHaWKhtkFF7RcBwYPM8Su5P3gOogEtvGq
b3d5gOfy5kFirR22yE+ipoor8EFWqMiYGPl4hA+MIS8qH8MPYB7ksvilPboZnKC6
TlJb1jdVsI80+Z6uoEAmHVFbDjsKlXKpxDzVBYM+EvT8cXojxbo3WD5iwijkAOii
PA9lueT8ngmXTRpN+CtbDQl+AWZehOBloSW+ENewyckGAWb9cIYKKfd2cIkiBwKl
hy7lwqlBavFajpgmuLivYedPrdztrQS/ZGULSTvR6bwaKM7gUKEki4SB569qaIzt
dgxkxOUy6hJEuddzyzoJ+aPMaAXEiIGMfhtpqIYDYof8KggxUZMTyToRlJ3CB6td
oYasqL4Sf718ihLv4ChKowL0ErHKSPJBLfWXw0q5H+aSgPxpKboQuxnLeCncwMTu
bAYr0F9famhnJp7oXaMdEgqimpvRbdBljQ+VudUnXp6EvHyiLVSXW8TS+feVCTAm
pLvuWUWtM3rpOenRGFUiZQ5k+OFPa/RCtBzjt2VIV68TN7bAV9Nlq5fJV4jRJwu4
iH4JlI/OkmtArG/EatAZvSaRSQUT9boOwa84Vn+3aL3eoTVGGcNNLigGJ6pCNMT8
20T6WMWbhNnDZvlqDUi1XKdigNg4flG7EWDWHZOA/dnvft9McH81UKAOp55LkB7R
LZkUtegjpVZhVCZUi7/TGVz79Rc8W16lTsKJLfua4XIcmS4gZeuW5DnHP5o7H36M
AY6coKTrVhU3RQFmzL1DZi4OW+tp7ziwPpMkGokcg5dVryF8zGdTSqq7Bu4t6zo5
PzHKewyf6YmAGLntoYAFTJKvBrh4cb/6IKdD3KrS4oeUz1ux4a1xLVWi/HD+X2bD
ZQLwDh3/rF7tu/05DMb6btN41Y2HbPhpl6eNf44q1YjreAjql8fyyIHcKU5vTs1v
i2Qh4QL2oHOFe9kKfc1PzhYqXCPlm0azWyVlmceoXNoX4OucZFBqtXFepdy3j0C7
LjpthUYLZEJCuJF9vRxKFJDZGWEiw7Euf+5Os+JmCuJ4Fab8GsuYycqe2GozhT1a
9Oh0BnLyH3UxeKIMjQf4Qba3qXifK6R4+QDKF27utlKcFRsN7V/XYX/I+i6/rwYI
FnFWJaPMTi3x5A7k3rlSwWlD9mB4GgY5omASgrT2g+fSJlVd+p02sqhXJu31fsgJ
mhROgGZ5wKo62KBTZaC+4Q9CFc7NGiox7qpYMNe++0xKNK4Xd6VTRCff31Rt5ge3
neM+kI+OmApEG9dAPNOQ2vwRnGpfJUFYueteVlpti+QViUceqOkjk6QDxbkubHaD
sK0yonvfBjHfEZRC2qePhYUlizK2q4/0ztPZDZZYHhOcF2wAcwlHCI+3JUUfIKCt
8nxMPombYqToEacqiJStdGCUysyzgv/UWE67UvzNJlGkzGTS7SPq8Bt5eQ2pryIt
7DkO6lqOA2sj7N2jMoZUlMBAtAzvHG1Ns0OFKvo6BDJm67ys01mwr/2ZXndXykmm
dwUdDACV2myMnnIYW9PW3bw/3KYW/eOX5dewW4w83+Mj0UmgT7oMTztlW7VaGuS1
4EqjI9oN/Yd366v56xHrebdm+YzvrNMqb3cd+ohZ5AAAvU7ZSi5cjC7Ic++Tf1YY
4ax2MNIqSTBwEuRsFPWFHAPTSCzrcVWTPfXjnu+LnWD8q4CeKn7vbjDg13jjc9ir
Y1evP/JxSnIl+fJ2dl8jf150QS7g58W9LAojkZB9W06xaRw0kwhsth9xQD/prq0y
dlm7yNZFHIb+EkhfunOgtKUoA7DoA+ShsnsYzrzupyGMsU7+E8HHFTAE6BvPiflc
AMEs0zD2YOvU3olyEo1+k7grcW8QgAbpkrj0P9Ec3EiEn6D3ynGL/p6PwXSDbw3L
GqQq6uMUS6ME5IYYmXv7h7YAyjZAphP3JT5KRsPs4HcTxxGOPUeMyac4l/VKcx+3
8fJeQYxNRZr+wje/mLOcpnIbrg36+7rM7Ezt/iHSJY+8Pn8L/REoM9bxFxf9XzY5
KQ7x5K1B6pBaCxLHhWpRbm7bNdwwUQul7lv5uYmIZM9jHEpPHCuQ28juY0Lt38yY
N1WO6ty025jAnU1vHAg1MfS7t33VYnCVG7gO0jteO1ylNXHIzgtXJkvtHMMSvmK9
ZwW+SRiKPBkjYoIxaKNYGa4oWlHCqKXDKYt6Mf0V9LsZLr8tNhrnfisTdF/oiTes
g/r4M/uSfoD9VwHC4+HJJEev4IAKVxRSYLjUC/GkSyy+2Yg7qjE/N8geH+ocp4Rc
sLN4CkXmDbJh4AICONsXJR0A9HdS6He9mbn3PwJrjGboQMICGvxXfgmKv+qwpQyC
Bmf5tcFU868fmYnif3r5gqr0EWVi1YEsBzJFrGnUP5p3Z2iqXEkaVMzOzY5hjvSR
F0EkRUfPEnzaz16FSo0LpwDrfK0gJDROUgmMKj8/Uw0+cbmVcpgpuJ5NrOuOmz+z
MTdh13c3pvRwvOpg9+Ki+acdWuT+9PiYLphPHFxwGJhJYUW9OUfgKLC8wlVkdiOD
mtA0h2MC0JWPruoZNfRm3P9ic7g7iRsDeRPPdHJrEmCXB0aQK7IawxkRaYh+KUmV
Mjs1Pr5AkkgsmWD9S4sqIRY9CVujKZDhISQ7SsL0Q9L4/iwLRui2+H2dDibezV4e
GYrQLYAp2E3gSiDQp+mhRXOLUIX/TQJW2cP0cKCs90rLjH1qAw13nI9TVq5GKoX2
MPJxjt9TWplopJWkcfTB+jze9aVNWxdJcS3GghOr5SxnzJG2RRNO0WVcqk1yOSWr
nEdwXLqlTJufD28TyXNOo2lHePv3/lNX+om+4ajjARK0wqNTEah4xQEhtR34+wpT
ekLPDXUfNKIbqfEkGQuocfizO+ufmM5IxTFh5V4RcgPV5T2nEq/YBGkLweJtyAUX
Uh4PtrLocknaMymw1J7r1AbvRtZmWZiGCyck3Quq20AsKUSKvZ8lvNVHPdNFjsJ/
PGyMzca+5aNq9QNz174l0h2IIB+H7eIztXWbiAakJmFv+KaUvAy0PvHSWHmZDfNo
9d3R3S36EP1DHi0vZ0GnlkUbEW1L1p9/JzEZYcdbY3kEj+NZ+s8fC38D+UP+drK2
/bCTSuk7RRJkMSQLSwwkQLVzXmiG9FczpEBoaRgjb8R1Vv6ZpgBiU3PzrZHxk7cU
CgymF0coQELKlNwaFIXzkyieROCbq3/XMyhcJpkjg3WIanpqD6hUqeKxw/QZtod8
GG73f8cjJroWH8VEa8Etl5qkMpQXYCwOh/WnycLRxRs+j83ei0Vp5mwVVfHmvuAx
b5VPJWBaCOT1IOMoQol5Lkw8FBSy+XW/h8fvCmprQVCRDPzl3Udi8PmfznGdNbzY
mxfUwi+qPH+IRUQMcO4h7IrACDzp0Vn3y/L9UvyW5FY33h91khQfcG2NI+7qwTDe
MQ8GuQk59dFL2GIBmWnrHJgcfDoaB2rBL0Dnkh779/1QM3Z4ahQqaoh7nY1z/Ybd
3aPBPnm3cmU7+j8rh28QgsHX4OCyoL/Mx5MEMvQo/wGl3B6KpoesjTzRZyVOxt6K
yrpl4hRKEta3f53fa3IYDVYkFwYh4jxiE0xdyILKmufcNaF+qdRJhaXXtHwSKECs
+TzIyfaXtNjxS8ynyV1IlSXJLhWTuzaOWAr53AHjEiW5/TnKo41elFF/C6BkXagq
sJsKZAYze/BxYLTtCbXe4Xgo/oXIT8ZSxiq22dex2Cj6yVOfxMuOdZLbQJnQ2rjA
4JuFDFvVlx5+MwXSyx+prPuJMpf8iw+VUaMuwALMvGv6RXtf/ZDA+rKsZZt1MMAD
6g7vdphxqwsFSHzYmGwPk3XKvojgluY+Ao/Oq75Vkc2nTktEjOpdgtKdWQfaMfoD
RRXbN89nO95zURVVptcORblSdSgB26kEgVFIvvqZcoiQGXbbNerl3rawq3AYeeuN
0XHzunc/OERGngvOe+fSB5XrujDiP/CrNbvpiPdMIo1FRVDfISmIqp4jF7xLK1tL
Mwlriyd9O6UVYTcrtcgTA20GSjWhfpIcduvaoiziQ8K7PPGxExk4STDIARXvpR8a
axBBCzcn7B88yCUGCbGNi6y6selhtQGXXQWFjZIgswQjVf6suYERuMKHWPw3vMAl
55t8x0371vaCHSUxDbChma+6o/3oq7ism0awRhlF6iGnKquacBu6n7GOtY8AD8Yr
6T0OgZqIdAL4rhqnKvf9lDiA8lCjhNZezgqb7ScISNj5J00SezN0AYCivCc8+CzD
CW0Lc5x4yBmBDzAIcbzZZ4QmBNR2MuMZBjtSkRXdzID5k/okjRnmH0PEpmfQvzaC
XZAT7EIJUTcKvBL+OtfCTbDqorW0QRGcuVY1IF+ssglFZ2SwqW+uDiM4XYX5ul0Y
QYe3qieFAvAlHvMEroqOE1oYki5xolxBiIMQdm0DkxpKiT92jbPNScMCww1Ya/IS
HeFHrNPG1ZxnAOa/leQqTFpRT4gVAIZvwmhK36TdNzBFGepckSX7UtwvasyE3IQV
SAVgUfkFzzE+3RIzieA9t1cnjpSk1DXtgb0XzBO8V7XTHbmmVCIqETWvB1n7maYQ
bHly2zjsFNn8h1TEEfzIfVGuKKC0snshLRsxX8EQv98NvShZ5cODM+9946VPjkFo
kBYLUUcKKKvKFbzWBCUun52pDbVy7wDTgV6u5Xxbr9vmPV2VLhEXhkpP5CnrodFP
BdCNPLPb/JuWDjVXdm6z52uIydrN7hHzINlf87WrGxSfUYUUhsKejaNzWa3vcVGK
8Kb7QrU4RVVMqgEvb5L3H9Y8lRK7VQGhoOyR0BfvdgnXGAVbm+ZBvEWN1xh/dYuF
/NwsA1hsp0uaqnVT7bxvqG3WbdfaMAj3LarJSrQc6tea3LqMiA4peQK74KOU0SpI
K2RhxkqiIv+CMwoIw7gFy7uQpCHPGtEVBGYd5xSF5hyggApdHK92UyrypwG1nM4M
+hR2WM0XXbIIshmTf/hfNABB0UkHDSutmFwJ40eO+7DK5piy5fEvn1ggmyzjJQI6
ZGcJe5Trlqh/xLoeY1aniOUWsH6WBuCacGSfA5qHnIVQFmHyOjhK/nr1psafU2YD
kb5OQXz2yWweQbHmunQI89fhS5RYr95fHmIX6N7qkHavDDmZe4g61bjhSRQ4PSH4
4UNG+QzD0sGqMRbFV3WpWu5LLYeYZjKoajNmKqdhMhe7mrJkrWvLYWFy3Os+/ZW/
mNcTojNnodHPdA7cEoELkeoIurUOQrgbyerILncBxkKu8PikmrIFxFvPj8tr9Ani
3u4lu+S4syYbx2yzdB3ayb32FfTxinUnvwpWw8MgeIbB/R2Au7Ll8jOyz0yk+op8
te+esC2yvQCAqbONAZPoYHqsvyQtuLmbN8wXQ4BMZbRdNEbOCbThQj4ktha8t1Zj
tY5NJ2ptQnU3PDEKDvh9IOfRCPV3ldF3UlhgYVdoN9+aIbqmExvVsY7v3ipnJVBN
ZWnplXZx7015a3vJzY2Rp7gUqezn0x0xamQKED7mfWYvnTUx2IJniZmsP+d2xYaG
DZfIeYJPyFUWI97QpDCI+QBePAIDKJ+TO/nNPHG3EiXpE9/EILsoAJaqTMX27r6R
MaQmm2cWM2C/5/3RAmx2b/c+3ILinGZgopg0W6Jeyei6I3PtmCt7F2f8b57FTGtM
5ThAQsDRbkFXmbCN3M2UQK1SrxsNhT5eY/3jRot4mkdKvfr1qZ6RBpDeb9SBS1tV
BR7jlByrZjNTx+QNiszVKJFF5974NXPxco6RhgHS827qNMzNJHIQCbgrgSFAJ6Rq
KD7jqDMft5EiPk62ukozh82K5tP9shEDxhl6HkwpLy2Vx5tDv8qisxntAgHFjO0q
emuvnJUdTDV0OzlxvKy+3rOTFUgtoahv5T2y4TwzcA2Mykw3FGbbj1EvYeBZJ/Vb
xY27Sbc3mSSk3vvUWKzjl+uTyrG2c+hA/P6W3ej9e+87QyWIZvrgw0Kf+vL4T9l7
IMUzQ87AUPc+TlshZLIx2xP8k/u7/S9p/AXDLXRzsvQs4PTgoeCQvZDmvJZ49hPR
PVR96V0juDhZc0zUGj2YZP3ObfvL/uN7kiY1qGDQuXRPexRooR7cO8rOJU8hrKfq
UdaEgr3JToKXMXYVUVX8Xvw4UihCaW4bWzMTvc9mNePshsSi/s2sdpT66cajRGYA
zYQX2kAjWBI7WVlPQEgyOk/d9DeTxnOLSSta63oxYGiR5HfzDqj3ClQQ6pZiaKW/
8k6ek3wL+5Ry90ZPj1bu2Iz3MpeWe3UojhONyD5xwNWtBALk/7FpUkpPJJvb17Jw
6jurPkG/sOIvI/BVqTDSab3/MjWRWBtbsef77vtvYnJGheODOjCVmtRacFBtRmbM
52uo9nOWy7ns5AqBP24eoTyrTKYPurtXXBh3hpP62sM4E7YeBBT4cZX6fjsUphPE
ackdLwFlALFErnsKGCnWXjX+lT8YVhm/sgVUedxriohMYWu+CAGNlNFew15ikV57
GkFASHHS/mW+0rJ2wbscfoDUhDiN8l2Jht6nYesvpGvRIbKwBUqckbJ8Mc5RPL0a
0G8OV6thlcct2LwEckOdqi0L93SSesUGyWSViTiEpaR6YLam3KNICGhwpEj/Pw15
5S0HoH5WChjsRhimABEqZpwV5yLNbrba1sWSRfQXuDfyCD1Q/WVHnRuqELgVR5hd
gVRtHS2DBNWdWfOwLEyyO1v1XdE+x7E5fLNbvRl0DY19pZrRXhIEfp4eLUcy/6wM
3k6MUiXdrwZwzHqx78Sy91PGhQZnSO3q3juj8qf4mMMZVh3e+Av3dILsWz/bryei
ZK/RS45ml5/Br+0J5vv+SeULoRclcoKm8qQ4X0HFQEjGg7xd+69fsjfxITD8D+wQ
ef32KZMMPhvo3bFcq5GiMG1ms++tHkX3WFGGTB75bsGrN/gl9S2FXQPik3D2YzAi
KhcgJq3yTAixZ9+uYxJccDA/0CYZNxZ+HtULxQP8UdHUo8LYr+QYzCY/6HdoiZbc
Tm7Lxn75BouhcGx2v53mY57lQYpvu/mgas4aOU4ELgp4W8uc+wlZLsB1+GOH7VnL
tlPOB9W5jHqGVgxzUMfqIG3iiJziMM7DvT3wOoS7fY8LL4JHJRg3MZGEo4kUEjwr
DWQ5JJtzF7vtoJmW6lWyhxhyc+xf+2VoPdzYV8e2rcENmDF41Z2cGHc0szDqpPq8
PDrdJpCpbpn/9j5bktHGthY6ohAQ0js9TuNNaZKTlWjKcmYqGC8Tq5Z5c4cmoJUq
TYJoooAMe0fCdZ8GidEEjy3AR07w+eGWosjYnzPlM8RLULxwdwHwgKQnUfF5TOmj
pHAAVoA/x6LD+TCVbqdheAO1pOBuagCmE9DB+8DaK1ex0bKPqB1Sg4gi0V537cez
m+5kbz2l07pLvFabOV2YJLX3LN0qdvICeFFhr7ww496oZNQij20WC0iiN0b49d/S
YA6dVVdCZnKGjCfq41rC+/KLhYVSZ5qvspPSOw3M/4dpetaDs4SSDJMHTdAJz3VQ
UF360qPEY+CAU9qn6KPUF7LGd2+3Oa620eFIUjCNEvSQcQqk0VMnorOLkODgnZ38
He+bkM83P6uApoJ7p6VO9mauc6pjQXzGQ6KY1J5sr9MfKlPC5+eOYgYF2A2jNjbx
SCtT3rlDyV3k+FYKZF97Ox999dp5VAuHa3AD9egBesg3kAvHdNWQ223KM0sIykLA
R9qWrsd46loSOxwTO+tSsE8dTLGu/JSabW5RXT9O/Y4spd5BbN1/N9Y2HkgCZDyQ
h6aGEFzL6C3P7yp9V2VXkojSUhT0A3qVAHadZ3zZO5akb69cVHv1NCt+J74EVfOD
Y9c9EBAtQfbJaOqxq2WqILFl90rpagRpvjvW94oaoaMgNlSJ+7aSJDurLz8rlJbG
AhDPaxyYmBTcjJV6cdIy6mD7PTdVaeOdXt6PRBgpCQz9hutMhmvVGGgMAi3cv4Jo
na8NvYhw2joloxtmquCL5ejLE9OXo+ySEl2rekiviM3b0bbPOi+LnaXHTeQur0oZ
EOS6OZsFzCGVESUTIiOCZ5SVZVNxV3H+Dix7ck65OTOXkHHxCcFU9JbiwJtCis8C
iDrxcVln+P6YF1nCWJBABg+V4UlWELc2mKOS8I4KU5aCvDeMw4OY0QJ9EeV7nv/z
3ic+kCRG+EIaa7BJAnLPba18UoSrAvfoT+8LD0laOE1OQS1Lf418v8a6ViivJN3H
PghyHT23Fm7Cq+l9n1S9gBzS5Oi6ljX7HWWgRFESnNpK1Y2/xceoHXhJiVN1DWVU
2NFTDI4ZsytGbjtMHImfYfK0EkvbCMv9C8CeJUMAUekFZ98FzE7ZLAK+b6xoSM4z
Gc1P9EBWKqBOnXqIh1OjrVGeQYKBdxrWjNYhBKV3N9CDm5c5OZaEJ7EXzHFMwQt8
FtC31as4fvmBR4wPoNX/jjekKKgblyd/YfQWuyQ+7C4Fs1bXSMJeoNfLCJNIC+Rp
Llx8N0/gy1+ZLezEoU3DExreRzaULrBVsKhTvUczZzexaKqTFTzyLmiP5rXqmPGd
L03yqlIjQFvB1Yt6r8n4ZkPVynFTI4dPHDiY1Ph3//NPSvxc/wNYdGtJhUMwr2mI
oipq+nbWvhO/DHBSIXvDhTf36xttSUHX0YSY5PP3E66lDSdvokMjXj0kkVDsYCqd
+kkmdWT+VI9nFD0ar8q2rq4SdAMZR2CfC9kRdOOvFFpxhUZ9m31zJLto2ciRvLxm
jT+lj8u/VfbmqHaDAyFdEXsa7o69u/8gLCR9FX+q9ra6M21pfhsQUd1OLC3aP4Tt
hh1pBqVE84vOi/6UKyRk3tbs5F/mSw/StV/N5k81MlvnAezAX59FEdpraJZ85UKK
NvzeYg8LUYUlcGmchpD+mrWPObxp1sSlV4tsnsJkB2IUhkx9QwVPc0l5AfvpKl66
NgTMJPrs+bLqg69Dz094DO45de1+W4l1gppnyWbosfAPqVk8JoMaP3BqLwhXe6Me
0wN2TlysSJm4MuMs6pshNopO2AwbnCbVIi0cMmDJjDfSzooA/UF2t00zyPeECz50
VsBbH2MuU2SC/aCCr/DlTEe3uePQJeY5EoP47+VKSI58R34an+mBRklZzR9yV6kj
1vY6HYPCPR9sOxIWUtP4JyGKHntfN6zRLpIYdgzCkjqByy8JdCjKOz8pj6MjWysr
FpDrxeBLDH5PekHQSfNkGC2E6/xCmKdWueAZRpCN2wr2cC1wT+J0F/jfeYPBFXnC
IXAKhUyU5vLGotW6bDY8LH32Y4qM59zmlYgfpSos+5AseYFOj0WCGA8Bttt6FQZQ
G9IflLMJwUdfRnVvuXq/kcIXO4JH33JqqTG8CzPLwsTiQqQ722aL9lnEET2lUgUn
pVQOCo2W+9g0um4/4lETskLzoE+IZfhOPryZPr0wqJ6zboBZL7pBiFJ9NhdMOJqR
EfiEkYcuh2iQygpiWroFpjZ9sWFUh7GJzcz2NaOzxxyOOzHOHtvA25ArM4UNYJDp
5b9GsVpkFGjDq2lINcLss4gexFhGaEhLEPhQl0trv+KeNWJs8OVjQa8AtExjMNl5
yLiHhRnHtAaf3QetOMYMNUx4GhgbIru4x7R+WdDckxlSFs2W2MD2QVV+ZGrm+MzR
Z6oohVDdPMVtoNHnxZB4XmR7MSdx9NII5sw7YiQZsQE0AAFVTMyo2fBp1t8yBOTi
g3MR6rp8Fz7OYs5EZCbOAfmFnjJawv33AAOLSm2I6Zb/nmwCr3R3UtALimXEqIms
WxiQMDyj+NBeBsuQ0+fgK8GfzWRrgalNeukk/bYatX3m5qcD8Xk+W/3NLynssl97
JNtbxqqYgtiNPKhC8u6SlZDZLP7ZT8IGv4XyEtGBmPL0J1tlPl2Q3HCKl7yCqnNN
KSTEq66BZh9WN11PYq7EyZYAEetkiMJQXuEOMQFwDNFCg0jiCo00SW1I+RGEMiGR
BCTYRxQ1InneJuXClh7CPQL0gJMctrxP6tBs5mDknOiI2Mf2m7SLKns1Y+zkD5AR
YXmA3RiDE1ANbljYzqSEwe8Eb2+zR1TBy7KZ8ahR3qne3t5XR73jcYWAYh955VH1
YA5lL0HD7RH8Et9uS/LRAPjYBcjbdSsEiQxZO+hSqe64zPj5TpOABxB7MtMePxTO
nAXZwKwm6JwfpVPFUvmEthtN5Hj5JxYrIONqFHsNvyzR8eX8SjwmC/5aWQmbJjkg
PwSwtpQaNVMsTEIxDq305r0sAvl9G+ZVmgen+9CagrFlgYMZWDXvLKeKmbqc5tlR
PzXqxQgXWXQRjQKNZTDAdOYP1+cca+tnpuQg6jCedUL/LtP2lkWvhMGLRmcqnR4N
5GvtLckwaLkb//TmQLGbVTwLaM/Y18Btw1BZBiYFPNOsMCkDpXftvOfCFfSthIqH
FntG/kNx65I5SHU8zlbv4zOwY7RfArxlTahwaHqpBNnQFKOWrW4eAULb65rgAMuu
jLxv/fhxdtlNXZvwY17v3/tsnFUlM5zabfPaz4GYXzqiRmamGiRnroRNhXr4pJsx
S84mvQOPWtrHbyCV3foozFC3yqD6AI2rqT9GwPc885/PEhggv/YmeCFSG/UOARnT
CgRiYuAr7L8Xfe/f2vNtevp4wKtOgMD3HtELO198xSc=
//pragma protect end_data_block
//pragma protect digest_block
ksK2i/B3gZT2AqWXl5Jy5EGCxnM=
//pragma protect end_digest_block
//pragma protect end_protected
