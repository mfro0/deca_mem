// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:41:07 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lnrOVimJ+YYoRqrc/PpFs/TYtoQLbyW0qwMTPz+PXoeuV3+GvPKw+XKFHQATOv+z
QAXqxFy8G/s+hj30EcQo8gf2BQOJlrXIaPpmyvNoL5t1WbChNhaUFIJLwsbKdUEr
oRnbFIyR2UFAowrioMXmqAeg924TcnPNuKWGRppWzXg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31984)
aUZKz/lckBjc6tp8GkJvcwr3IgWCOGInFwyGdYnbceGIH1/eHYZ6dfhviiOtG+t2
v1J510dFlfb9lQ3zKiEAYu+AD2X4ClPNvtzocnJtpIBC8zd/J3HkDF21PApo6HKZ
uA/4Hcrf8PG7BlIPWVs42j2dwMaddOZrA+aA7N19ZHGRV/t8UleUngoRXV+0rLf3
t3DX+9xoHhc8pwTSx5up42AOJ1uSgiHK6THi6miVBP74bsSRrzemGv6PpHwUbAk+
CoTWM9RdieIO+CCbUvv40QIoLPqRsqI2cS9LaFfmvy/wwOOnR3uHtG53+F+rvSkA
l0rfTTcHn+6ak4ohbbzeENqkAdetmXpgmwMfKND0LBBEujL3bBCq7kQ2Dza+4Hei
beDThSYHl08MPmITnPpaAnU8rcg82llQPAeG0PKg6w6B1Sz5y0FTyLOPc2RrbIP3
TvclUMMP4QehJktEZ5VNgJhgkWaku16jboDRcS4HI1sEQMmZ+4aDg52bbSI6tAGl
AMtssn8NJSOBSxlbWyKI5r+i+FaR0DxCcJdVCjBKZEpoWhh4lxSFDrnyS/bXnqdW
aVXnNV+ete6r5FWLjWOZWSYGXW7wslMOZKnLtb21n+u24Zll1DuPOjFvKAWzg/tO
RuvkmDVHF9mRjDpOUgkhTopuysh5fqNFqpZrEIewQd2rF87+XWxPnuqlOPMZ5+4R
gQN99z8KErD537NVTbfXUcrY5HdRB2JloBTeXZEoyqzZPe4jCqgm9wiz4FNJk441
STjtR15HQctlQWCpwvJTv7Ty4IoeNpuCXHNwnPxi9z5ZfhDtXPE2+kcEjxNCJoIS
IPtKvnOroVu07NcC9/DLZJptOt618pro8eFEeytzMyJ0UB1tclXDJwoeo4qFSWAa
EgaqgGafwZ9zzC7jEIyNDl3GjRoE0YjSdpJw1ztcZZ759Yxz9zeol/YRgoHkdU3M
s9pZXr9LjO5ft4v9kdvnjUPRUXXnEksL3JTTL+jrvCIKw+Cb/EMI2roG8Z1sY3A6
hL3oRGTAgFvV+n4GHy2yEMOldd2G/Znd1h2JMR9u20IYEwzIi57uMNKVhYsW/tI/
XnoNcgWC0hq0cVW1e59sQNRAN2dlUdOxdpv6t/HHLy58xONU7BKqtEEERroIcPmh
rvm6dpb32LNnV9jyMShsRQrbmKlSDT6piMQqI9LK6VBrWBG0/9r4/JOsaj52rWMQ
EFrbVB4TSYP1sv2HaN2CXMOWuqLfpIdPs/CHGuUbjdIK1iZNfSmnyUytqxMRpWCo
kZI+41r2HxeyljMzaFx0fynfWwyWCjW2PqtaaavNqedwlpr8+yjf6u71iSFETluV
B403jFtEffTlGkNH7zGoHiPqRU+jB6AQxPfJccuFXlLpaoELmlh+adbcC8gTSidB
4AIU74fsFVAfhoMv5xbUtBorM+/j6NBo4SyL4HWkmgDooY04jN7OnqCu//xn7Hcj
cuuR7I6o7tGK9bcOf9W22CQbSq52ZhggjaWucwJBDCguTmsesQ7ulTPYcfV06qq6
X2LfhvyQ2R8r+Jmpzow1i5c8xNpDTvAl1xHPTaSAlhRJCNsnekn0FDY9CxpvytSz
PjQ2XutmVkZ1ZtvfxQey/0/iZnR49PjS0MGHpP2nl7vTW6vsKCeroONt68GI4ozV
ecZ/SCKyG0gD0g1YbX2q6E4MuNXEBkSnilA2DcKjsbsvQL9hA0a7f8LtM5MEVWkQ
wOmp+q64RAr5Cp//A0c+9iVzeBGlRwew5nL7NszOUzZRb7ga0S+ua6t8aS2os1W6
NjE2k1/f1qX4ILnDFpinr1SJQSTwQld8rJK8Wr8XPtnj2lX5SjdbZHXIpGfBD2Tz
X+Qjoz1kLORR8KK6YZkqG2ZSi3K7yAPsj1y6kkmkxizY/m4u87egq+DB4TXGGUtj
QxXWgUkk4YiHmJMqz8LdqZOUsQYEySU6T7JSxlJHtEA92p/a4wuNGvOh5oyPhwSb
K9XRkKjxogNhtkLgz1/u181nDZcQLZF8dC1ae+KQJlZkkkoAuAxHZ01PtDFWmIpe
3yfau4jbtdoUuPRDH0knkIVDEhl7IOx3hEEMWqwloUoDd8uZ+AAoLJtnF3w8eB1Q
TgJWXaX5zJFJznVU7uhj6iBMb8IXNlhKubW0ncC5CsALqNJpqbRAzIacz/wjlioN
FyzQ6PHAZxVe41a9+Hh3R3F5KLaWi2HWvX9+okwrstxIK3wO1I7R+JxYoPZaW+VD
s1STU+qyToFcc3vXwNPtGL5NJIXvdU7rlrfHKcGPPt1XpRTWwxlsPQCWpyIk44LE
KsTc52dHyuZup7cWyAaDxxCx/aeZ4jAl5i0ornynzv5teNRdgR38v6vTgrOf4ZQh
F6rgswpCXJS9JY/oARvVw4sEtmTnh5HE9waErt6GuhJEi/YSrjG5JCZmt4PdXtf+
yTIR2ZvGEXFQJxwQ8Kl722840Xx9zbaxfAzE1XhLNAJ/OKePdaqF2waTcL1PXDPS
rzZ//qCDCuipIALjLR33oz+6RjGcrM8yj0GLrZk4npOV4q7Fq5Ltr4ZTVN1hZEuM
MacJTNu9B8f5Q8QaNj32ba7oW7c1UqZVyDgMnhPKM+1XL3pSGhya+xeiKg148ZEk
YK8ojW+aqMvGBJHYzpl0pSTTnPwZSaeDMnll5V1VdFE9Ywh/uFOiCFbS2SwduO09
Pbgm4ht/AI3qiQWyqp3pHbfDUG4FxiC9x98ZBBGBbiZF9k3QXFUcGh5X4SNA6emG
SeZpwGmxHLFJWbCnQKNQ/9SfjJm460cenuvfVXDouVuaB6JZHgtUUodAFDs2//68
w+QW8sPc7rdhidCiMpkRcN/e0ISx4zrz31bH6uqeEs0B385lOIIiBpdXLloPKJXz
w84HrGTRkU8WyciP832tRs2FN94BJDHZrLF4R7rIq7NagpTMTxRDf37b6S844lq4
BX/29AIpgIMXjm959nIOYl4USlqLBu5N9ZHsZjHCB1U9SXAWA1VJWpEhmxYmGa0s
pE64GFUBjUT2du94J0HVXi2QYOxSrqBxw7Tbmvkzyv3dHx8OWrCNrDJQwH+UMAMQ
11tRSsu1tYAjA7FmOeWdaEpn/wudRzItXjzrfsxu3hbLxQkK8zx5Q0oktmLpQDbE
fp4qtJobnhOg9IOUphWAaPJJBiFaKsUJMFycluvmP01LBE2YcoNwgRPhc6+gefA/
guhDWM5xlhiJnJa6zRx7AO4YpjkSmhScgtrQVYtQUK17QfxzkNss4RC8KFXuy1ih
4QNbouG0x8goinSuDeMFKIT77N3m032L8oyljiXyjUE+2927K0yaQtNibULznNEv
NCc35M9ruoqg0ZFK6ucIcd4BygBi2HqbOkWVgrdflmj2kEldM8potsghll2pxbln
aNmDxXy/PdsNn7Yksc/tdEvWqQfCj31lA6uw+0BHrSau5Dueh/cjYImsbNRTNG2B
cJ/C+rL6Mh6rKMsuX+VcQJsBEBYIYNu2ZMwXkXNh5v69Im9LGNnv65BIah2Ky/Bm
MUEFlIDk9xU7afu/x6cLS9zDJGRqERfsSEOAKoRNGQlk7cKO0+d8Gabbtic/WwTA
4bDG2DTxg0dGT7K1bnvruEZX1+aUlHG4LrQz4z+ERQzgrTBFkb/eEReRqtTjdcMG
HrPMuyz9ejJZbYmFerTnbnauhhm50EOuqicc1Y2Jq/1QPTN8qrNWTzNGEf2mybNg
lHcY0Pk4zy1tszjFXtSV0l1jQoH0hI0JdhspZO18eRqa6m78W+tTPylp+jDpochO
C4GXIrmKtoCOA4scKmdxcRnGjDOzl5F/wt2EU8+2jhpP6YWuLd+I+8ttw3oi2Npl
IJrVHOCpsoR/IPfPMlol1EOI13LIc4oafmreykeySsoF/gu6yCmWz1rlMbpX13gm
DohnKgyu29XMIHN7EHnMeUylocsyngvd1JwX5ICoxlmpyTRJoy7xzZj5OdxnTE37
TTXaPte2Fmsr1kSTV0eCNsFHMctuKll30gd3HZafx8yHdKSQ1R+rvLojT6iY1jEu
DWufNUMGgH/uoGbE3dWr0bdiqAc+PW4oZn8kkJtD4OUq4XlYZxk5nLHYzG8dJH1L
9siCeNlVxX9h8Ol1mx5mSQ/M1oE3Qllu6fjHFvG47rNMGogIPLL/lhDXkmulsfPF
wlbZY393pOEtmZ/zqEkovCy5vJX/8tPTez1Hrsvf8K3gLgYovySHXjTeZuUflAcN
sqQ8PgiZdbon7Lfm27/ZrW30QooUr/OgYUEHRU/n87K3Xl5/ARcUW4hxHojaS/7/
qvlDWYAOZ7vTU4/vyprtdE9q3+KvnAUl8PBjOZpgHtY9gKBruTjxzvCvyDfw4L8c
8bd++AtLlPZa5Cz5MKEOXNtJAGZz/trLiEGSHAi4saOYHKDm7eXbx/mqP6UIcazO
pt4/dFsIQO54FJgduMeE1i+Zj8qIkYNeiI7ORhH7PCIuF5BHjzlUBFqKnSzOt4q3
sUNTSA32BeRQI5OJVQhV+upJCPhGyPWCJoHUovlogEpAGRYDhv9snIBM33XGWm0H
9AtaLp6g/LhFAAbRnhTMuDwww5GW/2aHbkNl0bbE0UcIjli80ySVNZ291Vl1dKO0
CDWtJNymz/eUY7kuYN78HLlD92+AGVVGyPowt/kkyP1QW/WzMWv+IMCkStrmp4As
kqY7UW9Gi5wOzbetaaxkxvpHRcxJT29KUlZEU7EIwnDaOe614BXG0TDR4Hm4OruO
vb7ylidf7Q29AZ12AoKPu5k/abUCahUNZQvp+tn4Oabt7kHTzQx5Z48hhXIbEwsJ
r7kgFuTEnm+7ThIA54tCm72SXrajgJLViJzSHNv3XfjPQBTvNyobQ08EKQBibY7W
+OHe125x67hmUWZUBd7j+GIsvX1Ak5lU/7BdF/AKdeaTBFMIzWbw8eq/Xy544eQt
4gtLuJAr8SdoEx3u3wWwV2Wn6jmGX6nke3nVLU4KNiY1nIpGN79WN48sXafcu1Zw
xXjcs2CSX6rgbgvREBu7eEGF8CD90+0O0nh9HpLmvuCdNDrrgRhKAyFXrh/rGTnb
6f5KLGP8dbM1g/tkVtp5gCyDhtVsmrnWLil3eewCRJMjo/uwbkwGFYpiK3LzeiB/
baCqtCucqqFPKdhB8XWqj+ChhtPMPdNE2JhD+1C4pPsGe4ZINrhPPtPblr5wLSlJ
6dfpXp+RkMavAXUo8i4zaNhgolLHPeAIIeXr+DJdHSXfG0nqTOSVkBoQ26O3JUGd
Hf7rJ9FjPr7JG0eZUWTaXVZq+QIW+LNdWxmSNs4RoqzeaVI7oI5MCvbs9f65AbpS
4k/CVD2UjC3HxKX84LvxyGi4yGqb5xwTGJHwrrEilyAVKtTUojVr9WrYu1hmWZwf
JszKgMRwCkIYggaqlFL0iuxUVQsQlnLLDXlTctVNNlMVW5sLoXoE2JxED61QRMMU
U6lo4IoSGtQy71pAq6x6IxpLolbure24AE97HdrJ5YDutX/zK/Y709cpD7ZLGZfJ
d1LTghhCmQ6CWL+YtMHaCUQ90SUDB5arXWb2iDcJhR0Sk0F8G0fyLrD5xi937e3O
XFrO5XB/XbCWgMqVd475J4Oy1FxCE81DuocMsmmwtuzoCItvzfiu5P864ECPpO7d
SfiNNwKu6LXhVhkXpX9LKLT5hKQmEOszNHaUtoIxm9qnGv/HC4v6qekmAEaPugJb
Y49TrbwO6dzNSjgX1fdAeLGDf1xxrqrG5kl5kYO/UKIW68jI2sYYuRhFu3kj/ZOb
FfGO5sFyipQdydUPJG+UjqpyeakiNn2ZMpo3Y49MJ28XG++JRYGpygpOT4lpixRo
9m/rmTgeThT7j6jsX1BtGseRX+axxcbli3e1d+kFM+evQsTnrnWchfSfmveKXaxG
Kay791xHJubsxZUpjCOr53J+xAgArfLiqhuBTPsnIjeP5Au9soPyxR5RkDiVO63F
I1Ma/XCFz3qBXLBKPqO3RN4DIsiUZGM60953dH5uRVRm/xiX3Pt8wk0x/ZMLHjgW
VSBMbBYw5QeSOAREXoubL5N7qAXshY20uC1EiW2xIvcyrNVUZ+u8Z7KkoU4ZUklV
NfFdFvsgMVesHlmGiKJgmEWl62FUqAtb5/8YK2KuawvmxNeV7RQliPf7jITmYIVi
8zyrEAb+RM+vGQVapxzcGjGU+R7hdLKHUAoYX9OFCZH+GQYGBgq/97vzVKF/iuqs
a9xQQWQcIbeFCAi5dDC0oYnmfsLTqsiPzLq1KQEmuPjNyMGX9SQM4EwUS18DZwvH
H0Cn6w3SVqcUwmcFdgoWJBdh6pK2lGaHEEFO9+iUJrPZASYdyIC4JbDMold5FC/2
5txqu58x7TZB7KwPSqMIgsH7gamVl5SdWhS6V3h2vwfBuhJJxVtwqTK5SOf8VnXy
4/lAz235EwFOqAb/t6N+f3/iuIZMrBtgTDecvtIsUbEmI/p7buH+XSVt1RGEG73W
ZCHDZkhwDeEO1kXT8Qkj4SC4MirmTfuJPSlE7arnmYLxbytW+RFgbyqkHImfp7Pq
aA36stQmPbCJpDS37Sn1EXHTzLsg8ZJ2DbullQYzrUU6HSeIm1DmVJ+jSlSOaOYz
7GF5ZmBK9jBoOg4scq5c0FLJHwEYiOQ+Ix6BsooPjOIegUGHL4q42TNsTRWPy2/z
IwJEog4KfmrDopD4GoQ23whVzXXrg6t17jCRbYT2/aGItzg3/GQfYtUyImBe4DSC
aET8EhO+IKqgfFVpM45TPttlFurbIzftSaNutYQmgIJutPdCFW+7ZAp5A7+HMOwC
dDo03R0LyJwZ+9/Et+uN7NDeQJGhMQFakVxR0tos0s0EvfxmA40+/slR/1qepHiI
Gl8pwte2v7dkAE0UvGAFGJE3vOHzYSvzaitt2MoMkYZnyuFt5fK3cd8xbEaIVeA1
t3fBhd+AWI4knl+hO4vE79agOke5Tar1VfjCQnT+XELgk2AMzh6iMTXQAPHkbt7j
PYgkxUv89GuYEkqem7RQYQnnr1+ovOOFhGAX+A++K03o+rpH9AA1YxtG1kcihIDt
EEx0XHg4gDYQ/oSrx58c8o/HI+ihU/ANUUu/qJUTf3qDTWt0AVz6lT5x3qNS0AP/
8A/LWty8lt22wpYNn/jJbo74Lcds/YUayZKWTVBgbqnh0uyKqTR3U32VQ5mr+08m
k3dEAtMElKeDl63YGmukr1MTq0NM0xX8pUSEs/L5674LUxG/glF/r49IuaNnRxu0
SPVbZ0rmpvuxsW5v2EF9mmLkBuoVJpbk5hvlUCgzTzf/SxlkYIWSHtDmnxAt4e/K
W43N7DljQj7gL52Sxg6c2xGqijz6oA6LpMNA1HnWxNYxigplzNubxU+4aYuJf+4d
nraHxMtyj+RiWUwav4fypExdDNioru/mLEP6JvCY4zh1k1j/cHxPDaMGJgvINdAs
xdBUg505yo28fEOD7xhTdM0h2yc54Wjl1337RXOvU1IYHw3tP2ClohgPnEDVF8WB
/3EzbxqgDxK1EMV5aa+bHcYeJSCtBI+bBRe6zMp+KGN1zsMg0O3YsfctsxPHeACs
H+jihqTn2TwH8eoX3o6Qj5XwjH6sM18bCEm9i8eFDEdrf/5grSYlyYTdm3ZqmgjD
S75/3o2lfsbIjZHiv5Z4WTTjogzoe4vl1+7KziFZ7nB9d9M3vbyWMLqm6aW6ILd+
TamPQT8Nxo4SyVzxNJoRkUdf+zkrgXFwZY0VeuBbRwddZe1N45UzKyUTjL4qfbVq
Rat7zF93q3t5qFAI8p0OPkFE/dLVS0JCoeAKZubgl5jYnzd5RiKpBbN8PWYUr+TS
QHO1BLCp9QDSZIDphg0om84M/dQ4o6jSOrhGB1s7Lg7hTljerC7i0DqmrDLv1wTQ
fVcYziTnqqZSGhKQNK0r+l9pnMvdMvUAS8rOpNP5nkTJFpR2M1i7H1D8/jVWeTK1
L4LjoVDDucprHJ3opuxjtuMUPZNWSqT2r6CLmntzIG9XeH9OzbA7VgcYf0DAsJOn
9/2G4+biuZ1UqeeeIqkUg/nOl7kEhh4x7evBoRrn1CiAE3J4awFcVikSp8uF3+B7
1lzeTBqlIdlvP7IC+61W5yrwaQZrI32PBcV9fxioaLTPQkGJIi3Oz762Xav5fE/K
cTU4BbLpA5HnfXFItbHXUxh1jm75GxXZa+Ap3oDmhXFZZse/vVIiFKtPEStysxoD
H6sV46bDJjRwWd7Ob+fpdwyk3v4r7DZZjWSi0K2onrdVnVKfxIhwRKG+x22bo4V8
sxPgUZm4tHFOAWiYzLj/0b/YojX/wYHZIwtek+MpmMzldzoiZbAORA15QW56ig5u
s9ZBEtNn2z/34vHafkfCnWGqX+isNXHdYLDR/yUNG7RMKV09ICX+qDa39Ta/tbDq
bxBfeaRzByXwn1u+shXknHipn5jGx+ZCrDeI93Uj79xSM3zJEfLnAmjqNSsk4+by
9UU7qReBVkwxJGbV9i2bMSwvvYhKEFMsf3W4z06nZ8AHR8ZOe486Jx1N80Eac1+j
9tGr0g7w405WFUaFY+0UrGV2HL+dY9Tt8ZL+C+SO0zJj54BUyWKDHgb+bfXolkpN
jYdrNXprULNVIzORlJJpyUuxT8q/v0HCoJehyblQKiJqjpBQ0TMS07HdgO/mJTR2
8QQzaob7JxYjTAd36Wbq4GOqAXIcX+AC63mo9kdmbg8+3lJ8Wx+dEwLry9OSUPXd
5alc7MqO5ADqwx+y62l60flL6jPc/iioC3Mhw6SClPlKiWPdILXVksUPJDrRJKxX
nTwTcBuv2wOuIIjCpchZkY59duChkgCLJAg+YO5d6Etl7ca9deqZ9SedWr2jtJvY
X+THeieVdBgTAScqJANsV2WEm6g9psGeL/KzHjPfRyjTiEmIGCQL1OSZ0iaGMWuw
8VrmIBXv3w6BhVFwoDMMgcTJLpF6XHKJ7tWcw7QC7JxkTqUhvmOzanniH++gPpNY
MvqydgH4EOpm8/4VKjxxY5qvR11rGYqqd47zGd8w97FQEOPpQAVZ8tWki8y/7gTP
EnnPfKNBnbkCEWYd/0tV89qF30WuRZSo5AWucYEuSFOQIp8QiozH7XLQVfkyY41N
B2L8qZ7w3Y8unFe+Q/LAl0B6QyUNlHncfuhLdOxUMXVurNG6AGUx/2z/y/oE+EL8
yNSc6DUXkUDr/YCNXLG/WoIjlVStQ+iayA0HyPYQvV3Jwetv68hvZPbclkoPtNgP
Ipe2ujZrDwCCQxFyvFs0ERa6B962Q9vxj5jAb+OX8qtOluphBW7Wvd0xguR39SlE
SV6DXIG28keQQm4zyrl/YUWT3zCpZp129WbfYbKsXoF4rU1js4SeO8wAZ/f2yz/Y
/PuhorIWGqhZk84F44t5B1Q5G2slL8sNCY/So85uBsum2LQj2S9EnbJJ6Bwf+haB
D3f2XzsM2oZ6TGaeIWx4Ycznt6ffUrsIOT7V7IP0EHbhceT0VVhxSzHEiRNVLfTw
6sFm+9fJUBVy/3nJqaOQbEjYg7FExJ5cMlnqEw2wkxnGHN8eYU/T6mWkrA/E0tmo
attbL7qhbIiA+6OsCTZtCmxrinoPb5cg9uVYvLwtOJIkwp4sKK3GNkVbUy+Yvlfh
b1f+P3Xt2qjCqXVzWPfW8vzoQFUP4giJIxiY+iwdme7AYf9p3awaTO0/ibUiewXw
IwL2qzZSRBpT4TF1AoAyYU4cpNPU1ikc0+rnIDsMgdUq6qHBBGSDwdv04Blwj5B7
/8uKyxBe90kOjDr67QzCl7WDJYbjqcOOazNlpydR9p2pa7ht9pSbqCOKvy1iVI1j
7mHQd7iK1I2e3SwhIOcfqEtl9Cx0AHWwlhJr2ztMh/THEkEDRCreP5iTuR07Y8nW
o0Ou3F7dhks47npSbqjLYaObwjscwaVyndhLHDJFZu1yHaMB93UTjTTgEG2VCyOO
NmwEzoH7yni1yKwAXFVXUgUd9tT6th24fQ+lgewyUoQndusEIW3RlulLdUqsGSdz
A76Raq8BWVw5ZPai+8EHs3L21ZTAQ6+fL+LKwXIpz3MvoLKraKH+HzW1WmMlMn+v
KMQo1zDUCWAGokCsgM8PG1quLu5IKZvWDQ2mA3ei54nvnIB7/gUel7pG/h1NXs++
8hK0jVIGKjdll/3NiU178fRC1RkkbqeJVn7UZhBIEawwORnZnHLxR7fScKUXuvu1
Q1w4cjRPQHzZZ5cHnsOgW5L3NFHToGQsKQDca+xV4fHsZssMqtINqrMw692q8ELp
JT5wkrAyOS+aA2AIoCYvBZhvhcqlP8BhvuNXzcQtf3z4w8o7GWmDfPvTOsTchj5Q
9Gj4wV7/N5I4yYulFRIYe7QjxTy/3rhsgAAOYEVP8zHwsC6i9iyvatB8KUsrSXA5
y/zcVToSod34XromcKYt2fGluGGinyksubk8Wc+Kx2b4YSzXkHHaQcGq0O8GRxYh
AsDCW8VZTjIX/FzPtkOYMKhcqCuRmv202vmt2lbEG5E/hJGm5lanOkLKbzHCaDT5
JH5LEMEDCQSWhJUqaOegt7Lsd2reNwYhIpEQk/30L4/25frmG4f8Nn1iQszKrwK9
PMHyGYHWkGP/BAaeC4Wyuwc61ivP6/012Oep7u/6HrOvDGnWhcT8FVpWdp7IAaMr
R/ltN/L1Fzw/Ttt0zwSQKksFrCdV+wIK5WkSi0QquceJeUWOTttu/JfJo4Aa8WMZ
RUZsbkA+FIXHXCmyJpfpnhtYnQ5gSpPurmIGt+bCm2CUa+moLjHxNWnusg2x0zqP
437WKgS+Wp/ML+lYhByjrZauLqe4l2HanjL/lnpW1YoR4srOFtqpNYM9TvPdHHEw
UvL2/jLqrJKgtI+553OWLC2vTFhpsh/wiCwKf/4N0M8ev9ZyQ7IFJOZBTzn1amX7
hEFeYQvzLmGWCys3kEClMATLSpRUFBLsTeljniT4ffL0c7Vv2Oo+n0enJ1wbJ+W3
irZih3ci2ucXKgluymsg9iZOQaUKh29kna5yAYArlch9f+kBVw7WJc1EesuL6Gal
6rvk5wSRoxCUWMYMurFsJ5WBtcQH8N4R6E9k0qRpLaNI7cYqojC/FWtmXHjKqF2Y
moK0/wv8gyXuApKk8w3F78xyFMXaQ2k7Y4p+dTpWR1RN2Nhhjv/ubIV4Bj/59GiE
8CQGJPuGhiWzYznWVvU6za60p86EvackmsgKJ8/Wc2NbllG+vwyAE20911gzjCwb
bTp0KjmGFxAY3xZYI4Z1x0axFMi8WIbLtIGTt/EDt79oT1ESF3/dUKfHfD2+c6MM
ZOt7rjpa+R2KpayRwSRic2eW247H2ibEYZjjv9/4v0NYRbnn5OWj5egZX5FhEswR
nTbmYGuKq4DgaRoSC7+17ZSwC7vRPj7ZmstVqxyvyUiGplnFlBFWWvosCjsoSx89
006tGc7FjqqPvynPYffx2qm32WLPKHeLZ7CsYZ7wyOyGsZiN3x5GctgICMnf+qmO
PYuN0XVDiZVCc06RfwL4V8t2X1OJqmVS4QoU/s3lCtyEQohlv+dqGmLi+K2xU8DB
/szaRtMaHBvA33qb8nDXj8TQqlIRK5WG7yPk32T7vf23CnsZoEPNxVrt9Vpul7Cz
/Fd7sBXtB8cgbnH56+nnEfPakpkZR9VYnO0AxqZ6qS4dMBjmj1RkskLNA2uZGeLY
LQoEOCJ59ID3L/e9bnyQ02TNzuS4MH6NnFfsw02CjhdzXiN1YCLi7ku6hm5sj04D
f4K3XtusNvu4om4e9hRIe3YNqrB45Rg4YlLwTcxzuge5MRw4z9CvNyDbIj3SMZb3
5lbWbSrT27jqYC+whRFlEw5bFaj6z8uf3Nk12gY+ygExnxVaj9RIlGxxEUScxdlu
PSQjfuStjlJs0cCNyy+lu/phg0UocHEgbMDTKdO1iGLsjWXnE7FHgNal8HYW299G
ykUSoPi/YLvJjoTVF4cDILI2o/NFev5/S53dXchdHOJkXUpeAfB3Y5GRZg7ZHr2v
wiRUV3ZeHLVtcmgrtW0mvjiaMAUxF/0pM8JaPyURPFQa9PYgB5xwLfzvqJJOxPYH
YNU55sp5jXL4ahDYjNup9K9YkdexrVUgWTFkHCwLUJquTBaGILfGI0Td19gUWZTK
sk0PpRwZwESI5RUG2oj8MtjHgbCsr/DulCveMxySFXM58E2ZhqROJPtdW/zUENc5
9anjj24UqLu6eqKKMEyzhjPhmbIh7vQkzAg/ntAAqKVy/2wD3y21XQQ1lzI6uQt3
IkDeRCO8f5pLX2/EWvebQjViE++PS4UtkWYxZdG0uC+Rt+AZEWBf59xWdbNM8sTb
Q07Wl6IgAlqTZKXu2mxNe/i3QC2i8bMVs1hbHUUA3GcYuXVSHiZIGndJ/3jLX/Xw
3WauMEMPgzpUp3WQfvvvD8wiHwJ8GC2VDW5TAa9pwiu7Av8VtMaV+tKkR3XkX+Ik
hWdsGMfCVAAiGRuxS/mYe08a6Ewm3sVdhaqM3ZrF6yToVGRuX+hlBw/5SPstrscm
YnJ88LDPRNKIhaHhdEXdF/Nlv9r4pmm97Q3w01E4vWWMbNt85z4ePRc1Y5mdvn6q
5OshZ++vH5x7S+W9dnz3IRPK4OBqrJvMQAKonuvO/WFqJ2YeO7HeYzVQjTSFjJ2A
sFTe4lsAPat4HQzT0QNz+6fZs0CexY6FAGRJE+LiF+8uOkVPtbFV16o8ggGalm05
uXg8EgtzFGX6Fy2OeAfFr8PUzooLPfKk81VKvqCwBJoc/B/mbnMpsq1cagBkgcs5
oUFv6dPlZBOPPt6epHvXPUu8RV+t+XRKRSONxU+HWwCd9SBw5C1hWTMsX3NAEbpv
Bc8AgYZrZZkTcVg4MfAFKRvizFv/ljgvO4AkpK95mYegsGlPC0xpylYIp6zrynJI
KATSXx72miShcTkS69shdzciW1TTZ4ck/bJqw0h+pTodDBFa7vsazSvFU4ECUPNb
qZluHtKK7+c43jjmftOOsbGxyN+A6WKv+PUo5af+GLjumQ0BtSTTY5CZC5cRsPd8
or7DkKqbpsnHSG0UuSBGwZlopRAz15EPzgejm+sbMoSlWcIYL797Xe2LA6GfQbxS
QPIVXoSvSlw7N/FWlvMz7zP9XMxUbrTr18932Jqgi2idmZzcpWYXAWHrwgoYs+es
S8c5pi/kI89aUUhb/syFHTnHymEYu9WX73MxL1CgZ5qN+yrj08Ka1lhH5TZZG+FD
b/5XoPY1Tx/Y+gT4HGyBsmsbXDxxEBWinXi+DlTwkbmR3B8LQMUIF2mtWfR/e+CJ
YhWtE+zFZNLfwn9h0oJvybSvpGMbPGPsZu+aDl9XfaKLkkE9PvDf3/qV3vXAAxTr
NNMHwQMra2033SbLVwJKvfTRKBNRuk10mG8C+85gTrk1YEED/UbJgnRF4t74RzRI
GotPfSeotmsm/pVBK8aIBm91xUZvBbw76rrAS2E+PntUC3x6sHrd1VUsNM7+F/JH
QI2dZHNefJs6QFAmSk9yBbRDuLp6SXNYRCKVAVFXmHq3khB70cliIk3jSf2Wka0i
5XzV9c8rIN6tbyvcR2rRLqiI2EJspla3BfV6t5M8QIgxp69KmTgb7wdCqe6ZsohG
OG2I0I1ZWatGkt1e5eqlznsPH4sswT/oRlk0/GenNKtVNpfQyTCxDkEe2K8z3R74
nkvWK4+qTJOintZ7VP9AAwHdNOeJJskNqOVIrgTlwamMjDd4MQVMd0NyQoFhj6A/
MUCNMHOUA3kZzzm/lAdVJZ0NVgIh9J0RWxL5TqcWNuBNrAkX0hKArFBYZcp1DtnV
4m6FNXMCOrTwTViLz89UhDCO/oxdG1z3jzMEPTmx2QLa2AsmVLH3/n1/MleBQ1Sq
P3OQ36AgwXyJ3p5CHDQZENNxisdojekks5JQfirQr72hjkIvrS8gR7SQK0Zzcsmk
QPA5oCLiLedjgEvjIA+o7vQidKBfQGlTST11tyv5ttIFVhIL1j9FhhuK8BXWFWIC
rcuIEd0Gv28VGqf2HcUMtxLMLJo1E1unI8LNSyigE1NL6dEEd80Gkcg2DmL7xv0o
PHyH19OKy9KXi8ywnsLKItQ9BiUnhTxPGH102UhEY59tlsc5s9lQR4EtZtta0OPc
7tS0bvL8E41zOT5dL0hbTo3GW4gbxpXAny9rqzr3n+yOM/mIPB2sFCRILLRB/3bz
eU5AN4vStaUXuP8DhXXtj+DqKl7XJlVFJRBWUi7nAy/CZXZpA+U8CKw7WWdinEx8
+ymYDkhZtzrm6eLvO0+yd3ImAm1YpclxKHV8GxHmQIMvFkCnOTYy4/I5yoQt4uS9
gizHb/94u1vQlibQybCv2DxQ7bv/yAEw1ll2/XXtsNz58QSSGuhj3PaSx462gj/7
y7j3aH4v1nvcKLTVmp57ev+2x7F8VnApdl8cWG87/deF9wnTNvGgf//rl6pThfP8
h3uczm4EaAaeb2bOE68bAovkklNIGoiZQLYKMKTK1mIBC3m81s4og8A54vU4uhHj
+6yM0JojcJm13QyYTQljbRNU9LCHBeKOakIy5Kte4oOSXCaNH+Or6gib7tO1fX/w
oQsSSOuQAP/no1rVEqIh6e/u58O71fp55dYCXk6/Tr7C6gfpSGbJPlj+HNhryYtC
4jYVYOx3szGrwtvhGwwdcWIkB20Kv4JnwIEjxtSIDtmXM5f9q9icYl4r+fToV8VF
OpjpUEOIKBNWYPKoC9u5+46S/E1RsyTHyuF2VwWmQxYvW+8l0BZ6UFrj8zxfWTCg
/kNREX7teeBQyg8RadyqY+mbbPqN+aX+AdtNKqATCnI74I6G4+x1jkz3pyWEUysr
fy41lqU+e/st9P9tjUjdlZw9tnQYaxMVsul1RLCaDKZ+adJghRmosJeoaabHeyf1
lgQ7etHn0qJer7sqkQKU1NIIG0XNARPf38ld3CZ2ZkCZ383TGQaq5tj1bqU43xWe
Lm/EJsZSQLhA0g6XoUDRcQ3WStO7JrBwS4qDWJH/tkKbL6WnkZ42hx6ChrzpY6fn
VF0sOLhvWaa5IVrpJ9dbDy3fMEUZwY87x4JifuP0mGRBdK+8FYRfkx/tGELiEnM1
P9k9F2iOx5nrE0RQ1kqRsITX1+lJR4o3yhSEC9r1A0tmJ0usvEfDfRsc1Zi4dWOa
2IF04csh7nRkiPtXJ6icV1hhE5UQuDDjQP1wxAJk0ZdxhWPNOY1kEVjW3TZ9Venq
sjf8TnfQ7/ca0W2Lm9YNQ3gazpwQcljaqAVxfVfkOLk749nYGP/34PSb5Q2GsBYL
GLZ5Ce7Y0oHhmXArzRc111EK76Zcw9iL5i2KX5Ec5xCYMnrK3FcaRhePUD/y9WpP
svnyfH63ot/pL39eRCtB4abkkI2CHoi0rvggdiY4IWJjlxZnBF11cT20ufsRZLH3
p5tMkDVq0LvvE91S9Qdwml3q3yl+IrhbxbdHyQr388IxWtSBdVQA7e/Hz28qM3hh
DUhGjzYWvlTCacOA2vCSFfLL5lJFaEvOn0cfpLzEkUvsGVZbAVkBRKUw7rVc4w/n
58gm0VB3v7C95L4e0Q042rL80kg3zbZTYVc6IHbkNMugRw2A4IHaB+D5no+A3kMS
/PR2ezxfYJQJChQMiEDDLAyobaqqBVxWKDomMeEiBndyvu1koHeufZtdV+oEnCJv
PcQVj/H+q2ofxYRpaoYM4EoR+dgZGgE8RL6SFVoHkv/WbGMb8LAZ/gc8Owu1Flce
8Z2qf05Tssz3hFZn3FDEOUgfwRTmThE6lb8lp+ZN4HFt5a+WZp5yAurhTF5VClSI
G1asAK7vNYLkUN6jA7IQIk3IqnsjBa2IvFp6gAM86aGxuWf7HNa27/+WjfngChYC
jiLhFHB0QdfzJv38AiG972evS7RnwBHdemocodrGnCGQjwHQ9e9o5mqiRHaHUOlg
x4MoRag4r19VXWeiM354NveTU7YBvGF6PKeGuNf+I/g3Whr5riadMfXaq5CwUYDj
uCAoR+9yo1J4k2hmzS9+hl44W18V2FLRxX0jYAMTWQfDA398WzDzKoS9lOHYCwU3
CBYiG88AYV6PbfmQHeKkp9knezb+eg7UcjAVnOEwMebUaPbwy0XsBvnFhLTm4OxE
e20qV0hMuYX0riAksaY+K8Fi13aJAKWGENE1ScyH0bRXMR+JQUeqZPqBwotsH2he
7Q+VT/atTsJoa6VVszxG+TUAow9ri5qYHVt9D8Pgrrb8EzANlYSPCPmnX2ZQfL6Q
+ZTkIl5kwzUiFtDQNcOuFNRO4nISRLhopnxZbCbcVSCH/cQp6rZ3Gmh+l18Mosoy
pSFKSKSnWxJOtJpKk89e2iVnW+kA9128X3PqYGUuZyupgFrBoW4Toa1rsBmv1Je4
hm2PV1GVSEvKW8ZTJgz/UBpP3eUG4s6t9FP66LOL+Lu+CNxmdIHywkyKMCYEJWTO
M+eK44M5VNNpoI7PBLt2RuLqGnKWXRMYW3zTAdZTlN6xFGTDwAin1YphUXqr9MxB
ZoAVhlnp5AgNAdq9e9Q2X10W861httg7BHKPV2eeEsrjzRQFQ+D+m2ki71cAmmw8
beHt+jw9uQf3Ys8HZDOz8Z+YE023FUg7fme1arRD9B9ci3e+O2sVvwdUquorHC3V
vBFrLxDRw/fH7pvUVMNoovBBBNRBs4Vgw/djG1zHcuIsqDbkG3V7+9i4ybrUQmnY
3QR/Ue4OQlwqhWEVDM0V1aGQh3Yf/73jip3Zk/jaPNvIZpVhi3JO/vMIHrjQDQFT
pl8P4MCRO7m8NIzhVso21yImECUfHy67pmKxm3cDhsrciv+X9AmHzbsFLXNo2jNm
QUjymH7Or3diSGj5OySLlNI9PsAK8Q3DqSuA3Dj2vqO4IEsIY2S7CHWCEqGLeq3l
6s2hTcxgo7flfrkp9nSAZE2U3r/CRKp9AyOg7COJwu48xUwOPwqbkXk4Sqs0Rxli
o0mu311WpJa6HKqGAsvh7IVwyKtGDU7dO2f5zqV1Vb8Q8toT7BTkVrH0i1WLSGak
k5vzzUUClCRRyyPJad8CMdcoiOfi+N0SeYTy1nRyJLDt59t5u8+odVjagYh0zjLT
SRsbXbgKVBz+ecno4KJwbVSwFTOT85NwaBqRSAg5jijrwtKavN6YmSM3sduIqUpb
seOgMskx3Pt/NusMqYO1Ej7RZa5klMSITqX2ODx+oP2rfADjwQawz8u2GHn4PzGP
hAefY1Hh35vqmlAzquSxLpO77xDoUD0AftbF6vOxpJHwHaP45XwvjgeYo7CsD5hT
EINgpGM6lbFfAVYYTuK/LE2sX7MNYmptLRZJ11EbF8S162WCNqEe9ZuFVRajQRgv
LEpqq+0EknAKzsE3vqK0YIfNVmYQv0KpRM15TzH6w2X50NF1D5LaKVNznteyIK+w
uVBf4JZWaeJF4KGpyHceWtA6guvEu2bpW60AgegoD+kM7G7lIj7QP5W9ay+QeyK5
J1K7KNNtxgr8rHaLyMDRAu3rMUn0aHKfgTkXGbmIGnSr7RJzF6M+MZOaED97Stge
/uYv5ApIzKKcYF89GrND0XA+f2NCHWIbm+MJECFFEMitz2MU+E5OKkRRWSJEAst6
kDMxOAIoJvFcwZfOqQGS7YzZ/hoskcA7LpmKtX3ESx1nq+jDfviIJbb+0J1hXHAj
s4gih3+5pHjD/R8qHGNhsEzPAwoKJsV8TwZNzUj+T/SJt6HtooU+0jZD9RHI9WkI
Wc/sNv6yf/gt3TTZ3pdVWg9gd19PsR3Hmu3OH/gf50NuTP8+PFxtzPSV2NrWE9Ac
klXFG8nbDfyBRrnvNaMrYb5DH++jcTfXHarY+MrJ1Huj3UThDTl0D0WfCYW9jHWi
dGDxoBB7iQMED7Wy7DvwQJW3E4kAnuDt9TgSbeqJwMrY3UfTTsDb/YYixWaoDr4t
bte4+BhE3cYMIxItp3/Ky9LyZxEKhSzIl6XShQSurXKM389KwpNMgGD4u2v9wr71
f509e5lgQByRy2Py7WYjPFVZIHnNDpLhdeM+ja6hFPiLKkcq1RhCoLp8G3YNnJzL
kUxhu0puc3RtET4XvJHEoOhdMOPOW3236FlctqXmR6DA9GImsJL0aA1YobFi+uM3
Vbnf5HbdDsz37yRG3KbVWgoOuAFDnyve+LV4+zzgHQ0g6Zl+ZtjfbZoseRj327jv
a1dfuXkbIyRBD8Y/o1wQwOBAovxKwGPsu2V4c/iqpAJxFeYQ7zXFMmYJcEzBUDGS
J2AYgdaXakK1Bc2miSL5/RQHc0yhEV8ylLTIOATUgGtrhNrteSlbg+qTjrRZIPas
sV6FujhFQ0UZcaiaTjQP5MeRSd9n4YnRNs1SzYNaWYOPSzp89ZMKX6kCjEet+cNA
lNmm1AaPM/Grf+5ZBJ82NOgibaZHYlain8biaG8fnf1bV4qmtZ7s5b3c9nzUBF9p
5HMlkmLX9WM7mVE62Gwk3Vd7yybtUQhh4CMm4l+LgbsErwfe+goz+WEIa2E86StU
kqFI2oWd4BFYhn007y0rpzAOz77CZjApA9aT1tvwEp3k1qBrq9FpBnlPjchZ9Dxo
5sEWqh7Y2qor17FeehWoOQOzZXHsed/Xw0v4ZdiZ9/rDJHQdSUMM+ntQgkYwywsk
5hMQvVIkQHzrbCSb8vp7t5KzsUKEIvVOeoIaBrHXslPN8wyCHs+umSlIaGqTj7un
O6/1MhMy7SNjSvpcgVfjKl0mm3xAnT3WECeCTJHrvn9bUqfn3VXUisdjt+PEXefZ
VhAN1mS84ulJJQ6y7IYFSK8FAlS/3fQnsePOh46X4ADoDLEDhnDI6bXKQC+2Y8TU
Pb6+jLC0APH67DeekvmM8ZkPadbm7uJa93MsBf6vZTQ4ckLNbzMxW05WQRhHzUMb
/bymVy9YKE/JPETuOWas0+1AANmSyHMItva8swKz8djbLPhWiuA9XbcgRv5r23H2
JABWb84ebsuVFOmYlivhROnFIuH5bLBNwiHfohAebSqS6wavAjYpIODMrRW703xI
md7yhRKHE800IfFZgJMkvnGpeQtCESpYIacsOzi/E587fDN7zB/Jb1gClkvM5aM3
bbOFnMFOA5Ht2FNkHeZkuDuT10kWU9lTXPPZSbXMv8mxag1oxzhc/s8kuhHvIS9q
Qi0EcPRvMgJJclja15/Z/El8tevUo5xDoGJGos9lP5M8L7KPYr7EHiHTNN1nB5zd
qwy5b3tTzMy6wD3LrEfMf1J8nFkx9bSfii8Uumk1XdVRTRcjW0kqtlDbinKibk6m
MTz+6v65yAiu9njpmgp9+fgyrtlQsxEpLJuLgkYoO3635a5X9p/ujxCQ5hxT6WWb
kOyX8w8e+OAyIQcvTI/5FDcSQRKAoN4M+LwKbGWPxWx86gRwACdZQdizKggXNzjG
iprKnAHUO2iDdk4+i482gLiHHVp4EoxqEZ9wioHGxwb00erUCauUJcEqjmI6r/An
hzQKXbScy2QBIZ6P+jsWzD2eY6hJUjcO1KgIF+Wr3H+XL9JP38j7d1Du9HbMCRv2
rcEsgCXQ1qmB9qRK8qPIxqlIR3dYTMoo98S2wsJpyBwMX4cYqxoRM5Vv3OW3pl0i
ljAYvuciPyORgpWLQm74SmtXEnXjvZmB4XB6qhIfuZrUo4YyptBlqRvF73f9VMav
gEdEGAg0VMt6mCoH4M86Xt7ZkW0HOV324k52sGiEDHbjayQiZ8wg7e8vpRTt73j5
dGUEkY7pDRaAjqAuIKVH0eY2Le1hxQ+yolx1V5PPn5mTkH011fUOZF6HLYB1WGlL
9dVB7ChEeeJ/TVV5CVC+hpdAzfqF37bU7lqNI+syonMt4mqYekxMMgfuKuP6Nvyx
TkpmmXK9JVZtJ7ZVHaetbjn6TCTcCqXOpGthGRl9HI1F9Nb8d43+gI8IK3+FWF65
ht4/CbYu6VaKpXrCWyf/Q29snZT0K7XUwEggT2vYxYuhrY5gJmYMY2arU9cfiP1i
fL3GKc4VzJ1WkvPnrC0khNO8nyXljJxBzCsJQgK62ROPlaDy1Q971/1QADbGz9Km
6Y12E30/0iAomN8q60VUYkFaJE+F5k8hgouEXNmzPTzaruyBVCAMK0LStt/aQAOL
vuoadvrRjnth+JZ/RzWss2Jk4hQLRrPt2dOoS8CrbKlevWwujTM3n0xS5tRvHLbS
ptGzIyjFtin7SxsgOnNRp8XnEKUhNWUzT9hBm0dfub0EZyzPnLJwF0oPCjD+QF1Q
0xMp7ydKr0tDui870dnbv1XJBEc+z7fjO917bXL9BzSCP+v7sqWQ/+2LMnEHJdk2
tjOFJVpbCxTHd65yr5Hfeoo+2/iLe+WgVPPRmIvxcr1YuaAw1d76UG/KXq7869Dw
oQn0gO4KLTOrL2zOZD0X5xyA13NwsXSZS1S+y0BMXmzEA6A+NFBhiMT197o+W9th
oEyCdJPetgiPm6yQ7h8tjMoDqbz8eNCyjkWiTX3KOq5ysHGN2Zs/bUc0EdCtEV9k
sAc0LRNyPnMbloxEm1wHbPPAsPCvM69NlIUCSenNTaCqUeSQsX09GWor1d8RVa2H
jXBF79cz40kkqsSqxat2RGNrEUBBYlys7wltsWzp3vc+IL3cYBg5j2WkBMnXQhea
GcQ1Xg6C4sm80Ha0ixfUNN5VHkFkMXxntW8caBLYWJ9zc0WxuEz5LCR1lIZjYPxa
GetwGc6zNSm75VNhRe+g23HJIL2mNQxghhdrydYp3TLhk/LrbqRKGIAgyh49onLu
SL68VG8DPJoA6aXYNb6tVKRhDJUCAMuUj2wbZnwsggoPXksTK7mthkRNX2/3txiA
rAo71zm+izIjfJXd7xw+I7LdntHc9G7x1D/bLK8mz8lDnquwto8s7Xk5lYVAZg+0
0gKXm08KakBG+Mu+UjA5vhNnUGe/+a80Y2ez5XLT+dc6IQXQa2+PH8MZf3844TTZ
/FCnO8wf0XFqgvU0Vp2Jqb0GjycvNSnuZg90uQTgsm/mPc/0baDrvsYMvZCvQZ5v
10ciOnbN8D0yvRCqSR4Fssvw+ms6PiAk4/ObBcTLJPYkdvAGAX8SJKJE32rKYNQd
7mfSvbHiOnoPmhMAMMSoKJY6DzxHs2HBxtR7K9w1C1dl/ihkmonUd1k0DhwMt4vV
mGxljAIF/WFx5yf4ag3AF7TDLzgOlMJfrsXxYZvPI4GPDHfu39AKIZ5Dxn6xkdKF
PQzHjNFYu+gfYcQ3zbGRnItr8BIuSsu8gSVvXtpLcnPO8CqQjvwh2x2WDop/QpoX
dyjH/pwK9bKvdNE+2sCO2VrVEmv1fGYdhCejzsfsXu3iOZojIMvAI/jssWpk8d40
nig/rbIQM8EYuC1uq5OfIDOLKUHqUhYVsH/6RrtFLEm2w+llkeUlYaW3nXW6AfJs
i/u+1qnoNHwAhCCNIwE75W8jkmSvWqPiiMWPE3lQLMKDk4rHnYUbBfiTQhcwgXRr
u40NhXi6BXHbuaVwux0sLPi6qWEpL7WkO2ZfAHMz+KPH4T5nIOFGZStM0Q5WNFcb
aiNsZtT4qGfW6r3B3anbNerejrYg8FtHYujspWUErye2Lgln5X29pmnaXyrkDz/Y
y6MESiUnnUldJnhHk9CzeOICqPaFFO5aWwU7W42UZ16etugkB7e/8O9AsfEcHWlS
9GM4JVhAvRcKcPj7M4DLsg/J2aMarNP4iMU25z0Vpci+fHu0L+jIT9bR/2atW5eu
I4KFmlZou5iR5YluGSEVjkm4HpQ4tyVmB6Yi/caEyDqlfQJ+yDcYIL446Nlnvc8l
9epQRXdck9GQprZFT8DZG93yqBinY6VZUmuyO6vXTfm7NV2lqv5ErGAjlRJF2Pdm
EbMgi075MPuBBTm7LvT/yi0u1Q5WALdOnpU5QI9pk8xjkgn3D8uXjYCsiTwtma2t
PI7tT7H2fDaX+PAw9bhHghVCfeBu37japR+M0jAuEmBfFsrTYDakaZyfzUUto0ko
kgGA3U3FS1qK+MCBUj7oTqytREcRe6+xmWzjkr296z6E/H+IdgFh/Fw/4J74iwGk
HiOLVfIvOsNXMG5Jv4bNnt+o+7yWVicmTYTmYPEu9cxihjGngOLsAfyMMW1M+umA
EcBmFO40Qa1Jsb3CwRb/od0/tKD7E/BWQS3nLPOR8MpHunbh5QPtLtliUISzbBGY
Tnq3WQ5nRBMVe03f5qAENmdgg2/eEQbMJsWhF9Ol9GeebpIxc7rfSQh1oWGDP4ZO
9JJ6cnYD8+V27+zttxsGnrlFQFwVGVJgA5fQJ3Tm/Xt3bUcuZGX2hCV5LsRU7r3G
i31uDH6aZ32y/jvKI15YDfIEP1A3rdHR61lHw0Gwo0gYHBRIyaA2dPoqvk0I5cJI
iEksSidTpOIoZtQwWbzyID0SoRIZTa8CykA0cKNG88OuJ85vogMohbipqTtrHyyV
Ev/sYN/AiO8ys9Cimps8uHAfXQi3IOwgABfJbrH3nL2f4Q2D5ctuFLDbNhd0Xj8O
zmNpvirrW7mgClcVhqiOdnbaE/rK4q8XZ2bmWArUK9hPVI6Bwexe60uo07wj5Ctn
yD0Xv5KfzH4T5ad85RqTYbdV9qhNP1HUP+f87kznQJa6TSHZqpKrIk50+M5dxvdt
mjFcC4ZUzaM+6kEFB+a8ujj5HjGtL+DPZKg6IKvlIeYFM/oRW8fXH03mxcatjaEk
LvWH4kXoxnc6LCJdA9w5xMsDpkkunhCOXJlXHVFj0Rgk8o9XW9vr+ZLOg7I6LIPq
TDeQYLGTQ/Q774Q7+KOfHw3wS6m9w8g03xH0updpAk9sILnt952NgOsX1gNmGLSQ
Zfy7BZPngUtntM/SPzDfxLWaenGL2vZ9+lDpE1sSrbPKUYW85QAgs3huIgBvjNAd
19cCGEUlctOZGnEkPbTS69LZnubtodcl/MENl1ANd/ZndBcUfDrcfVVgymWN9u3W
PVaI1fkRKvLBeKOZqbk9y7SmlRJVnNlXAJO8M8/fH1Cf5/9ES8G+6mY9ps5CYtZg
czOgvEAe0j1B8l/5+UaX7zZk0TWbMNHggSZ7dA55AAkoBmep0nrJrOK7A3XAGHDJ
0BFvEAYOAf2SdiOFw815T9To+y+FURFLK9Hnmyy/Vt27MrIEFsgQtO8FaE+AstU/
s2bbgaGJ33cqgq4AD68ZXZzJfNuAJutMq7R42lPJKc31Y7GtWOCkktMk7JtIK9ua
qb6Qo5xTGYCKVgZZdsfUvszks5/TufzHN5LUWQxGbYmWmKBLW1HsU5JqhTigHCe8
7FOT5aUmeET32eA4KBPX1jg4+QwLNcY6u501+dTC0NDZszP3gxV7SSLVhr5KKCma
EEzTtMzohpsbramEpXSZOUJnZS/GLTlxDZh0qnOFlP5B0/mRXeWoQ0Tb9iOhJf5d
NUyIMkCQG3ulZm1FwuJyblAdYVXgzzOQC2FNTMxLq5KdfAZ+1MToSurliZmOc41A
Xo2OxFN6qg1/hXnTygJMN0XsPHS2nQ0NRcqXQkxw/+c0gnUMR13XrtOyPFLMN+SS
3gSIoDKMkdnduO79R8bmLWFKqrojW0sY0mfRPcd2f7VFQrLIjW/lkjXqI4SkrlBE
CuXUCDJTbjLOENHEoKsYSEidhmprETOol8ZfclFd/bEmtAfrpEarSMtmE33HFe8Y
A0SIj5rO3AYaDXKBwKLnMDYW3uvaed0U7mOaZJ9YnaIeQ2G92ut37RV4Ec5AQVLC
J6+hOY3VfMeoNxHI8SVA/anlnezbUhfWVPuZzQsZTqf6uGEO0grkyTpPprxYSp+5
Wx5JA3FVpnM96FkI9b1+/fScX2M52CM65eWqzEZYAkasXJlFDYNqsmn7Riex1Ltx
N50sRCWxXORrdZxODtR2AQTz2DLdqEkDoyYKRCbiOKU29NYXsIDsnbolTqtgz04Z
1dFitPzbRM69nGzKMoVrJP2Rfd07lX1TO7ryaMv+2QG8dixhRvdGy9RJjgdjE8HA
z+KwMjSJj/GK1KFirIdECAAsY+zzAwEZYvtptHk/26Xciem14CWSs2ng/ulaqCyq
ypIBZZhcsg+s4/uQqDJfcevZD5/NYE/oJXWX9zrNrmABiDJZmHpn9YS+2UQX2r9g
YaKEbFnPYpbMMO2QPlCXjgy1YVHbY++9YLa4VIJrVJnisEWehc193IiZ1x3DSj6k
auOZJvjZU/TbJJ2gLtJaUBYazg26HDNQFJ817huI5Ik4fLXR6ER1aj4xg15UZP4L
EctCaMsRqpOUdlaExQ1frUroAFp4yax9JWHId43RkwAcQh3p9ZGb77kT0gkLwZpN
J7fHmf1JcrGMh+txYwUV65MG9Uyscg70U3cLX4JR3Xax5xzhLl2mq6Nj/YdusQ+a
99kpqiLvSyp++QIxkUTdAzjTh0DGFSh8hNKXX5BR+yzVQqqqBo+hA5mcaCD1IjSX
vUPGqWDu8RPHuiiK9STlMJGCai5F4Bou1Am7D7jCOoNXUzLLcUkCohaKVKI16fEU
FneBZ/YDX+vJtPkVe/xDX3VyLcXnvGNBuSr8G5Q2ZI0oIc9W+uTCN2rR57LYhX5C
9ceWOPKmm3IztQ0nz/wuSdHmvT3TaPmkCt0gnUN8EkuhoKJFLS4/C1Y4fTIAA45F
JV3qra6FR7LvPWbeBSeaqrcOcZVbAZHy4Typ5qRWLNRSs6aGWC3pVUAGbs7xTTda
EUEEpbNVHPuwOgPaPkckkFquL+7fPWJqYriURxL4CCXIKTtk+kIjIgBGcpiSpMZ/
l0inpAoIJfYRqkl8c9pjzDe89aR9/hTm/6iLt7hZGoXbC1DeUCkdMQrmStoMVQUs
j7RJqjX2mqTWQ2aSvRyIVCE5m+EcOyOJ4eSYeMyz3SSrNkmP6HEIGKAveimn8jqT
TexJA/vnVnb0RNLRAZWjHO8IIX/2PQAGH8xAcqvzB/Hr+jZ7z6c4rfrkfFINdDTq
2z09oBVHg2Ijp/kjBV6WQaYKXwTxT5ILuB9intuZHHTz+MVwcG0S+juU7C4HhDvg
tj45eK4MSN250VSa9t2SAYFN+CISscleRgZ1tOfWRsxmYX3wYdhmZbAxfOyqtIpZ
u66Fapu/hFrxerjAWhbo3toAPk38M2066RxMczI6wl4AxzGVhvwbCeGLNyq10FFb
3Kt/q74Zl46JETP+YpchcC/vSZnLFEG8vP3t2gUKbKO/hRARLBYNgw2/qU45lr/0
aO2y9/WUJZN4fpNUUG5IVQPEnvff8MJLou0Ujd7rmiWiJQ/vmCTTikJ5x8Ba3jni
WHhTd/64PP7O8/KVWaA+SvY8qbcqKvGK4umsiHujzQyJyat6UItLx+LjNZJEctvx
gDVC0PDY2dmILT76f5Z1FXHHwkd4+33S0s8PDvjC3dfMHtdTyWoMEwExp/D5CUYp
GDfJitx3UFOPD480ycM1+Ra0UjbMsjdF0ywfj2jWNnDiWleSTyCJ9IZXP5IsbLTI
IHE1EgBT5U4H1BAVwFGI2wX25ER8fjrcDPaXh2a/gjpU8zu6+WFXlXMix0dUCnfc
irYQtG9Vv4uEsBWb72CASu1/IM+Bkn6+vbSV91hc6xLUcGEWSEcsoKlguxWoBTzV
GsOd+XeFkFepuTITz8P81wZv9XHiEXIEPSKlnJnagIUFcaMAMcaby+TH26IbtjEr
yS0hWa0WgR5YCm55YAxPJaP/l/aI7u9awwyinIk7o/W910G65xb7sVXEZ+5MfvXA
XyWJ41Jy02N0DUvwqXtA5djgrpdw+j7A/T/RGCrEvYND5Y4/RAd7eDo6nzrmLn93
MMo4A3W0IjBDmpE9mW9Bcl/IW/UOcithyTbZxvMnIZUk94pybMHypgJ+O9HdY6Wr
kYUYXrrWuAeQE4CzsyrtCF2qEkQyZPQcgUW2MExHGP83WORMl8Plk+C9xF4i7hn4
XBfymZcuZ42P85IGeC0gBDP7kVL4bQzUcVcG26J5tlD0Yf2ui5VjpcTDnaJVBcb7
q9/V4npRejhk+L59uK0CrXM8r7uZxtOswu+Zitp0mYlkqkfxj/DWqKYvQZ8Db4iB
S7sxenKszAbhy/SdeYBWVV9AAKNGDO5VoGmuX5AsuCpDks8UnDQ6fWHpA4TfUmqK
C9xvE5/iXVU+erz4/nWjIJuwEgvHKXM6B+zr+ywLFc9tj6w+dS4yzh9teoGQzKq9
QHIPooNG0VuexIDqyqNqL/rXrem4shMsCcwAlxSod+JY5RvwaFPq/yrPBQNmX5Bb
P2OvwT+4aYyJrxq6YwGhvH70nFOXjSHgInl9bQBDkMiehLAMnhdPwCFJtoQPWScC
ZAUWapSbUeBgn+GdaQRKxXnYAJ+gXthX2EJxNKvJs+68WaSrRb0z2Q1tc+oRnZ68
SdxRtRvyHbo5uyb/RQDLl3gOjq4iGd2ZH3Xt7lmAkJbd4W2Hm39D8KVtrI7YCP5n
CUcmBZNzwgzJ1wlkwPIqJeshsOXS7ZhTaHJbNxoxvVN9L+BJFWlwPXIibDg7O41T
vfeJW/YaBxf5K+rfjIotSCzl6QQ6dYngP10/BorGMFigbBYKNl6Tj6ylFcpYzngZ
gytsucriLhCSClLGReRRUAy8zcN7e+d/3UyVebEOxGslw52GChfpID9tV9bPQBQR
2mLGNujVmH/QKC+m1Q1u9GZoVd1ly/DILAjRQbeiqEgPsUoda9XfnehyjWUpfech
+01J4PgxvCQOlZKucaUL+qZ3CURVdN3ncU55rf3AIRURQqDD2TQxwHT+nANEcd9a
yhsJorJmamytWung/vFCTEaJWcZZe3Ps8UNkq6p+Y2wXuAd+1xEVepnxtNKz5r4S
DBiu1ylqdXjK9eVC3rWSWSS7aNoeawGXl4oq+or9s1drxzaGRqqBD39ubwA+tCRI
wI5jDrziB8Zq3aEyZXylRb/sxTKIu6RyYW/BgTFG53dgOhiIHzQ2X5L/uhgikC3x
938Ruj/vqGQx/YS9Cp4cSSPMFVT+qyBPEUTakd9QrZUjzbABcTHUf+otNucm7tDu
pUWe0b50HP7uyLlpGwQS4cZmZ22jxEh5xWpTR1AV2++co7tQJASP3PKPLULxIPdZ
v4wYNXLK8PXBEWPIdabDcxXwtKPodlltsrG7G9lqhtPavsdosI9SP+3u6y75Ul+8
WZQElH84540QiS6/ZdadsnxUQzJABkFKrskdHMvged28LUPf7gDsrpPbETLWWs6V
LP5VvOqGhdi8pVx6+l5vWuE5M7ks9KnwFDY8zWGEe04DnShQZAU37XghvSqrhr1C
Hp/TQ/I72z5XGOw83yqyBhwHIBPe2P3Db2M5YIBXISrufGVXXca4E2kIJBxWG9bm
ht0w6qtaOXz7FJF0lokDxonroYu3lb0WVhOF0H4Mlmn2l85nzOm76pnOctQJ9Yvb
M0p5aoZj6nEi67g9DIPIN0+HNy1DIB2+YKAScjGAjrKMfWXQoNYdkpxrUPcUm4xe
fxrMDVgVO6tkc6yqVGtO9qEGTTVNeNhVwCIepfkZtSMx98eB1DOFwOidsVf1kRqi
iExMH0hvWEOTXs9odBwIqvL0/e1Kqti5mkA7dixGnB5qQ/wGfwtSvtV6pgaMtgWo
KRZMmSlITP5d78n5l/WNR6cKi2kZuR9d2VvOcwc3Fm6Gm6QdiZjRq8WNyjIBfeoY
RDFl1AFuLC1XJloahbmmw63PFtgfpW2tmqR7Ai7ELqos/POjym3Ff4n6tx++XOD2
tFfgb9y4KiPT71g+EOxks2A7WVJza5hyGqgSlN7j43VM/elWDcwUpQf+SsZQ3XWd
MqNlWZZ9lqn0EWv9LKL0sTTEcptH62MYq09x4kI1ib5auGf0udWtMoRFdoBeZieG
Mn6wIDSdOpDDw8XUQ3BzZwBUBtvf2jQQugxGI9kElX2kKb9jmb4bfMUt2q0VG5VK
KqETbWhdlCzTnWWCc93ecprNXWfBHrJXQYIc1yCSU5ZZ91t97DHHyW3Ie53w0WKs
BWv1VoNWzqY+QQkfSUP5B3bYL3qTPx9FxDY8cuWcMuhfvp2W7V3/TXByDlp96Ef/
kE0Sfi3IqcCQpmmlqMi911hBoL71zubQc/Kwt8wlZY5N2nNYkkd5G64SIEvH4hmq
8grNC5A0aCiWx6Hh91mFpEUVNs3e2s7X99J4I7BiD79W6ai2X/sGlqFx3mNTKsvU
IR4o91zg8zVhFPR3BPFCSmPfHrbmztswvyWGElLFLX5K2LS0AeNxmxQd3IBXui5m
wGEgX9T1LDR8zAiYJhZpyRpOchrHOzLUkjKM2zRSJmxhztYP2yGosAMmMjXeEnzO
uxL9vMpzZT9NTOgsLPaWGVSWH6j7gF4b30Y8MpdKvE6eODf6snlxAZKWDFh82UC5
OMGF9baTdDOdhPcbf0cHoMzvmM9c9vblOjY3YblPH3J7Vxk++/uq6MfCq5Y1HPd4
UI1Mxplc0RqaPRoBwpOj3K8KhNYJTOkXUwcmSjcu5oGQ6ouUOlXUKDONDrE9EdjU
6kTybGLaZ1PTJYhs1SMd5bXC+7wEYgpL7gZtBMpTmWUCfTdEGdNUTnQ2pym6bDY8
N8J9qTuK0b+/BFgGW8bxvyxdtWLSkTyUc1tsFhkyBl1rl7ryySydbjZvKft0b0ed
/sVfP746CFXx06VDGHLrCHXa89lKCba0pVPaaG+fgOdit3k6cAPd+YL1RV401Ns7
+DiEtieEIiDaUzK82ea+PYDbkztmFWiyg4WgFwtjF9oeBcz5At/EOfppUzZ3zJg8
VkUpmO/d5qUJ43pJqjURc1g/5rV1gwRfw/t86pgtIjXxvSTs0tVitlJwdPYBv59b
NdseSGwMV3O36SwXVbWwXQozLOG/nVFoPkEvEZSX3yORhOtDgE182tOfcXLREkSL
jGD/SzHSTvQmZHojrGiYAt5C/01RpHkx9sZuXpXLCgzVdrQz4lddji+lZ/yZSPVg
FB7m6no/rE9DN1byP7H9NFHZN9kedJdV4O8EvrAfeHF9a/JyOE8XeqRp/MulW9W9
fFv3slFCcdqelDxqKpFF1HcS14ikoPSwOQI6HPeijR0YelPBnVa6fqTgWnORhURa
Kf5s6EPRKNzauwtWZzwrjXaCproIOM12tWDOCJtoM0NkMkiSGLmEHilXWvvJ6LE6
Xo8Shl0zSPpSRNVDq24toihv4PQaB331gDwsydKEUzmdDbu8MFFmXRZtuSJLrWJg
YYttzGZPAuCGJJLyP5a/FZ3l+sx6J+2gpHzpEVm9SUvMru9snHs+rRArYWmKN7gE
OudHwFWQ705sF0oCBE/D91/R0Dtg0K0jRlpg3hJ8ElJhinLrGCSCyi6RorHQioi7
OX+uo392TzToV+hFtWA3uO9X2rNLROmvSv3DV9eOkqsNCuTfI+8av5r1ArVozi4m
6cUCS/J3cD/AanL1MEoCiAphIEGKfZZTUC88Omo7fx8MiZ3yfIsvGWw6vEsB5ikM
PiFWuwXJj/4OxN3RJnXq3eRLNKxdnVRETgvhV/LVjGhGvAcJhBdMNXdTFjJ3cuzA
/ezXKVsWPCSnGk9khd0uvs/Z1RzJV/8A2xtNRneTNFU3eZu4ZcxK4H6qt1ULNZxF
TzLi78PkNRI8c1byQ4F1SNq7sG1J5qBnpb93Can/kCJR59BeELRF3MmJ2fAuI0hc
gaT4SPJG0zc9m3O+vcwxbdb6b3BJXKFEsSZTujvzzMkzErpyi/Eov+eLAw4lCATf
KUPepwkjIwcLLguSc94A8zzEBb1xO697REm/F7T1tfNAO2Q4rfWjMV0S1g8YndPa
es7XayzAPgl+ypX0Gt/MTDsudVJxsm6NHySvueWFEz1XKCn7ZuQHpraPN+hn2Kfd
eHfTjN3FZjJgd0C1mTfIwBwGAbb6e4rzraKV85vchuSY3TchTSoQC9vo2sp9JLfa
GbyoZABmZoYCnfKB410k8iX66KQkW5V2OvpYCr0Tx+SejHkL/gKq4rXx89fHkPwL
5k2IyWhvMWOvSqe2HlhJ5NntcNwVpOfe0910Q6Y0vLqTu/mU3EOjElba1p9XNMkg
FQ7tNPUp8EqDkL17NFPL04lGSUo2PjHrWv2rie7yrRchN4oUZ1phDXxUDPXgsy2f
ND8+qalhoUk3XTo2ILhOO2aJFRnyBe/hKka+1Kb3ip/q7h1GTUKX6wCVYyCdBLWB
MzV4aVj/S4+aqEvJhWhn0kSEf2B3c/uvBJurR6rxAg4v9JJ62liNlseZDE5owjNY
M7GVgJBLW///UTWp0Xt4PlOZ0sTbjA3g4eZds+aq51RJ61bhqzJmO/jV2khqy89E
KQn+uvCzXrHhVCJjU4tlNaxuEc1fsuWcfNoLYxoYmxbDityINbVF5fZ/p0XzrAi0
iqlTKvYUgWrsxIL0f3lqrluFWbYeX6erqUoOnr4WIKMxsntl6VZx5ck1BktTOzTT
8gtacud6JhRePWEoXBpzJjl9hV6k8L/NEe/6xtUDRBCr88+yuN1BT+qNpb2s9dAF
7y0mjtijbn83LWBaGW12zdz0Cf44/18BkJCTGDIydUlUUeuwcdLyH1Z1TYJBp4S8
opH2RAN1HHENBpS76fOpkcbEA2WxEI+aTHuvq+XSQlsXqo0RRr0uQQoX0IH0LYIJ
GiCb3PF0UR1FJYLPYD4U3GhZWLqnzLebe+GVnwNTDa8U7/O0Evb7cju3BKKah0hO
jcjpLt63X6S7epWwa6xhDhDq4bK2/sZblRhDmzUjEBVZJdEAK0cT35TGXv2UZtia
FCpSqEd0iz/4gg1seD2HYmw3Pklo9DjqNGs30oRcNIBeybYkWaFMuX0p0BE2bJx2
rpM3sCWLyRKr0zcjadVuundpWPyTK9k8jhp9X0QfyVuJdnQSlnkDPExsvYl3n4+Z
6k55KkRJ7KYGj4XLGDuaNqGD+rGtRQpnSdzQo6Bi7AWNAbhEFY8yizgI9XiUFT65
T8vmmD8g/WjHJ2W8SDsUdbQlksR1SieXThR/U7/7rCR4o3+jKw5ekdAuHYWYQJVD
aU9nCmxNd899KdLiLFDj58Jrrk/duF6FyeKnXNDem5EJItUUeEKviUqEkSiZJbZc
wsLrAEkkfrp7zjj4CiXKUa3FlN1R7RWbA8KwY8BNPjeYJ3/NUeiLe9ixtHcjPsHx
2JpZ5DVf35ErVdu/oDdXUCIt15gdzhK9crqLqSOCV7XYlySiYbHbnPip04kYYYzk
6YGhd5y6znHbV1bJkd0pY72XPHNGBd+asyPNLelOl3BK8RGmSbkOYtrUdtIlo35d
ivtM/sKXPZMpVJ++zFDjuu3613y/OOzQArLXsIBIELeNe2Xk7Vbd0dBzAyJJNNQ5
RTrlRGpNgDraW3F+Apnp45gDWVHt5HUzb0NLpGg+wGF4HYy1McrNTHp0bd0uvaBY
68dYdOiTFi/ta84/heWGBXfb8g0x4dolCb9LcsTdB0bwgE2ZFUHLT71PA+4SBReU
2488+Z30X/+6a/0zXcqViNiN3OXGufCydPEXjvUAzOIfW98Y5T16O7717dhDIa9P
xWN7+B7VFkGoSXGftL0YKy/sjeK41hhnnPIbivDw4rY1PRMEcXIuuK1y6j1e5Y6z
OEp9NaSUaIZUya3jNNtw1oTLuCrtL8lQ1vGGLj0F+GtBjG/CunYcWFlREqTS04Cm
xEP1DQV4kSTwa/mTOWgcZONk0bqMdtqqYicQK+PiYV1EGEL4xmje1rquDCK5hN3E
KD805iHvQaol+QYqu7sNt85BZqJTtkoHCcea9tLMEp5DSqaUKA9JMuDdfI4NF5iQ
g65fhra9wAdW3VJ0fu8c1F5WvPP7ulpR54m8zTwzPHwAO6X/V7TaVcMVNazBl8b/
ylvBeVDCEPA7t6kXmUnF9EPlFcE4fLNqusexOdQ/D8TeM3IaeXLX3+VQoyumMdsS
pbDaI9Nvtw6dbFbR4HnzwkHhWGT5Zp+U4F46RHBcw3fMYKfOCeCHu0V72qe3JucH
LsDDx/oHuN6Lq+hdgC0PPr0jqOctfBrYNRPTrTZuSTjvx55CXz6P/eDWnhkqCdm+
Oo74prr1et4s43mJARCEGSXR3FSLeZrUFM+JooxkydGEccpDj/L1Wb23l/UAq92u
jtGNF11UDDhZt4NdzpcC3d+MZOnHsND1KQbe6wZQ4R0yRO4i/YF/b2Ah3hAVByFM
iZ4W/YIcqdihFh7HlHOtNb3Uql4g5+KjqEywiEjBPoASZvF1fA/Mi1FSDnPWr1/B
pQ91fhRQ+/mC/ALF46X4LHnTZtb1a10p7kRKW1IEduSmgmuB7aDbns4LOIGT8zWm
zgtAxGBJtKTQZ8YJZxxdLpPuQQvs+2fomxOUgCX79bHtIjlzkZ81jHU6jciyYbrY
/xSSeWc7i6QM9cGyJ7uYo2Mw4bkwYzyKg0M9vWJlewkkJ8RafRqlLxPlp/QABo0c
tD7w/3lJKDxLN8Swmym9zDveZU6e2mnUb9bpVnOiViDgB7uX38m/rEfRXLDxPwxc
VOGCZ66rR/hTJ3baLWlfFToMcdDs2eTsnN0CqE38poxC5qu7iBpea2rM4vIJTgwR
hmqXwRP+NzovfZw1As8r4jEXN24SR4TaqZf9aM2dW7Ed9Cs03Cwe9AKrNXW5tU4M
zIE20M8vzHC5KMcxE3MGNkaVcZ5kAZh0CYG46du9k8JVwiooLiRMcTPoE6g7i5Be
gSGeM/nApjOBxLzW1PKCKrD3vwg/Ma7ivNf9W7mPl/14ZQGDGoLRYAhxO54JEywN
T7Y0s6Z13sVT+5Txd+Xb0VlcHuQ9mS4I83YPchuzXtRhhQO6DAKa70eM26h7Btb/
+fdHCJw/shQUGPeLMz2Q9HJRIklIDRtzjq95EAMlJ+0NzB7Xz/K5WjEwzbMG8yfY
QUdgLuOwmOymuTKrFZui70hO4uNibW/wWV9gdNByfrcTuamE7skNx0i8/W+R9csF
FgfA7TAKlLoX3fj87fOYUOIChlZZkyO1ZwmMXQpmz8QwUMd3XFAzVv4eU4sZGLEd
XTRbn5+e2RTMvrou3jUVicogw9cHiMmhgIMuJDTjoWxJKivzkSBFC5ORZW11++Hu
Vg00Ht5KvDnYb97sdQ1QmFIkdz7XAF1jAVVYL5L8FOA8iWHC94BsuVCTiY2UnjFI
IjC2G9uW06EVKwmSCeiOZDgMz048B9B+DaJB0NmbHepQ3hlLZIFwcxzzT2YpcwbK
BLqXn07EtSRuQM087LBASR9eDbe8aw+uoow1ES3I4A0+RZf1MjzS+fQaJn6lGv1l
z+7Qo6euCsqq2I7J2XUfTHdUF/hzyUxIheZHVXlaHErhzWgNOgMpnvILom6M2C9q
A79SeZMEv7ZHCBWO2+C04Khjee1Ng4j20d+Y3h7twiRjpy8R+Jch7ddmrtb9/WB6
zapaY9eiXPy5yXnQjteLSBLS1PtUBEIDFX62gRv18qFTA5tdUQn3/FmZvbPTCdR4
Z8oz/xTHp5R3hOkoSso4put3zr9cHio6qSmexrAaeRnTue+JOQmRIsQXS+AQ/vlt
Ysh6N0gYd5VVCUIbsfikMx7N/kp7GCGpshi9eThEVlaIHyBOwS+7WD42Fpypgc+d
Uq0dYufuGniwQrBEEWLISJsPEpefGJrunFM7ZRi2NyysvGo1WtDsKmRax/q222kC
SsQEtQjhM9aKRBj77g8SsgMQf42ezcBgttWOJAdzBptcBHXh/J8L4Ys8CSuQvscG
SdYaXiZcStXVaatVrcGhkpEusJaltMqeTilKR1Xy5KqCH+osDxYwxmSIA7dde26h
NNOcIlDHAY92CxNe1SYR5XWfpw/ArvR7BdlPuv0DaiYgYUvnhvE1K8PIsAxZN/IA
OWPueKNYuILpFa6QOFpzfaR9ycdsA/bPm8NjSDA15GLYvbAOBKt/ofQ+C25vFDSa
pGmWwOd13i+wMVT0hIrUzkfVc0Yt6thhDXPsHoKhiLeSEaqV5xu330AL9y9U9icD
izdGFCL7oG7NEywP2/iO6jhtvFSC2zSLcLWyTAGI/E+hjz5sBUzJle3++A9UB+W+
DxEpD7BJZp+hP0S5ccGpFVZp4a29os0GSBKkxUJkpAh+QccNlLAJpkE016BeyiQT
0kPH7zs6tvGM57VBAlTx3NHiNPALNBaLOk0c3s0sLGbyhTfdLA3FwP28vdDM5h32
lOUvXLUdQFpDozw56oee37KlAWlpk6R86HV1SV9ZHZDmGJpP4AlFYLepRWMlKswb
TngR24WBv+BmXoOcuUUxsnf8M2IgKp2udcYltqtytm3uwXQUsgBsqP6IoK4rsl2Y
e3ppfYZSQifC8hz7dbQf5URurpPv83VJYvJN+kB3Wl9PBF+GIlkD3UGHraC75zDP
xmZ2SpPBAmiyTm0NXQHH95uTWDpR6L9MxphWsT+YaEWwVdrJeUP0lWwZEI78ZRh8
PB3Nl6TrEu8kUZByEEFHa1JRDGvwemc0seZQDXMnADfDOdtwQ8lWUecjz+vAi48a
xu9Cj3PsP37lKaQL/G8qC3T8mfUb+E2+nL+T6zX229r5KEM+BuoqNoJY4k28f2bG
1vQ7ABqducdCrEf5Ehc/wq+k1OEf3KzG0a4LNp7IAbyXbLYzjqM1Ysf9E2aWnFpf
V2LN8S/jl+0HGqJmAKFX2SP0NHpnT84cVYvjd4lFi+mYRuMOk8ayiZD8ED6d9s5g
nH2quzgVKN//V6XEpRG1M+kLcUIkEdVbM59n0TMfNjC0g/NcN1HqJP7Uw1sDEO5f
ju/Kx89/qN8Fy46EGTAef1im9lKJAZcXqarqZr530DyhM0GifIlIry44ioi7ARpi
BCtda0iR/PSaZ+JyxnNNCJNU11rgq/TjmJh33eAHV4e07a17xoSXSHL7hND+E2Bc
MNqojwZKACA45hDVVoI3YQIFEoiZHnJmVyqxZMyFLt5bbXoyM4dbHLUl2phhYeO6
TP8yw2KxeFDmqxiryJ/UFtvCiWFo4q/eGOSVH9z5HpV4kyh4VDWCu0mfHaSM/cSn
aDONW0xKVF8hvRl+yQ8ApRrXYdZFOr8jUv150Lqr79Lmjk6ikAstdebukNTrPb5c
evc/+VEaWdc89B5dFkxiXxqiREMnBDM6V09v6IMw8RRLEJd9VgM41ID0iKEPg1D4
PdLmq7s1/EgBWvuvgkNwJ6ZLIc0TDvHJ397zhwEGRbXeoxr+Ub16REQnpLfaGEyq
iRLF4ByUgKJcMCkeEKgjZr5nJ4n9Mr97wlgIxOGbigoDsOTDQtIJ1YuEbgSBifns
7JTqJdcnZZoEGqc/uNWKp/oFm1EyDPaJ1yGw79K1emFu+nBZpyaJ4txu3twunDi/
Z9JKV+ITU1lhwnGVPvR1sRTSk3pfu7aPJMU9by9mYF19VAaaOAaZxLVkvhp9VRLK
mQSzdU3wmW1SR/kRC8ATZnXzPby7Ao4MqEqt01FLAVVUJNTgHQaZT7wvdtVJwYjY
M+BmEc+RL5gyNylHcPiFM4uxxg4Y1dKA9oQ1hrfErIonIlIQRTE3em+Jk1ey8Cg0
0tGFB06fEtzyTJRvwhjiORByZEebMAGoS5cemilosgouKNHmVmPe6vRSbJ4TUyAq
sL5kz1AX1ZL8nXvL/KDUoQuwQDX5aqUzw+++RqM1ZajT4Zfe6FtYDB7Za/9KbDcx
RYWk9hqV7E+bLG2EwAzQvWlsyI8RqPDGwB3FTgXqrlqYA00BsYH6Pr+vz8yfvxlN
2JJm/VKOJLZkyuEzPAxiHg+luUx1y3mRABRB8g6buvgoGMNkZSc7hSx+EWdyg8NO
e/V76gYqvKHNn93vcPLUtGlzGKZXJOcukm2NmDSVgNiXn9SkHBNML9STTC2Na0ll
Hvs7TSrwWa5JfXyrgp0F9tahM11PfURHhf5DBGeDik6tdNx2VyCLelSesLDFSGV7
Y2zaL9vsHyeLo/hJr9X70ibdeXT6NUvRFiNS0JuLumbjZxIqZCjMvMSQ515j1QUH
fkPqgSa5t7KSPauXyLlJ8zPFPVMVJUSjVlAN8b0TZ0twYSjxrfM8upBMFV/BjibY
yYLzMA14wjC6Sau5zosENTw8sFfAZ1l93Ka1V8if2pPgvUDGX51fFS1RPrPCq+If
SPbv4vIpNGv4F9QHwEnVi0G/PG+MeClgB09apfKXnoIGvJeCrba363F5o3SNdvhl
qcRiwNA5KG2fStboJeoF79V0oMG2x8JQJ3y8jQbOZBtIl5LgeZUSHP1UGZ8ly2i4
98rtWoasxOnc4FRQ6cI2i4TNAEVqD10xkg4xslM42yS3VfycKs9Ygzs8yxZnsk0Y
pk+CJWc02/9pfqvlJMn2SLPk08xzat23/RrsFPv/GhYsQvDm5okHuqHAsbDrRyRZ
GEPkAkKi8vDvcFhoBybOfqeYTi/BXWrzj7VVNxVerFUD69SRDk/OMY8adcu7BDnB
CzKVNivavDgWKiOxgi76+MSJ67EjLoFYuKsEzL9aAuFtOSLalI7Qi65cRnW5mQs+
4ybnQZi2yusRzy16fzQZv3bHh97m3RfEVNmK6e3eKwO70pPGMVULCxinAWY9UVNe
VfEzzRscSLHT6Gs7r0+DKmC/gkUiTbhz0B6ytmNt5VWCvt9o2v0yza5ldELlOPbE
3gRTjroez8+SDG0H/6x10VDH47oTb5bIdbNddX282hEFpY0Sjnb5xzD8E2BVfLho
oq3emkO1oC0Ga3PWkC8zbs1Ad5FfknhBzquaNWq0WzS0AGp7GlHID00BxOSUUsBr
Tp0yxne2D8dM9EiNSucI0fFyHJ5GLj03Ycn/tlqYH0pPDKDM+ynylvbzXWRxFOUj
84ViBshuJDWk7VJ6zlz4ZhR7VwrzcvqidyMbPG+y90PWwJ3B4jatiWpuy31kZhLU
OxcFf2qHpm0WqDv57xOwLf8MN0akosRwu50/E+i+qW+6I6qTaCEjUZWVdKUMOPFe
n6gCnWsPqnHEWccbczB6Fy8SjQcpFTzmLJ0rZ/utCmZRyNF0KK6OgWDA1SV8S+t2
ReNjlwIOXid8yYyoUPfxXz+PLYfBMUzBSk1ovkxpsPAzxcUZiZwmEqrTdf5GuTH9
vOeVuEnun6S+cgx2CHbjHl0uYlUC8J31jJ60zGkL1nGZWGKh2ruqbQ2A1WoWQtdk
lE7L2eFni13A8Kac201a1J0qI05vhFydp9rmG7voNTsWoj8502srR6+uaK9ytR49
iJrG8SecvrtyhK63swaH6FG52+qYusLwVgP1UXF0nkwOaMSgDB1V+e8zKVTdoiFg
pHllmm6Pi4u/g6z5/agAiyt6yIYaU7A7jsKttow2Ja7IOMxAuLJLCDcxFzJqwfO/
AuLB6BAp9VcNITh04UFJBSax760yF3qwP0acBBsJV9t8NDdV5dQoT+FouSGgz+rc
GKFBjRDzFonWY1Z7r7RH2LIpVYn4UGYGYNd/fDrE0hY+FHvgyzj8+BZWipF5qT+I
lccxaZgIinv4oGsSZ+N5B5QSVBCKazVbMoccILdwXxXCsgYWQEMf40fQsoGwn4K7
M3RBya0l5KpwF0pYZWS8IUuuT8hDznV2U52NhAkgdvBnfXCt8J61BFFlcBUKbp2r
HEBmTmo+qq4V17E9/Wp1P/PeN4SMnkY+7QSNrwpnKPv/W3lJLA5Kf+tfH0sJ13SK
BGYf7m8inohTo8csDxlcl1WOElnO3oigM8kn68odZIZr6d7qa3dsGOha4oGPjGF1
ToiflLT3eUk8ZTSd+A/OQZsBqQOyK2BEZ17Z2vW3AWuOUpTZGAwvH5f1bxvR3PNJ
btQ5g3HLWG1q/kFTGaQn3qvz4UROEfKmq7cfffojrfiBkdQKP2yqYIylh/gMd8uj
1YcTq1xqNBqWVOTWwcH9fT4YoUMzOFuW/bdZ6Z+WUmIjP1fTBWDAAkoS/EOknU00
Y8MfIItqOtGcf0MfhbY8IxBJ3H3k48SDcHYGhUPZYGvTD4kLwWZE/2HAIzRTXclJ
aY9sqftyCnT2zY1VFA9gM8yXOMVi/5ryHDSggERtY1fejMIAyAFmIXxjarbzg3Ty
vONjtlG+Ffikv7b5JqfEaWSaShxQr76ZKVxDR9ZPYH/o7pGLFrAyOFjzTU6Ugh8g
1OsfcS06v4+5RzqPODVkUKW4krLiT0un1lZp0CF+scCQKvJTLJFcSIt5PNeA1Cob
M5O7GsvNFo9A3JOjzQ+tdIlz5OfzrWX7drNJmZeEvFYcJCCOWsW3jXUZ8JpM/jMr
6ZTk9MrCi2I+0nyEbxjeOS2ZMACpwnQX5JzklUIOyyURnNiNcF575pO6YHAh5sGE
y2JKPid2vziGT84+INUCO1uJZ+hKIVhr0dI2pWO/IWKDhjj7n8xJALbEGr2gXJhw
CWyhogI2x6pPQtGTZL4+lowWFT+UTr0lLON77QF4fYUefbUiy9slsMr47juEl5Um
MC7Oq0U6ePnJaU4naYN8fpW/Gcn17kHrBJYnnAf11Mf1fFCaeXjq/oSMuoO5mNZn
TsurX5T1wKQc81XsT7i/LbYchFE3pAZa64PED6oKHSd3WT/CdNfKE4uIW9P4MjDi
5jMyZleFIwgL4SJbF67QV0pu061f5ZqfBSYEv8/H3l1qNlXQEN/RUp7xTCMPGAqv
w2jD9Taaw/EDREr9B4DBf1RmntF5myIcLXrbXN2Oiy2yq8F7DIx6M3TjHkGzj9BF
6mMs+bf1VdXhH2KiW+sT0Zhk/UjpP+ub+blmVRhjgcavewoDVIUurAoI7Z+F2JcO
4uNmy92PtcxwbLffaQW40u7qTtQ5j3uNIO5H7fxhijAt+RvpbA5w3OZ//Eknqs+k
IZYvycTgrt0M+tgwwRkg9mFQ/wuNxX9Bwkd3ccnsxPNbV+LCkoTa1ZKHvTwNXRZ6
+dHICPTLTsIWCQWWq4NI4nT70daumIzMnw7Q/S+pYkC+N3qr42KOdSzqNKzvwZwI
AroO2QAPNHaWwf97AA1FasSqz/ZNCvz1bN2qgDQAFIFf2IvMxZSnpB7AbOQCIwqb
q2fjosUyBOQkTos4GbHS6IeyqrurX9m14df/saQl9DSS4LZNpnhZacj+/uALusDz
E52mCGDJYMjd9koS2GTqSLK7tZ4lVrihFirXUhv0Gk8uH8749WIAfLK7OorBoAuI
UJ5yO+OOFoLekt8D47Mxsxy4P5CidGZKkaQNdOhJU0JWiTG1isx3zMFa9BuSVODW
LpvxQLBIVp1wZw9ZXvW38tym4ILKAaIkfIZydaEBOltLdeNgfVbBdaku65vhrTGe
YiYX8Y03Pu1tX/GMF5fKVgBv2i21NCyVZU6T/tPvCUZ8dTFLc8KtCXd5CWrO6EM0
yZvK1A2qht2W7JDyj21I/jDoAexvnbd84gfC45TZ/WutyxbKqPFQKI4yQWg6XT4H
xjGyRkc8QOGpUAEA3XjXQIWzFYVrRz04XyIwXKwnNi0wB5KsWnRjiptbliQfibDP
YclW2NEBFaGSZPoWZyDZFestoHeYfraZL4V8E7P/jVw0Si/lFz1GnBPvitkAYL1E
He2HXzLgR0xUzEhJuZ16GodlXFiWL0pzHSIVc7HEqECRS/uv/PrxkqbcLqEfZDfV
vrrAwcz9m5qhREggL+ifePhEvVH5X4tljbiadsLf7m5adyjr79TxH5vtvojVHmMT
yHWQi8VFT5LGAG42Om7AzMZwbclv8tTJy1A5ZLf7kBz2qUhqMIvgxyEzQ2BMYQYv
NnA/PDVw1l9rO+MIwYT/Y1AZPWdwCoo0ARzIHxZ9mieR259UbkGTukoAtzdeGyds
NhKWCNuEqfoA0EYApw4ytZISUFi7LC8uHJ1FhRNcQlNbXFvqIqiKcuIynKZWzbzy
Yf/1PFkgNORF1ICa7jnTHSY4pw9Mv0+xIvn6NcAdzpyttB3tg/bPaBptawvXAQr7
ROdqZwkP4aixXNFdWHdon+38BxsKZopjJfx1PgtuVzFU010t2m1PrWPIoJQmGshi
GPA0mo79kY1ouOQONLjRGeFlpob+anBFoa4xro+KOId3PRwHdhuxDMW4eFO2Mb0W
qUTX9EUS9KrLrYUbG0PFDKR0h8Q3QvcRK5/o/AtNd+drKfppBa65g3fUcLe2jXYM
Ce7WyjfJXWiPblqiTpQpo9R+5WFgUMzytx9Kplbr1yZMvjHE/zGflmSjxKDVGNmC
+q3UuaCss1WA6Pua5aY7/LDBJh0dB3hv7km1HIlFJo82F2nT6K9IyBqEJVLnTIsY
9KphRdINMnnbWiUvU9VJgOs1y1f3QRvjCtxyubJIQ49G4mEy460qBMFH9+xojpgB
cxchQEca0vX0VmKAhYDvJqqnIWKuGncOTy6WbJ8ZUjWojnJZKkCfg1+3GDqRP4Tw
bRZLYohoTVfAaTRyHLtagfxfiQmRwOaAr+WLSHYZHhUw59WZHr3IU31imbk8IScf
nbQ/hfN63PIEb9vZdjDv4GUn1g/SmMbyXxaGLPwQQTNAOmIpYbCGkDva/9dnSJC+
4tWYWqG+VMl5JHRKnIde0Q8OV/SrHIFsIoDxn6YZ+5mTQdVRuWtQ0drnvHlXE4pg
nqfm/AULDzmroWqb/tG4G1SInWgjMhID/JZB9Ft9ttGrrVEKucU4fywoiMEQE5eU
UadzruABPTWpdLp+YIJb9iTmcHwMh/SBrv31EpeoRTw+HH8bjkDVtVxWBeXYjymK
VjZGjBr0wK0sONoZiO+sHJ1mOOFGxP4yOqqKYD8IAPmqkMnyNciY3xIrjlsfNzjt
2sft5SPX9IzRNSj8Hd/ox+9orj/0APY985Jb+mkZaIiQP1M6eAfzt5LvyM+RjnhO
YtbaiYPOPpuWCtk/jfzgPcoWDZfQJFzppp7gumcJ3aOSt/uo84t6UZLLaU0bx4Ww
vAXvY5ilW4PEvw2/eDGqNzedYIy1XTUUpdcty9z4iippWnv8VwGcmsQPB/LGCaZc
rlG/BmGPE7EIKfU/38rmqIcrZbyc7jWbexTOt4LNlkwJNB+YmM4xVT9AIPofY193
8EpD2Exmt2nn2+q2u/PK1zQOTPE06QgYj+zt9o8h4lcBtVTl6S4u85LU5djGkhkE
/JPy63Ofl5T35CYW3NailULEh7yXzb0fDzbwoM+SRzLqTSm/9Oj0q01JlevnlF0y
0Yg1UMlC+AZhFFnQXqFhK6lAX0n5TqZa8AZnuX+8aXoumRUI7lPfXCdE9qTMnIwa
/qRTc+2uzsGNlS8575aeIfnGxUX0fk2SmfNrq/+syrOUG3bhHs82PV+CVRJ0eA/h
R4Ok5bGtrNzqzJHwferQJ72SWp/xc04GDRPAgapo18mi0SJQQgE3bARou6XpBXkx
337HCm7Gr1947a/U5rlxUSEgQ1WU56brdLj/wANMZzn2fNg/fzIUqbISeoxEhVjP
V5owSR4QAVz+x7XH+l3HyDkUn0JDHNGLtfs0gJG4OLKMpBu2NksNZTe20s6wUAjQ
tix6MZPcp/ZozmpkkxNhd8ldPs20OV99dwB/xVsFwC08KZrPs3100Cb9CQghw1Lc
+DwpCAH/kaXt3GtlMr6XaV2TyorVlr8BnDxnbACPDnlWME+BKxpMHlgBCyDIsx2H
iS3Cbp9TgkWHekSb+MFadVUW1ER5NNTBMAZEE8PvpBKHM3GWw8px6sS+P+H8lMIT
H12vOjl9pktT/AAJ8m2g7dqy8qHp1WfJ3u39U3Lm+tHiysPj8Ul9K2AXJTE0G/PO
ph+rDA5iBqoR17G/Wim31ppqvrBidJfBPV6pDgjlNjXva/29Ga0Mp8hQJRHS/5TC
yauAGgWzfETKw3fN8DRORWfPuib/wm01LjaEOR3zYy+FcUopFOI9ANleBlsHyoUN
9aMwlwGtjKcCLYyHV/n70fJGDsgSEvnQohg1H18jdN670Cc+hYLBgg7rpxXzCquA
wg1cB2jfhfPmLpyYra548Sj7X0g0+EM8k6EyOWgMb4rUKtXyjZjXgLzyQZ+nUvoF
SBHPvPNZ/u6mxWJiZzCcCNiFJd3UQjcgMIbiWsJ5hxlWr6BztNsSUXlJDtqUm56s
DK+ghQIc7QrzO02yYXfrIIzmxUAYDwlYyci7OHaModmeVyGaxvv/F4RSe4eqSpjp
DI9z5Nt37wbVy/dYo3oYOR9rpSK3MS6exOlL5DyJcRcAopMXfwf0jJtz2FTwdqUH
W0QDLFvUA2TS5bP6LdfNiwstL3RQ6nZdPT1QRbckSP6Zo1iwzhv4hFXHaTIC+BSK
U67gzsI2qJ0dHZLUyl2hyDH4mhCnEzw9xbpPuUz50t4jSxUQzLQh/Mc8eKy9UzIw
q5Kpmisn05orynmFTsODVka0kq3kPYj5YPTUbHSRGjK1fjOEe90z82KM5mmV3Zh2
S6FwxO6Og4JQuTGc4vFC5tTQTEmPBSVzLr8Ce62N5HjOdEcNvG3eHee6B7RAEXtB
JDZULh+ddG+5/YrlLNfIveRCvHOjhpt8lYwdHxNYbG8uJYyM+369X7lO9KwiHx45
M129pY9KlyCDjOXoMaNge3roZyiHHPKsfynWdhn6BJ1yWFwloTAAyrVLaRd09E/9
xeDcTqS3gbDBrrpgzJmSoFNtNdOnk87qX8sPa5o0qjRhm08YUPz/Qy0driVC0c/b
2rROiX3bJnbfM1lg3mT8YNcBHocTN15NRgXnQyKPOyrhKURqb78syZ0zIOo17CLy
Iz4M4Kd2mHYQvJmj/MID/6A95IPE+O+lqRAarM9XARGHV+DvX8n0lr0UusoRKHwm
YXL8pxre3q9aeKvOQ2Axnss8PQ0XSp2oy4dZd9kNF+cUQOtGwNiBPQsZwc+z+/ev
sRgLFsfX6o+Fi4XE0OW5ni19WklGgMgw6vfHYjrMGsYGz+lifBWGbh346keCAsxN
djsWjVoRueDS8D+J6Xz7Cw==
`pragma protect end_protected
