// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
inUzQe6iFE5Lts8ECGajvaJBYwEZ0FGY/tVi1XkdlgsSMDlpPrf2dZnGc1Ia4lv/
/0q/XeVUH4R3Sx9lxiTsXmnurGYDhFH62vzpeyfuUV+2CHxbBkzFN/h8px1rMjYo
UZ7c/0j0PMgcx2GjPWYuj6bDFABPD8PmOSMqE6fY/to=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16976)
Phplwu/fAC5iFNFGP/elxcS6QDtiEmxyLqC3wSX/2P4bLvGNk1g35X8QXJgg7Y65
0QFGrcmn2Y31Mcw9LPOxGjufU1QNcvwFKXDGXqhbsKL9Ej0fqjamIpZ0YhOJYJ4L
hAR4umKLcK27fw7pn0/tJGVEctjrdL4btK3eaErS/ZuNmCmUFy/CQHdVquaCypm+
B5tW1rLyD3z8a/mZlEQLZAsGirUm0cs32OW0kE88jfKesm6Z/8L2lSKeGe+fLaUZ
mhP85w9SWXwv8r8f5Ljn8ctM1fPDDPM3omUlcbZHZzlw+1Kvrk8MnNnjqW+ThZq4
spIX5F6psIcYz7w1eepIyVojFuphM4FvHqBOU0aXIo5Kjifqu3y9u2c6Gnc7/FCE
8rM1f02d3bbeMQexltFG4kZaiPhMZKTBA98v6oPGB2FK8ha6nrj58W9F3ebnPbOr
f37xWU6RLyd4PWUNp6qU/4V98M8/JjAFBq32ROCr9clfpWBBPwg8rdfSToOtUgud
V3e1YQ+cEpugwtKBFfGzswpX1S8is9AsUmgzeVamD2sRYpJL6YwID8G+YqHAcmsw
f71+cfJwj47fxqps1jTz0KZcVwRDxeENVKc9E4SFS3NN7/7q3XrX/obw5g8HGxqt
WKqM7mhOM9Ni3ouG1YNKeUPlpD6g1tEAbkX/fdiisTRqOUxLEotrPf2Wp1M1Dxcf
vbEbQkWWLznfGWjagb5gGGZPVvts0IvMjnNhXWNf8sbkNSztCClUKjdqcMglJCsl
a9WsLWtTUx9/wDHIz36QI8s4HFXqwD1g0ZNwUfglDz617CPHB5TWzuaFtCWxeO/7
Lvvw8cCH6MYe4gMlWHys+NqIgesMQZaIWGv/uo4U+yEujYsHkMxPs6jxbcO5Ndxo
SKTznBzmOMKKT/k8j1VdThIlUimHZ0qCbaTmM9+kB95/BU0LgPfw7Vu+i182vIKe
GaX2iWp+1itUK22YF8qgIQ/DIC+guHH+d8zfCOc9LOPOzMg/VILyyMZOhEeiCaqg
U3Qlutj2749W4fAh3D8q/py9S2+TFnLJlYtsubwSu3C+/MYfl0YozFd5xmdLGxM/
k5YhcO0bI6675UTn/cMh22pS9TD/R/CXi337lN70pdSZga3RR7kZSTJJPsgrKlbF
QNBlXYN8SFiU+o2PVoLcklieKo2p07yy5gTMZwOtxyFGyTV6Ho+y7589veNxqkLS
XbJwjuB5pW5UH9hWPYejC2lk7XKVwipJBG/xyqOa95IUd9YqhMWz6R1sNL41HrmV
S/h31Y4roPcrVTwVkFCaAJZNRaJXhR4m0ffKByyTcmxmNvJHFhuMh9CA1Dqadpp7
Mlc+uebw+ngRrkHqGqJmSRUcQxmrgmKRXFOh9oVaeWWEVAusun9z9tKxuXhx7dRh
yBzo7BR0BVHeX8439uEuSH80us8acPiRXTWW7YdUQR/WzYZE7NZdhtakVKrQtNHs
tovm0g89c7zUlcId1toLRZnRWTU8KvFleWmPGSjSQtl6XR6KCpGulZdofuCb766K
yzGWG2sDooxwd8TLPMuS0gm1TVsF+njdFEMPRkmf8t8b84QkN43i2Ptl0+51B3IO
kvLEcbMCDuMWc/cfC0zKLqyyo5+X9kSr/zJyHqh3IquQFtIS4mRHbGg1+eRsAEWe
TBt8X7r5zLDTbfFo9svKLvuyKYQSJUAJg6fAG80TP7UQF3lJH4u8WR+KAFDvX7Wr
DgLYoi0qg5Ziv+5BY/Tj9ZOR8NxP9MAhpe6OlIBnK/igzdX/NC3huHtyTPtihkTC
N6SqQ5f6AUHL6Q93ANoF8x8BjhAFvgUCBLPBaok4BzTiQ0p5siV/gDn7hIqiHOF9
08tfCn7WynaWUjXKys/010CIu8+vXCY07KocJMe67Y6QLXeakFd6rS4TmS2qSyPI
SctkrLLNXUJfNe6HJ3FuJoq/wO2gT9ta0D62zOfFhKIaORXmUfgr+3UWAu8bqUsp
jn85E0IC9W2iCTuBqz2yFs5A1vl25sGMtFuuYYv5LBN1Estzg6ed4qwgDRNgHC0w
3T15Csq7oj+GSTAPV5nUum5+/enf2T0WEnJ2raz9pWFRcL8duZ/8tJey/8DECTgE
hSALQEvhtM0g85hPMyw4sONe/nDTWsHI4Huph7SJ2Utyk9UIo7pKHnv39krmy5EL
pp/xMdg1oHPIW5cBHsdGfia7vAWocLcp1p/Zfu7d/lBiC1OlReC/K7KNUgJP74dW
RTE64S4PpkKdWe32wuu7/MMYvKAUWjLsp/Mp8+l87z4Czv6JGm+sk8WL31jGs1Iw
KxZS7VU52MGwQsGg3YYaY+d881ACg/fyuy2PdmX/Olq7d0lLK8Tt1tNEv7SlkEIK
dMQW0DV/DqfzvUZAbNylRqbrJpIUfq1V9JiBnu1g0RnDVilnexiRqfcfHrSiVhGY
8X2OI6o5mxz2pGcONbt9iAyH0JzGZrefwrU6uwl4lvZy76awoTyTWl575wUp0MNs
2f9Ct3dZUOH5yx6N6rSZUnO7jq8ARZlV8pF8ntyPvECpEpPzWPwVWlm856oq1khm
CZr2Lkz6fbfaaNk3jZ0sXujE0PIsjsO6G8p2zQi83ob20fc72PsVBpc9FLFHEhJn
DWQjiFCZUxfZR8bO3RrmJFmhLyzPEnUhQL8rhQD8sRK9MCPVFUkww1QVZytWUm1Q
opYXvma6OXesGl3Jcw9FdjnjTSeqPCZQBOcei9r1pEADjg8cOYqEVQWzRQc0kd/j
9dic2vSJuMdhQI6WxofN5+AfgOT2JPY0cxcRa7TmW1YTSzFpCCh3Qq5fpTTj5EjF
vAZXdo40wF9ftej0gYdMpcG3znE5cSYRK2iep7wu+Jpg7DW8i3DhZn0RRokyT19E
o+kh+e0AVgsz7OZrGl1spsTP0O+xBRvDzQn/KIdV69PZW2GVSR2QAwLhIeKrC1Xj
r8nKbPD11Xuy6v9iSyCYKKqg6T7gvgsEFeFveS7+sgoNzbJ3Z0W/liy1pcr/KMsY
SNS6g8cpNfg2+VUopZz8yIMhuDVc7J9wrHdJGUzjIR7hbXak2AkN84EMh2pWohlZ
eDYzMtrX6dUU190aJQvM2Gx0FMiAA6CXetlGM0/feOrYhafgUQXpl7rJrhrEAf+Y
r26d3E4rGPHG/Wu5nCcP8yZDKPMPD4D42f7h7dcbkjBn/6WKxLO4IAVucbuCekxO
KnNppdR1jU1Jct7zaKKAS5orQR5wrNEIEEDhcXrY3x+a0a5Dc9y0PToVnJaz+V5z
YsvyJvvkF34Xuv4Q8pKhcIGrO+bb5emj0CEnqf3BeNewX2v4dDN6ZduVckCzzFSV
BZOjf672CvDgK3ImLJGjhD2Socg9nqe7oUMywv3J8I2s8S8v/5D+usFLkB6WbAN/
B8onuVRtHdZCgo8FuXD9HlaCwTQPw2i6i5W5pvb83muhOGBF+vH1oxmZSNiBzbGp
aZ4NfuWtOYyiSFsTGK9X3SFNdlPlZRy5aediAs8AbHHkc2JHgcFZKuhuXxLGkjOr
xaySP4E3qpraS4C6/ZWbiDmxY41gJJTN/i/ZN6uzQ7LhIcwjLVxdHkewTpv/O8qz
ioNo9aTZFgSTNLoIOyoE/a+oq1m4CQSFkp9C/xntb5MXUn0J1MaVQ7hXiy2D55Pm
qfuRDrQgBlfyywKxEvEwFvyY1tMtgwUyRJ5SiXH2oFQMK3hS6E3SoJyHbBx+EdR7
Ty2fw/KNU0gscZpwmN1ocVNNLaQLY4GFfg2mV7C6bZv/anVk39+AJszDWkTBb7wL
/hlGGJROeinZS6rNXJ/5h6YutN17upl5Kw0uO6E/77hm+u1rxmG3pzcSu/T+NcND
ZhBhuTsl6Y0JlPqL5KuqDRKfZ7cxduxyFJxKBoc6gmhPuKlcwK0Lwe6rspKtY3oJ
fWz6fxCILqV9QvSTw1gEiGOow09JoTHbtANYGG7XdS+9rZU6RkymnE2RmWbuGJgE
GfjyRJEqmxOesCBuCoi+kHUQ5ujJ3YJVDfP0MpdHrbeV6Nn8zhPJMS3MxLoXYHQu
SN8KfgY19J+qTBavfrmIKHkxrp/7EodQnLtJpxwrlyPKrcjGRy0jh6blKaI4Z6qJ
ppKhvaUX+7kW21rBPb8xX2YhYrke1N0xSxGEGaXZqB6vRcuTsiUg2JdfJUGCwGl+
jhvmw7bLEjo8nw60gMuTS9mZT92Ter91Bi4258LXjc01ebhfZgZs9rfnJCKjfei6
LuuQCQyiwLHm++6fUwLGN/uqmLWq1wOkfUDPZ/57FavBrZkSp+/kL+yLHBqdMwPb
mfmyAXFEjpYD0gsWSULatHTbORTLcO33mVJDGZ1LQeebNgNplERBQQS0dO4sC0xM
onBXXmtBEtCKlOecfO8FQpO2zbS1Abch61hdCoyDHY7tO4xK+MXbo6JQe2serecL
qNtpGAWbv8B+QmsAGDCAJTi3IhQFp9atKYBdJceoR9XK65LQXUWlr/rNlbqzUsls
FMJQCh8RTKptgiD+tD4fuc4Fovt/hq4NqX8//wE39ki/TUmtn4RY1+HvlPm+I4fa
lr6L68ZkJPF2XB+hIVxSmDko55y//UDbYrNblvTGdN3QbQ/HF3VuejaDzyLKC3WK
WZhTyVJzBN7mtMu/6/95GUjwWi7XeBxwk4QE4kSeXjBVXmTXLm0+V3N/A9qxH1tl
X1TQfk5n+dDPgwPsMGHbjkXUpgVzZpQGv/UBqStPdWOmZwtFzxr9fdfOYQURMVEB
DOXyYlVhy+JEaoFZoKnJzUy1mEhgvHVJ7OB6bsJBqzZ2t0/uzmjoewJvmyHe8F5g
ft+lkHM8QPF1KGULDxKFAfhft//tAfRBKumNYvk8TAWb3rGLfeZUPuTwUraPcxZX
t9OFdJrs3wVVud3fPcSPChQ26RIHugpcEm2xaVo9jxeWEo91Ibiq/FPz0n/MaKzS
L/RIfOWwu5vTaSyqG4ZBgp42dJYVlvjuN971O/mrqfCxLc/VSwmjDyHE2pbT+MJl
xiQaZR45qpbXJjJINad71AJvi1VIivjyvvVxnx05BK+gpWx1QUNPAj99/PE1TyXD
5Lis2C0Jl+8r4f9fRsg1GSZRF44MYm8/B1GLNSCs9ybz6dpcESW/k8ex3bBznOy5
o8p1vSyH5YrtlOxII9OlfzdAdrxlm2YXGsHw/kF/Ba4XK7uhISqiCA5FcQxv94Vn
oMuW5Z3wjWdW2/cMm4+vPxjXS48D80BHW3PU+PiZC6hGJXcbp73RhTv13eL5uhWR
VbegBT91a19j2z4KwZw/hkbZulbyfBEgphkl58STRsauyI+pfu2ugYoFzTVvqCiC
z8lvDzcUtrNxrUgsqe78xgSCwlNwrFVhayqbNBiiMAN0yA4k0yVWCz+UHYqzajJh
ArFySijFcgzc2tFW/r/U5SzaflyOO7E5XWQP2yJqdUqOntnsaEYwINVNxouZK6QP
e2lI/coxIr+hPf8gW8DHrP6Yu66RQBLAI9bJZZwOFlMcr+9NbZwuVcHy4o9h70YQ
8RffTLI/10Ndj5TDjkR5FtTW+3B64QVQfsEHuQRl+cCKTBgkerWPPYsNscWo36u9
D5Innlh+uV2R4oaydUWSyBdrk/0xJakyx0oOGETtygRmIMzMJAegUeda1fH5MKu3
bAq+7LiZNacosaWm6/meS5BrFconrishPWr5NuvtHvgWb0zihMEAhgc9rlu7W1Du
eZVuotivA07jVSjT7Ocxught+/t7oW6qbXzGQytLNnizdIkonlp6JxuMWr0D156R
UXo5uhpuI4ej6mxZ/MXGKo1dhVK/7gGO2j7qX644bHFRdkqbc3lixXsLoUIITOYk
X379N3jQqUUyy4qLuDTYOvY+Dn3VYz7pkG7wtHCAn6HzPklT1YnkUOiEggXGMDkh
W/9TlyTS0K4mYM9cJdnJabNVvksK2E898c3HyjqqlMYN4/NbYo3EFMRMekCfNpqi
PmoC2AgAfzGxPRYrTt2+2A2sJ+1Dxcnu/jUCMPFwPRMYSG5tULvEoiEDgHSL/hDN
mwZiUakiDVdjFzg9D7GYPVij3e9jAneJ/mOxAQDSQM9oDDfAbpRAg3saptCS0TB+
KEjpKdZ6W2CtEAdCoEM0slb2rHn7m21L1IQ+AFL4hRfpOVNEHdgkEKxKxqwOtGQO
JM8WlaSZ2NHMeCCYOQYV+ENt/APdZaon5orpDpICqoSUzMISsXwK1qaGYfVJE5zw
gbqsxYeg0ycwieqOmH11sQZAWLX+CmMNY4lxxOlqohY/cTsiJGf6lRfqiV/CY11B
ljNbOMtpCmkotAs000qOkC7k1ZIP5L2jf+tq4wJR/XrLatqfxXTaosOq/Leggumg
BWaTFOMoKPdPoI2amYbhvKPpNwpBAFM1/NR+LUdVkk0o29Uc+y5GXZAhW8RuC35u
M5e3vdHg7cjz7O9aaOyHe6hGYNWbnWW3VWBR6sXq/PV1Lhf9sDDsiJO6ubh0PnIT
hT6m2ajQnyU7qSbPhXLXSfh9pSzMm85+9+FCjW/SrF8A9CEgFquofAd/eMSFkaqm
0ODZ2UshzS/oDvT611e2QCoaZ2anFCsMSBEEjhIlQaN+fTFdEl74FcW/xWQg/T5J
zzzDQuoNBgb7h25m7EcsKsRiK4P7qSXXUzKsabvVhy87F7uFoH0aznELx4lfV7ev
2OxXttKZ7U/r8WzXAgzjkK9+D6ayLyM6iV00pz3WksWMAfiBBPTQOLnxfPJUNy2M
py8jbI3Y/S9cFBG/W6xrIJkzDhUSnTl8GZ6EORAcLDJaws0Rr+93Mxk1G/IzA3wD
LeHxymds4O+HoHY+UpuIL2L8TmsHU/lozTMTjsaLRcDvYCCah96OZ9Ree61PwAM5
62SCLT9CatWb/YCQCKrMRBq73xi5I2IhqfhLuHQaWGyC57GyODZnWHBpsuQTV6uW
fM4LFTtkrzThTspYe8wMHQozjUufhGneD97Zd/UI/vOZNVk65BQSn+hqnMT1YNMg
b/g/54XmNA+fRHvH6VDWS6gjTr3WDUJAZTiNrY/hP013jUE0lVVC7iZ/HcotNvAK
Dw5jH+39J4lbUlypBiBB+H2OYOXx4st0E81VqrjbN8rQRd006jFK5+M7BhtLhr5L
W7S4lc/lEhmPiU45sXyBTQ9KXIr6N62a+4Hyfb1/xADgdLekp1jThbgzxggk/TVZ
GZnklFapmosiiF0pi0o2cUWSdpf8DaLuYBN+M65Bu463goBrYU5gJkE2ymqY8KI/
cLdtLLZX+TNovDNzYtcy0k8op27JHYS94/Kgz7VmUsJWQV40GPI2ym6iKNu/2iwK
FLjaXXSnWGGPBjMaiyD2bDIBDUS45XWPWnjBwyZ6yA/wr2J84UW9ppnfvYvqpivV
ptDDBRF4n37idjtR997al7OOMN7sNXy6V1sNmIxkEXipSSWMBfQK5kpOJ9en+Ypi
3ihrDTVxpbwcud5ywUwnk8N38/QtXYW3zHwOHhrJWr327V5vUGx6tVNkLlQFiwjr
iXlEsnfumDXw6QNEFhOtoNWYsf0GdilVNM4iZaTctjK3W6+KfTCURBMU2Ku54ICM
jigFWZbkGpJl69bCtHuCaLW9ER00VSrvSrslA/heATfNX2NSlb3cNz8EZtBmiLFW
SsZNSUUrts9iapGgsb97u/EaCIjZFQpsQ1yKTmpI4n66tu6iZjLlGyxpLx0V9OYE
lESx/BJDWR1hGWs1ZfmQS10UTt5KMQ0ixjpOspxye81y78hweMvVTyth5Gk2+Eah
ANHd78i3xOSp4tvtx7NTRtUIYWuQaQ5fB5uHVTLAGPxtV9oKgNRvyAwEh8VmEtpu
eInbOXEzQjlDZ7kTmglLPYYSHR9/YvYMJsvZ1RHnWL2gSO6ZDIka+sEWbQP7XT9s
ZdNftdI1afvSdcByKMMcXcehv5sgN9/opYTNaMe34x9uxrwT2Yh+15M91KjU8CWj
TPAJE4C/dE6/mMwiCTfiYeN67vCgmd7Zpm5Gi7MKILhgQoVdUaskvsigvP5sPkoX
GJDqjYkRgFLDWSnAcdn+66H4uLXDgRQbzjkT64PphRalXT9uayIIMYhqdWZ0lIMU
iGSIUrNavZId5/iG9WebEEbbaoIFGXsTeP2Uns+kpltbi5Wx4hHAEXy9AuZBEtLl
Ucife6bSlXG6XyUMufq0jUzODEm8LdGeC4KzYVheFhKu+Riezpszl2ZLP2i5U3cZ
MedkJOHT3KuTiC4KFaXBTuz+dJ5Xr5RYvxetlWIDF7NTi0BrAR+4uhxgrOa6vz9v
/q1FY7uP0qYRnpLQn7Fl0NcQ1GHA6E7BueHzN8CR+dUx2chWEhCGLTDG4NvDJSHz
zf8Rw8ftQT+E1hPXrPzlT+34nJcSQLr3fhIpXOg8PMaljNNrmmbXsUG85f+nytoE
Zf8k8c4RYZpcVJCh+Idpd1KVc6JbgtaDOt0K2oJM3tLrp31MjqoR/YujR5OcLF3Q
3G0UGRu5Mp5HscNELLC/3pVeGnh10jdjx+WQL4OUjnNEDTZfs+Iotq4QFtBtgJHm
uUGvH5t8UC9Pxe8fUcpaX/FNiUyyI1i9fQYGrwj+EJ96DT/9ulLuPhrqUo1sPwHS
i+DBPLyy27tFrSjlIA8zRzocjDqMDJxrq3LqlQuPKrRRHVcBTlQxclT2GVXVGMCd
hDHCpgFg+Zl1GON4CehljfFEIQrapy5isCcEHC49SnCPPmCRdlTtCaWZW0pvtgYc
y/9p1pmaHjL8btDNZK1FRrUGmYW/7dQo9DwgA0MtRnWsLaLYBn0Opt26YAUDLMwN
rzmyetqRa5jhGiYOBfsMJr04wV6YeXOqYLh00iViODtbk5P2ObSVKe4VSo/54oVf
hP/+lmGhDs13V7u9qhTENuu2+09DP9ulmh43Y5qzq/MrWZk3tn9VMnnWHCoV7TZo
e13P1//DKzZjtzZnexf/yA+QeS0GM8uWlZgGUuGAY9QsjtEHnnNPEV2yfpUrbULy
y4PmbpEsFtnQNcayY/89DKgakGtjh84tJDnAi4fSsfE8dG04YHvkqjMWDqecr/6G
xGqK3Dg1bLg9bFoVcCkyG/VOWDHbjmru/0htl6ICOj9TMJCbqK8crvyp+u3qoRAy
9t9+hr4IhXMx8IeWXb+4DiCLPJXW6ajkvzzDh8gvSE/Y5EY9R/8qvscUKQXdXLu6
S7P0+oaJiXX2IV7YYp4toFLB6ZmkRK/pLyosgu/bKE5Fdj+wu0PAJ9gOWm5l/V1S
u6oUKigUgEG24cqakO373nEsv6Iz30Rvtyjs5fiUTfN4nFhPjPL5+7sAmioEYgIq
YwhxwLi2XkoCUrQgciFG1jid8JXjS2cZZ6G8FWrf+utO5EciAPF3iu6H+Y3+MuSA
sGn1I9UJybW8hsv3CkMeql9xkEtJYfyagx5E2xckyGfZQh/f1ETx55e90289Szu9
Ml9NplsOKvu4JqR5C4oxP/Q77VVMfxxHBPb71xS4C1DzyYDfxfpy/W8SE7CVlRI5
zPgZ2+aZatwH0ywBbLNQakaq0ojEYx5zavD3B6In+Jkfik4J2OTwEgXUMGIQyV0T
he9TeeUA58jqxP4vde6PGS7J7ZwT+i/cG74J2x0g9b7VQHMSVTyYWS0xq6avlhty
QIwsggqBrqBQzQnCMUNs4Iyc2POnCTLdKXrMbsIC3YcdukyiTZ+PDIndmOvFv9+M
bVE5IwEeewoWZo6XeQmbFsHq902Uoq1livRjatUPcTXCGiGLOaVihkuHYJ13E0aA
27+M70ewwPZsdWHR08XFSa2IEWDBO5JDOjlQt7H4lQxDG38ew+qubqmbguDSmiFx
0Z17dZF0ba0oO6PTgS4x+dVzfhVcMPhA3/O/AIiAlssoWUdpeYct70tBZaLzgoBT
bZkP+q72H7TA532k2eEgZ1xCdeOKQeLdsKRMgPq52v+6Gykr3stqxYLOciCOaCxR
QGtpfxc/g4Xzn9gwyXihfQzhLkdcyCDQtkqEuP19X0QAhZURMINWrrbq9mBwzo+1
zEltL++VybVj4QPGoQ3I6AJ/s3J24S6dmfeT/kiYdQ4F2qoSb8Zb3bmY5UY0NTTR
icRKc7PlKUGNZVSq8XTG+RtYBcrrTuFqtKoJ4mEpg2PChgBZ0kSs0+Gc0vC/nAwG
6eT7Td+5On5h36qY+jcUs/mCw60N1YVvAZBDOD7vxHo5NQWTp0DCL4aGseZMqyso
4nS0eXKmBeJ2ZRT3+tFEMzr9Cw5+89Nu9sJG/fI/h+xiogk1yVHYv7IRDTvL9FuD
zW1PHo00dk7G6QGoxQ5Gbyx7fniPRl3KA8IFuRUeaTsBFXiUofyl3Ok31XMY3a+o
f9NwFT1FmInYivXId8epnYH5eu02/IFDsPsSty2PDOtVWalf26Yc8gnL22MABGXF
p1X4ScMp5jyS4FdOA25rzOvWKHi8uSeowE8swhSAv4I7+gIHNy0k1bjBtkdxXKwJ
pUqoJ+ptXazSDmumevM4g498NbFUFcxQTae81nLIDUEkjyYCAFndT6K7whm3T+08
jhbUDWPfQ6hUBOGRuc7Pm/xeCj4GPOs64Y01plYAeRiucNm8AOzJNPihtS/HutUE
0Y5xNuUzbNc1LKQlBSpVYdnnnIChiETzBHOBrS2TdQUVTLgLxWbk2/xFf2pQYqCc
kQ76fA8pPmR67Fc2s52NjkzDsIOVtw/eIdotXno/iHaMTbCEV9OzyjaNCIgoVZvT
EiJz3nmxZg3OPlPOHpC6y2EK4pN0YonvphYnE234Mbh2hRPe6nhb73KWGlKbESpl
U48Q8/SxsZp+stMXNF2g8tAhPBzBHHb77zcUfj9gipk7ee9ib3BvpOehp/eI1Km5
rskgnTqUI/Q7JQvoreBIUzUDiXXHLS2gABHzfrR9hVSwPKpXrtTSPlS5GbwZj8oG
q3lHw0rGP6YJj18UhfjwynLoxK01mrUIJOxQLcGqVUvlMmPbnTqwttDIh2NgQquz
amow0ltOGo53ltxZlFR8nZPnNBGexfpY/hFvbNKRl5aIlkRr+vwrjmFQJiWSlBGV
2/K6QR4qN+FZUIIYwk2oIigAF1vwqe9GbYZzpWfzLlV2lPdkU8Y03M02frS9VtZY
k6FjRK9+DLYOLq0xwr/F9dce1wGGvhqLKkzaazSX+OsuhNM1ptT6naf2bSfNH+U+
CMXc73qtx9/R03b1y9MS/0RdsvyClewd7yYRIyfmxS6ZXoUkwzFiXgF8GP+GTkE4
0xTUR+wfQ2kdpCA7CbZmEnp5sz3CGWLuHJRKmEf25tWdOSsFJSPbf8Y+dz0qQTgc
7IvgMlm5knoFqIxDNnbDDI4EKkg1UjsxqFv6KWf9saRk4pIOUkrpbmxl3Jov+M66
aG7V+ioDAyRhVJwN86J3SVo1LOiPwGsmvLtww7wjtQdDBFCJrJKU48Lbro7ODhQt
oJBkUltudmqUo4cGm/cDU1BQNu/hgU7XZqHWtxn0RF4p5hhyg+qKWDQUqUWeO1Cz
2Iw/kwn5OAiJRPcIQDib8pjFtOlexgMCXUVSZFory3sD4lrZol2SOFu1GUIPhsLY
JCkdUWdkx9XAvqS06kXa0F6gAWfVDs+O9xxsVSgfa48oEGKjgtJivorkF1F6ApYa
De6pqYEtis0Xe0ULrJf78tBoC5o9bTo0AoLvh5v3gYSW0T19uieXvnSTT14IuC4x
u2Vk9apu5HQux2sen/cgJNJuFjPeVK0nvkPVmwtxfdrypvWpw6oVTk1Ce896EXpp
Fj+wUc7cuGQuWiHfjI/IWaG+7rOTLHLqCizhX/QDCyhdQpmlfVHzdEYr7u/HNn04
82dcdyUTLVgTYXyiLl/XZ7/urGkrZgCUFdG+A9HxKH7/Pi5VJRlw7IUzycoTfOvc
NQg9SL47N9RtvVRyUMldphmv36rf+jeMUyPg5uXf6/kWumiCDcTz/JwSCTaaDck6
eBLJLiDmXFFLNAv3gQunzQU7bRGQdXJgK49agpak2xT6IXKeOC4EmfVmkw17Ypcj
5PajHuhLoDyPEQlHcuXrjUBcUCmLuoAsJg8t7NfBKtr1ag6A6ImmdrkqxDuxzAQW
ug15yOKQgS48bByKTAmUo1YWe3SLi8hweGvVz0Q1733IGU8ijRm1EXoYriOM7gEb
pHeVBA0nNKWmggOVu17NCNPr7BPupuohzdT1IXiHcOHHgYHTWm2gFxpaj0k1D8Hq
rihEbQD5eokQi5YLk11IWeNM1mr3LXi6zBFP5S9+UF+ufeLsyTltVNoBIGzKipgp
TKAnzcBW0+vb+A/oWaahJ7kgLy6D4AouozV4hsCuFLvRucrHRRX1zsRlPBUz3eUU
VMXZ9jZLBcYrNCfgPqf+QABQGDRrk09u/Xxvc1uUWjJLki9UKdCKWxzguYfMxsVu
D7mja6Hy75y9NB2/kV8k3Gs2wzadOSAQrz46BCtRWSBalcUtDXhTUEDZRQjy/A59
NKnHVQvMcOzlCBkQv2r80kKIZIVBbTPXFl3iqw3xf888/PnWly61gWL+n9uf408I
IwvPbvwc4um3MS+YrxWvZugx82pw7wA6bQkV9r+vXOg7fmsh0w9OaCWAbECb0u/r
47vAj1QLvrG+m4nh6AbUHf/fa/FUC0GufXyEPJybSfB1CiCDWlMivHZXE2150Iev
XlYTndjPhyLiCb0NOXIZx6ccMDuqYQ8fk5ypKCM8kkhDySqG1hQDE0QTC7e1CzS/
peW6w9QtYFIgp92rJdJ3Xuon/sEeN7Z0Zy1ZPEuLt+1MJ3A4FbeLptNN/g4izVto
LsfBppZyvc2V4oQGqPyOzIUGvl2LRrT8in83JEU5dR9gU8IHW4XhJTqEljrz5TES
vKeaECmXXU7HAzHY/sOUQD6U/8FfBL4zBpp2C5ZZs4lS04SYwt7SF9eO/AkhuLQX
b1sA6JZbKz+qhPdrJsDXFAYj/hSScbfPnjdM53abDJmCVkbj4wR93pVRBgCPna34
SFf3NBt35YXO7uYg6wY7UYDWCnG/aEC5CTfKcd/OxN4VOnW+KlvtTQkmaxMnN2h2
58j7kW2HhFjRcdpeZIEzmtX6Dr4w4jGI/jielBFq0E86EaKK305J+fbpetwPeuid
FOKJ2O8VmI3epqtu/cRBl9ThzQsDzl8Naq68ujzDj6c9aFpPXZFJ6Yifwk2mQA4g
roM1QlubLBXvPc4uC40RjEOGxdhtKU9iByK0J+CxVCU+UozV3ch/wes+Gn1rRdHk
Fg7KzvRxLH6DnTvvHo1D+yLTR21Zf0xZRnRUX2jPHv6ONhbpIwui5IuyivNMPDF7
DfjbgwIbeSJFtNzVuWXFDkE0OQu/lc3KghIFoCuGl4eVgTXf0rhGl9UelFFMxvpw
6OYGEioIGT9m3bIWA4GmqW25fe5VBMpNGJLmUSKtCr8wUcGQ8UcKbQFoSqlWsWJV
S+Rlw4FO39rYbqWaJ7uuHr63KDsEpDc3vJxXrjAY2mm3T5wUAggSR6YrqlqG2DKH
3IQWKdG3j5/vdvCnmEjld2ATw/hDTKWLCSbmnW+r3JL1zu5TdIsVBlcFyBNnn4b4
ICvXNGuoLL77tByNJdzTgFA517dQA+alkWaSO5Y6WnFB8JRnc4q7KGAv2dt1Iysx
M+RcQ7QieispZrf8mpCrBOeVf/Ns/+p31oQk7d/PvgaKizQACBYQ4UlBW01QBcDU
RWBp1RvmnRn/fFY7wPcxKxyvLXmGpBGgyjCAbHvYrN/HsyeuXarnKzMT+Rww6g00
ZnPDdUKfXn6sZMHnRPiOQPYJ2lPWuHLeD7wYcdUJIeD1bKzHrgRMfCVNyxIT9Vqi
2iHRA2Jygg6bIxlakhDvykioBemwFzbvdMTctk+KlOm0fkibuU5myA2P+9HJ1772
S8yFMFuM2tfgj+QNL53y9uKivuMP1NWfUlhlySNdFupxC5Cua+kbqPYhrVomhLJg
Mi8Thp09vXui9pvB/acZgkTY6VGGDxyiyQNh0gnyeenNI48CO4IOnbvSVb29D6Ov
o//xfPc5iB+pWwE9p+uX+eSgEOT3D5mt13JFlxqVMgCgOjLXk4AfxG8EotP0nM/D
wXeX88rgN6KrjvrmOZRVL4lIkuPwdL3Z0D1AlPioeiPRy6qsFDZtcZl7iu3vXJmA
AQTJ6cp5Fayoc/BVD3x2xBRyvkXQSqA/hI027Udm2jiMsafZTo+nBIrJ9bVrZVOC
E6JJbMvCSGI8ZoQd9uOj7GcipfLV5KbURWyPNiJrxPZv1KD9ih29MB02PcTj8Co+
z8MXduMAr/Hsii/thy2ScZ9mE7/I1dpaDYzJQ+laQ+UQwvak9xPl6aQdLFoUabcF
xnBeqZv0YNqPQW1N4OyNGfZrmXQgyrJRWv2VNEEWdapvmZ+vXmNZ/sbLIqRIugdE
x6A6SpR+vTUg4/tcQ1IlLA/afkXw3NttH5Acz6qD6BvGT/+2mPr0FXPnGHVMCQEJ
w7eE6MI8GjAHmpVH6Q90yP3DMhE19LzSvPmIJKkh4wubHPtrIrKbFTs79neFytiw
LFvpibdnBmoyy67YevcB/iNiFioxh4DudKOSID4ra4wesrzQnN1eoWOKgs5V8CVW
iXrrYkw2PjxGW6DF0F6CatolTss4Fp0Zv/2xl3IBPGAzbPsPi4i5OLpNVbGuC6Ej
9pXEsIFL12ANxdGwnQ9wyTy+7/hk4eOejzjW70SWPmj9F2qw6n+gBL57MO69ap9Z
dAlPrxt5hf7QGqZMmos16XEh5KNpF41qj0w7hEeWmYsi3YBnD3pyOa6+SLKahCGm
Aj1/27LTeoZU5NR+n6XZ1J0QYYg1/kesy7qKIpVwOkir1KyTDeG/h5uSIbsoAHV2
U/uS7lc+EQEdkluKKP37lfectQ6b67hdQOOthmD4xHivbRgRn5xT98omAiT4Fo5n
/YI3BtJBG8Cv1/qWIJkK3wTfMGqo5+y3IOmIKuCf1Jfoseeb3WuNFWGuSnCwS9PB
UuTPy4Mx113o5GvGgZI4mQwluxkbFGx9zNx6Pj8Vs6+obHxZ4j4aAjEB7+J5dJzf
PZ1cGNgzwhcdOhYd1kqXB0bWoOPnuGLNVPo3waa3LQR3mr57e4AxRFUG/BfOjyJ+
vz39WENqjjHY2264SWEWoalOXLEqWlEym6QE6FN37g1J/uratqD9S+eP27i38Rs7
VPkKHoFCeuBRW0ULdaCf4g63BGOeB9sV3YdOY1I0dcjijLaDtSI5ZmdNVo5RAefU
EOCyoEPsj6NUwJ7WhSe6G51jtSHCVdfvhMgvd/ftwEvY649gSAFvM9nLXYkun4gt
nBZux5ACYMtCn1KzUpGtHT9v4qeAfIf1xpAC87+njItl9EwbQuM0HKKFG+Txdypa
8n0pvu8XR57mWBFBqQ322IcueY8FRyojTUXyN4cSVDhTwYSbrlUVuGKErVqcqKuA
auPG1HGY4kxUin08kpkxZxWzXF3xkJzJzpe2B7xsfarKzGvWM5zxwGnnTGrBqhaO
9rqC0UpcjzzPPHjq+Wtd+46yrsSKAAEjEPLZ36botWv+ZpEIM7xJowpe/TR9KdF4
UEXLLrJvwSCoGkiiaFN/BnP2IqqvBElpQvVltn51cjPNJBJYhpFbSgfmJGbgb43c
1jkCWeLde0bJnU6m/4HFQ5e08xbRGIoYd6U7IqiAG5y20bZBmYrpZq2lEtLsed1y
Hlrnu1oP+mWvRFvA/2IF0D3OumlNZ4cLk5tERRuzuMaDYkjZ0m56QYERIMxMChEd
vlXucOGu2ZygR/hyYfqxpBxTxFnIkkPw7RgfheKIHv4r0flmh1oYe7uePUkeZtEl
QscOQPTk/9kxwvLaZc5iylLQWTBc/CjSO32jEEhwV5fqQvOtwDb1nTyv5RU4J+ME
7ICO371XvoIUG2tDOqPey+XNGmb1AIOodaBeaoYd2F39buWVG6yQil8HGDNm4ah+
59NhDwq/7JhcV8u4z2HKAF+8nZLeJtAtX3TKgu0DhRQBxFgNywmn+ReKtDtPp2Bc
5mZ0+vB/4/feaTDtG/1G/plW4EjFZwIoqI7sdhaxV5MAXnPpzT53k90tfTbXnArp
AHefxEDbyCcBiM+otS5gjtaE/KrLPy12gJtVpWSEbwcUBsqngFEqTBOWa2CSqwXc
VSkFkr33u+4hZC3j9dSJd2BqQoAFjsLKuZaakb65Y5K+OgO+Hkc7G/G7cYM08tMu
T1t5zMVmrVmlsGm9T4nsGCxWDR6DZWVNJoIZl6mzMQiY56HSrlB2zhxY/t31rpIi
xLzVpjZ6415C0ieKpNaA5VkDGXCjg3H8kUiUDvjbscxsGLP8gNo7dHXikiV9NzN7
HcCAAt+pc6/7m2R7sPJXSSgnv3xho8LC1Okgmye4WK8bXGHwEBwHVxllhZk1TjL2
RSvWKujzMEP5f7cQhTrNLlt8K2lySBM600CAZMTTtN7Xyf/U4uVd5BC9IBHJyOH2
58vHeJdn2cArqjSfm72o/2Pq5wXLmjXCzLQqzilvXx0C5d8tIfRO7WJcOqGLqrlh
J2461oef8mY1BJIIrmlqbRZqwA2oGflsn3B/hfBG1BMN7Y6Bk5fThUcd9qgmCCbX
7jdMmmFcXGdAccFMpypXUwjmWtPfZ8WCqNoXZRx1g6/knQP38cVyKxZZVO8dpY9y
3ioUemVONp213HLyOdADS5Ji9qo3NO7/whGDW/Dv1YP1T1QScFaGHmn8OgUjnNmp
Td5uFy1y1P8nVYBdYsDLJO4RpspBmu6gqpWPeAd7PNsMoH1bTuE7RjqpmTmOKgSp
GKeRpaaChmjJz0+rVnMBdVf2TfT2qn/GADMBKMMZIzF5fev/xi80kX51SzLiINb5
iWCzO5Mqow2Ar6jUoQniIn6aeLhBE0vTmdEwn1l3UnkKJ6WNHP5585Vyw/UAEGK6
OwpU4aEk1bkxRVyFKaEFEhSdmstp2WK0/1qnMnrEdQvVGMRzR6NfYywCH3yWahCw
qdAAk4/dh8Vok6JXiqwM9+rWFtJeGYKhEgwqb40GlkOUCTJVdRdLFjrPt5c9YJd5
qKuQEOVHcgef7aO5hzeFJ4ilqwXMUobpced4H2W44n5nudaOK76z/TQu5nZNbrRv
WisPrK6egGzFwD3UmWkTGk6+gJd+uAeNag2kCjP3x3MRkJe5HqeEHenUpGOSUbKZ
09d6lJI8XZtn+rICFrPLfej/K5XAXwoEtGSTevWOIdWmPgW9HJa2v6HRauwTMrNg
CPk+Eel54cDAnSwDR263cQA1dwc31DiqoQplN8zAOj7sBWwMRXHGCX8Pns/KwPR0
6OVnPmPX2oGCDLHu69J1kSi7y0SnvqekEVtIsxNM6vXGlEEJqgMh34yCkleihIWn
WPOCA5BOi94eneWzazBZ7I7lvmv87jnCv2t9T91QnBPO2L09LZlelSW56lrdGaCP
k+SZprhJyKoBtpUQTj7qV/p0jSgB7KyUl3oRL9QOyPxGAAcODwceFSOO7gX7JF/4
rPItfkkcggsaiJ3mtJF9zP0Lb90om7ttcSKQ85LAHTJ4nJVX24M+EldZj+JsVhN/
eTRzlXY+YVsXnd2rnbdf3EBT2HaBQaEyltlaIgseHvQbDcLNV2hVnUJwbikOYVlH
Lk8zO9aW+3Y+7LWdAbSRkI1h3SkoWZ1uNXsbK5kn7/oIgkZrbsFH5AGW6lmKMSnm
BhkNEglVTtsm3zF8IBKDaWOEFycvRdT3w4gJeQq2b5TeitZU2KqoNdxGlIGaNoeA
/2WtWiGyq8Gi1V3ohXyAzZ/SgRoR0WJcwsbBssPMaTeHFOFRityyojUSVRtxWmFa
tvf/x6ZF2HMedPYSoPR1T1o/UKWeyJW1q1H30Q3GNTQBnODDlKaOdiCn9GDsLd5M
cTzSYzK2+o25epQ5x7YZfEN4/neJw4KsBZvvt/Mm5Ig2vUXsc4gqvEAnt4z3hBAZ
LOMy/Qwl8ps5zKIE+K1DdbJcZU/ppzWm7r3ecmRk8PcRRE3fzeYuYHFE0EzMR1nC
eRkcO/PD6+tohzkbMeZqJxKnwq0GnKbiqOYpL9LkXiiUp4f2Pw66VMua/Yb7SVgb
equeeWFBLR87CEVWK138pyeCZmm8pjeGseZj/U3zxutKfC0Swe94g66HxTUbtJwU
mmTl8/rRnxTmUrqYIRUStFJOsIX1Cyx7/MGmdk1pGU97pzBuB4YIkMcdEfggrH7Y
tULp+i7q9zESMM9VsL0HRvH/qecC5xQgRmMJIut8Z9PX4QErzvrYQkZxxypO3h88
cqzHjZP2z4uo9Lwci7oy0LFyBM9PF64aJckKPtQzjORQtemQmOl27B83J/LBMcDP
HNNPm+y4BWf+sAev6AfJ7lQ0Ku2GQlK9OYOdvbSO3fJmruRR6MUaq8sHLG4x7CT/
OeuoLU3nZCn9j62wq81e7YFFeGmiE6ewdG+R4nvABU8KGXxHme7tsoB0YbIuR9eF
wqoR845tJaMgL/dsWqsgRM23gwYFmWW8LMsABuhuZ7PYxxlGFXu2NsYvPS83Dfhh
3xuc1VXWwvOYB/lMTubjkOBwQJDPucxvQ+0uIfcKgrYjUgPKsXUgJ2w/sZXek9Hf
E25GSrLgaBPHVpDtO5px5rkVwNo8vg21fkH5AGYy1IQ6SMSmPbf9+8XuOX80Vs4b
rkwciiHSKDYGiFOBtSCNSUiMZp6eQcHZ8TYQ2jiaLbQahrA3+i3h84RcY9mKiuIz
0HFlne+22sMlwLS0/39jr09mmFQYYCNigHZl24XDKsCnehgnAFDvMlIFTRIbDiTH
afXMeuf9BbLuN1yHlxdu5rh649ixycIb9Qf1TksjxfhWJhOO1tcsrWpgqmyiIwrh
nCtinREQWE9TzbDKyECHh9EgnK8rwhVm/Z9hL5sqWBPMg58cVN5MsAL2cVdV4lK/
/LC4pU6HHQgWY7N/hoaZu8Trc96Ubivts2gGOM8qV/GP027jR3Vg9sjE+bE7tRIh
ol/aSQ44Gpb1B76zgxn5DrBHLqJj+OrXhb5QpB6pqPy3/W9jMpVJMY/o86ZV9X7s
xUf0otIPaveFF8N9wVCM4qdVp7b2RSI90buk190C+Fj0RNRFrCivU0QjSG+5ykck
k+U20MdOpoBRv9W5X9hdyn+gjmEv3A6U+FaBz14FCz/zTKFbtX8LfCKj3+P2oKs8
3ZEQS+ELblr2CvceMQivxE8SprlwQuBeVSqKOknSfHj64RkS0pXDZKnJOoTSYwZS
ZMrCnE9EHddJIa9pPlSjGmrMx98zCT0de0uqcwIUDMIvTKRpiYTDxEwgMqmJktPl
4RFUnDbKR5jJg/S8zf2Logz0/0RAXem1pYJvofhveSx7i8r3e5h0Cczt2GOkoc7K
gM+zZS1oy4lB6AFdC12fTXlYQPw97AsvZkzYr5LjuBBd9NQhMZVNhI2Ssuh0wCQ1
O8C/nDUl7Zth5A++XSvGBci4bIGewsGKiUZlHiBPSGX06V47CACf23Hdptue4vGI
Wps4V/sOMdSaPLPyOprhsMVRgi23CXpWqYZe+aDBpa9giYj6/uS2mgFciVDqYUdK
yqnrBGu7xd/8PmHIuHSdmFOeK2dCJHthEOiXYDbxIVAQU/CYow4ZTyn++NUAba7H
pt/GquxeqjxKYSfebErYD8h9gPezJ8TYytmQp3In5RQLIAOdmcLArJGgtXq7063/
h6y8fIrvt9ILNc0n4f9FNIRgg9apGJ+s0KU/w3wI34LoNWCRL3RO3R1hy6mnS1sN
Zy1b8YfePP2JiytA4lba2D+NgpxgsihqrkMzbTPMNVjczxx55CxrfKpKbsnjjerp
3wkIQsshZamSIP8AK6uUBgNIpTxsg5ULLkvWCM47+KNdS5j8uvsyIrqdRbXI4Rx+
dOzzsb+hyxkNzOoqUFKvUK+DXmpOCZYoLYvsmv9dTqN5SpBPzwWoPfrf2+m8cbte
7ftrXUXklvZlKm8JnEqyzSOj4rTcVhdFkfsEyc8xW1pdfT6XYAumueiRPmHqtkjz
QdUM/PMvvfsVQU2BxSgKayf18RfpQA+/NoYO2TlGAFtG3xYN5cQW2+cVJiKGeYtk
mmrW9zbxlGX/UfcshOuZwUjl2F2Gkph2udLid8vwP0nBwX8W9ixUk0VSNRR4oYGO
mAfCv2k+ieKzidrpC0ekGit5Leh+3FysKXsD8OgvHx6LMlTsnRRE9B9Q5hJM3CjS
tLTsw/bEGRaLQALJ2d9UJy1Nt2wVTAYqO7aXAYFwr6Mp4wv7oXwVEZ9dbVNzLprk
wd96yV41rYoVhWTbd+cvGo7ZV4LtWWAd2ioucizGviS3Z/PMRWWvpVlTqTx5NZg8
dGT3iDdDYoEhd0gEO1Y81Ami0CIwzn9GqPdkOdBcSd+qv3MyHF/4pyy2YEYAqDZS
KMK56fDJy42W8Wtkb2xWyLe2yY6cdueJMYVD+ODJE+nZuGXEv3zFdGOqs6pQBWoY
UU166dkZi3diN1SWPEJV/QFfOm8N3QDQ85sepSlj9dk1kyKuqGw6NYwFh2XiOMnm
AXR0lVeVCchD5Gk+Od2TuL2WS1sOnRJVs5T8szLk2Udr5fvfHL4D+dOpleNu1xPM
8RdJoYHEMjC6iIk3kJxMPh1ekg1wyBUPOcyleL4MTIxyv2ZoCU7q2zY+uveaPvde
oRnhv48yRcYHKiL56KLlVjHYbQSMZ5v3AomxO5QKXJiFbc5KFs020zuM0Laurnjj
C0rpCEfKgN6issbIhCeFl12PcvUFT7AqIzuzhifV2PxmH5yzuFBNloArh5tnuvrc
devgq6hholj3fH25aeDRPQThV3TAsKImJ81IRi6kKM2UBjM/QRrUMzk2jBt0pGzS
rTadUuM344MdToexnJfLuMdb9aKO3Sze5d1CAjTt1gIUpMejuBWuRDPqxI3hpZWN
khM14v3Y/l+BFhWw4bWH5sXP8jfP8fxHZTKbDvrfQOw5tYUMwjq36hHE/5MQph1r
jSRwD36qs3rgYDLeOFm20qsjSoZ6EQH5n+u3N4/0dIAy3S1j8zwipCJYi+MOcnK8
RZ8FYvX6Rul8/xlFiBLHnsKKOskA0ABee0YrkV8pjnQyLorTesde2YibCox6vLSu
/5r0aN0iM7DFVpgVyQsJoyfMN6HkcFGouDQ+f0sjFrWa8LwQ2cy6TKZfffFMLdgP
gClq3GJhgCS+TFeq+3AqfU4/pm9Bu2w8izQBDgKsLaFUiF+I0GmFiEV+38ISKvSa
ESM4VKamD4rf281OKkQfiAqDiaufh9vonqE4vKfGvamkNb2/Yo6+GkAvofQBaSFv
s9t8cDkaPT1TmTpbSKdD5N5gg6H0L8SDo7rV3a541o845nJVZm3snuWYgnDdIAw0
xgKaOmpfy3jDtRKszEforHIzGCoa5rqHRzKfISGwOvRJww/ti5D9N6R3uEwmVfD3
AEGDiDDTbMjU1rGBY9zYE0JavGVp2wn9aB7IOYOVZ8lkW+Hn+4XbC8LjmkB4J6a3
p68gIHomOmOSDRHFZ5B+fQrOo346NxXKnIouVrS0W8rpP4c5hctKpZLuiwzvyJOK
ShVmqY3W9LkVdaXTDH+MIRCiiQhVGDLAT1GGeFZFJ/a5nN4H7d5zyod8kiaa194k
9QJ4KDtRMXvlbQ+IV7tx+8FI6pZFfVFwelryUiiPsJCRGK7ude5V4u4sOPNwJ9AZ
n9UIQG8cdgrxCfkASYXu7jLFV9XvLKzRab9q9I1TfmzvGBL3JUqAm50itDImFZsu
4Rblk+l3LF/GlYoaH/Z4liCAzocf96Ly9fNSMNX5adNw0eqh3S4+VT/SiySaznln
naX/kkKHCVHbfc90YL1q/Ar30AQsHoPI41bQy0dGSRlHfDMe4HAclCXi2vKWnVMq
FHEoHRz4ojRwNAghE2iYObqCkaHqMQPN2sd2GcNOFJkyuAPKS55disyfzVBBCxqa
+aROwID+my2Mq5V1HcRAjqNZio9TSgi0iK3gQnqVyf0j6OlO0qBp8FPXdLnXAfZs
ERaUjjfAcjEX/ImWlRBYxVvtC9Ah49V69+z6s8sm1XMqTuDEwvK9eqJnH0STXASz
IcOvdsUliusYFqXWLnWTD5Lk9s8zRyLXnrErIE9vdv3paNgyCm55duaCMmnEsGQd
Dt/vpCvsutLrTHGwoiCGgrxnOx9wCcFJAJ7xGuzrz+1ByxKufgCReyJ/D6ms911q
LMjQVd6BYhAmonXkMqDJutE+91fMcVLTdIVqVQet2R4l4UGUxPPe0aM5yl9ghAlv
/mL3TQ1Lykx/NkizcucFa8CeulE11+ZbJQWG1d3slyAmn2F/kQ//W6mH8aCh1FNT
RhXraN99rf6X5qYKMwdO8CfTB9ebFn/tmbQI15FQbP057iTX1fyD+pTL1xMC5q7P
42/veLpa5Odbj/yfXgfFBKbgt4yiuCyJh6ZbLoxEofrscF2mySCD8gvXqCXNQLvJ
c5CN0L5gHtt7eAgUYwDcByk8JxXIHXaZdhUBLCePqMt8OBcSOXAiOjcngA880qqm
OoySsKHN48ptihXRv9hYFzbznyyIr+ATIyKihWj/cX4N6u6a5egoiPEyGT8alkLH
AXahvze1fUveEB9ZagBzICbuPBBkTQaH047G7T7sKIi+M4bPVXjjuO/SGWOpQrJ4
BtBuDwjazQ8PigriBX8CyAQHc9QW8/mJuDDQq04fePV8sCW/ZchICZBS0yjqRPRE
cqR0KwzMXJzR6AThlxjD3aiW3ByEeWPAXWMMDdBcjkE=
`pragma protect end_protected
