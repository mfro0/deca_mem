// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HHEW8PZ F7<MW@45>57UEJ02J"=;)5;^;=<JRFTHM<WN^[KQ G_,)L@  
HU&[QX;^K]&X&\7>/XQI9*\8*M X0=:S0/!T<UDYHM(#<RJ*'A>FZSP  
HM@DSUV@"X%UA8R ,*K)4?"T%K\LW-UL=+B5D!YT)&'%('2CL1\:(*   
HE9CQ0I#\!,_2TY:>CEG)&=FSJI6HGTVXB"T 7G@=T6]EYV<N^[\=/0  
HT8$0N1V);FVJ>XOU_Y3HJU"NL9'!O-M2F>46),R[?G3(Q>+5:F)]%0  
`pragma protect encoding=(enctype="uuencode",bytes=19536       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@(RN ^ I]'88&K=%/RPP6TKKZ>I0L\J)^-K'B43*Y%'L 
@*CT6N=TH[V\ K4PV8UYANCCYWFQKM])XDW:5ZRWG0]\ 
@>6[RE5W4H*1H9 C<X0ZW@EY,UI%S%!TM7WO6!6,IL!D 
@.J6+?J1V<EM7U!P9!,@T9Z3;FK%"L9+5@/;V (P/P$( 
@"_".Y=9=WIV\\V$?2'I]>;^L;N$D4D_][()7.'RTN&@ 
@ VBY.+%LN&-V0+W/#'FB#BE>_-OE2^>.I?8DOQ#>]/D 
@W!G[-XV06'A68QRVKOYZ]]4C+[\9+[#0M3Y'C#8_<LT 
@*8E %9I, :&:?:_RC4X'<VXT&8;XBK)&MJ9L^I[O->  
@QP2P@X?(B&%J8;8+>K,BV!MN8V\27?C>C%DSTD0M1P@ 
@)Z.>6#M!&@T/N<RL=!I'FG]Y0"6P&-8>>"+.S[4UN?@ 
@A=7+#_$4Q@C&RG6V88,P8XIWT_J;S+S1P@5FHY,&X[0 
@R79GU,G->J]1%+%/EJ@*>""P9J_+%;$+[13&Y<<9Q1T 
@6GB8[\(;D!^4/8?"&/4$[<-5&WK%<L?U0U3K:LJJSU( 
@F;F?VEX3_2GB0DN=%@F)U"ZP>.R?!I;B2=*:/<[*0Q0 
@,>_)ZCQ_KA:]9)VR./H1%L9$)Z,E9W_DFZ(2:X@H_(T 
@F-DL[E7F%(T:E]HM+MM%(@H]:<E^=O+]%4L)^(ZO;RD 
@/ROMP]O 1*(I4TBH]>^@$J-"<4,Q=W\7_[(?&&Y?>@\ 
@I\V;59RNL\2&7/H>CJ6_MU$-^+)_@&,Y*42=6#0XQE4 
@6-/"_Z8MY?E3=:24*XK,Y)#BR#/H828E3]IKS,WCB(T 
@7-AP C*N3%#\&T+<U3@^9 :UCW0ZQ:; AL\W=0 ]MVD 
@5D9S=R2^G3XAU^=D:E<2E4:3"@-Y.T&7GU<] 'XO#W$ 
@*Q-!%,ES?W%G<'Y4EIYL9$RP!8Z9%CQ=>@B9H&K)E]H 
@2[V3PM,33A'S;0+]S'J+QX=X$1"==+050=BENWK_;1, 
@&\01)+T#=J<=>XFPHW=C1';@,!VI>"VCGB79.)6$_+8 
@T&A(J .;5#3^1QBF&Z,3OEN=JP>5?B[J8?.U)%4R_.4 
@6WN7V35<VOM>]ID\+N6*=*3/$8JDL*3K5@.4QK/:75X 
@U/T>S(K%SDN;JC]!D7@F8PBU >]$<K:Y<0;/ GW-=^$ 
@!HOX]1R:#YU'/T*2GO1EL8)+"U5H/0_C6.;F^K5LEL( 
@403U!M.S6[WIG]5+X2>"_95[ 1+80R>'[\3@2-4R3W( 
@S*C@<*][_."A5@"K5X_67?PA\[<AKB'O[6F"37>2H?< 
@>I9@;>LS30YC1S!M%8%"0R^&O)0PTQ5"%/=%-+TZZK< 
@O0*;XC &&6\O\:<\/D_];JE>UTE!F@!:7E2]_C<?=B$ 
@]M=;W=\&4AY?QL;[@?-^%DY(SF>+]END%/Z_KE!'TYX 
@%3YB(R";B_+"*M1B/%?+-C\_Q:P4_M6ST+Y%L%8&V"$ 
@S HB4T@H6A8A4).!HZS#'T[:1+]NQ;QG],.+@4_QZ?T 
@SBES&>UR0VDIO!5DI MIP_N8H?3';AW8K==B$"-@?#@ 
@RN_MN[02C4&O\SP\!^W]C99M?+"EL90$4','E#:9094 
@;4;+^2]GE>0J7X;/PN+G29H$W@#+BX;N:(66IA?TG P 
@?CRGK1_;(!->W^VWUVO\6G0G[_=+$-L=C+8I'W79M<0 
@7A"]N:ICR5_/<%NAJ-H%L;9F$H:LH*N@I.>]I)IFRWX 
@AV5,:$77OW./>J\ X".4ZI!6735/2<CC++4S:PYXC&L 
@ H.(Z_^[!9 U]6%; FAED>,WA2W;-Q'LW4X=[$FUF.< 
@!E ;U%?VU88IH"'WN^+W'@DVWVY=7<SEYW^O@+=?9/T 
@U3<K4!HHAY[^M 86N%\9"Q"/H\T&_/JFV=(TAHLE>N( 
@$>I?0$AR.2O(ZYE<='[%?=^S?/M(JFG1(.<6X,1&;_  
@JF%W> ]JCSU'VB7M^V<;JIHN.%3ULLM7M!K9@FK!1(  
@P\H,_?Y+ I:SO"Y*$ %X'+07?N(F>EF_^4EKBZG?C>0 
@C5:C3HDY0AA%/JG]S#/D\TY<:R"X=_;%9,BDS5J]73P 
@@WJ"9%A.WNC>4=D'IFM_X?YJ\@'A.\RMQTP7$NE53M, 
@ZBA--EU\]EXD.[+YG>D%F!BM8@3Z3.[YMY438:7NB1P 
@-.A;/#DS+E2[1PLO+(+.C@6_!#5IM0B@TB#!31&E;,$ 
@9GL%"-U#P%1F$E?E?HG> 795\,/,66;1 3FPRITT"<D 
@WGBX#GX6AL>(XTP/Y7E_E6S?20+3SQ<SH-* F-%A[*( 
@SAOO\=)4Z%UX%/[_!7>T]^$8=J.2G<,:PRM7LF4RK!  
@C%<GC() J $.A?&8!@-E">S_"DO_G+?2-QGNL2A?2'T 
@.1SM((M7P7?=&4[GI4Z/B"/\\$"WC!=,W.ZI,J)GTW0 
@Q0CX;'/6O6K@*?_6XG*O8IE(GBQ9?<O5M4*!/P PPNX 
@CG18)./[@NS"%N]>-6>40,=.&20]YO@7%=_*6:NHG'L 
@V A!#1W^6WLM;K4%Z[,M&0&F[NBT:P]$_I+;1H4U$]D 
@0W[E400H_,(D;=XY"[0W]C.Y\"F$+:[I"3*[QERQQ.X 
@L484>_*V1XVZB=</_#_UOU7W01S3T0,J\E2E)AMCC;, 
@X)-XKB1/GB5Q8V>::.@% 9/\DQ_S8T41HO0)@RPUM \ 
@71!QQ\[JLX4((E!G3L%T^5T/8NC=T(C#=+[H['Y4 7\ 
@#%& V#UD)V;_" K-^NQ(:K343F1\3W'6XQ/0JT8].<T 
@?N%DS$=G[QYBZ4D@,&LM[WI7(E9#I;D%"T6C:G*!WE$ 
@;-:$!;F^'3V\)E/!F^IR8\RZY^N=R^B9/L/@%/)=]3\ 
@GN DJA26=YB[E5]YBRE8@F$YUB\]>P*$0" XZ%G 7[L 
@PJ2%%_82KH JC]PS_7QC7D#P?1]=@7SMPU=#8*'C,@H 
@S)V:Z0YG;_H;U;K(\:>W*/;7'IM=D&MP59:+M6679&0 
@LL3P.GQ@7AM1WX$EN-K=Z$(.7KC JW((NJSG92WB;XX 
@+PPHE#RKS*2DZJ]C@1HZ+M+#AY3\D#YHS) 7DT1?(DT 
@ \=*NQQ[9'\ :22J6Q8I*EFLL(+X%<8I"D8Y<EI8T0( 
@QE9<]8T+,Q&&9A,/35^$#TIEB"9+^A:3BWR7CY*YN&4 
@U"M[W&5:-AI<6&]#2.G29O""\2/$2UUY[$.:U&[Y1=$ 
@^!2FFO=HDI?$2,M:R3Q$]X .68Q2),2^!RO8QP7N84( 
@##S<]N!/L2Y-:'CW#!,$ L4&:(28&\Y1P;WD>&[M.JX 
@9<3KSJX-9SAZ,=S?MQFK$ZM^@:,;+03+J$@OP2U[(?\ 
@,K([MJ6L((H_7JV;Z-V@2"L\Y8M_@EY6!Y7J0?OM($8 
@/UCW511&]TS8$46Y(==.=!13_.@Q#<C(N@N'!!@K<N\ 
@3=6E5QR[U46-&1^^.#%RS<4BYC-^',S !43:O4AJ:%< 
@L.(_5<M9=.@;C+^5I/J.Z>2-!ETD-D+I$ 789]4(HC, 
@H31&'P/@H]"["3,K5"8=L>[=TC()^_Z9XY88QSW:7IX 
@&0)U<KGBAM.+SK%AO.=F]'CEW1;A<S(='Q1_5N/$=L, 
@FS4:!1RLG:VG&U/"&8[E"AG:@00!<F/0ZZ XU?0WV7< 
@FM$CX?SY*)&^I;_Z8ZH8%EV>]& 9M]RU[8?LL$[R.9\ 
@I$ME*UX"--NAB.-R@I@FVU7:"^9@J;<EQE@6G"=-4P4 
@0BX6^*_5:4V-M6V^\FJQQWX?/$1QQNS ;.C':-BN5X( 
@D"67&D!@DIO60$W7W9]*@]4F5G0_F/@VAQL'W &V_'( 
@=QX75JS)XTN&POA<PE:G&V3MS_"P5B[?7^2G/2*>_;H 
@=D(%?U_V><U/P. X0<2)_;$56N?:V#I'6[4I\-I#^&$ 
@>R([B!FBM'>RG'V:+ZTD0G22K0>:?O>*[,=:R^H"^+P 
@<^PWVHU%[@H3Z3 G3L43^/23J:&JHTG1M8GND=A!$MD 
@FQ*J^_Y72PSKVS(13CP;L."^7&%"%%*O]M>(B(I7'L  
@^-^C]:BTP58QO=D>0Q1<E];JU/S]B2-T^#.J40'NW:H 
@F?GC"KZ.[DS*U>3W@")N:/DJFHHI'5$X/6D::=%QXE0 
@3MVCU;9->\8;Y9)?G3_AMKTB8T%7CN8NYB54=17)LQ  
@]D$QF&2!2=;10Q803@5+?1164<!G)P:UKO2BL29%"6@ 
@2<4X0E UG\(9<>8Q;G"I<E>LXVNRP$4?7-^J@/"$ N4 
@8"D]BWXO8&Y,894HCRYQ+U/9HHK>H(HT] ?:4 ;*;.  
@^%9LXM'!YS3)IH$-"!"@RZAO,29JM(3*SWOUW](.F54 
@/-DL@K).""L8T!@4;?U=\^B(O]S*7MO <D $':!+NU8 
@X1"2I$5LC<PJ;NR>B*<,RH: ;V</@() J9]L3K,74=L 
@Q@+J.KV"K$N62$K]P!O21KJ.6%S3_,3-N;UADH0L*%L 
@[:09[43>K%I,R8HG"DV)[!,6WC/-UX]T*O< YEI(4ZP 
@:0SD"BF=V9-E485!/'SR+S>WVQ82B.F#[57DL!^IN2@ 
@:7I^P:'_F)[Q?ID^6+8PG&4?<A4(9Q)T,L71ND;IAD< 
@H%PN<&4,5_D)Y0M8#YFDA1^D.Y&I:_F/Q)C#6>\O9-H 
@:DV>7SP0A(S9%#=*N-\O^/LB8:JO61[DYP42,^+>!H( 
@$\.J]"'(.H:JU9[6T,U-FXA14>X4Y1GU)(KC)":WU)4 
@KQU-7:6U>_>O<KYWQZ OQ_RG1V\L>/#V+A#:?*?TA#, 
@UV86^TI,UUX"LNY<0[0UL;GH"/43_Q\]LQ LL=O13IH 
@ 2E6-JQ/_>="*S";B%Y$3EA&.<M7VYA(^91XW2%6H:8 
@HQ3HG3319"I##:!)%<- X"\\BF7$8&"):OS2@W46)G0 
@4$O1 CH;3-H=/(8CR/PB81?R[95M^?.55@C*+[?H40  
@+]]7M,AU5EFK%D3X%G5R8;KY==!C<\4J:<F#Q[(96,L 
@)'?8( ,P6:LY]ON0P*.9?5WEQWJY@'1XD]-+B)QV'%L 
@10 7<BJH&!IEIT',MG"&2 C[2SG>'3&\/%B6O'3^8FT 
@J73'E&,L#K5?-))G:)O^4P8FCT@L5V&;^K @)L2SJ$( 
@,B.0Q9E0>N9SO^^VH5PG=DR04$- T]9M8G@$25^P'UL 
@A^.))81$LOG78RHG7O!4"S'VPG,ZAG3^*N8N6MN+>K@ 
@;\T]N3\@^H^ 9V' .#;RW(3^SMF.'MJXD,XN'\=4)A4 
@62=,#; /;Z65))MYE\:27JU)KLF556MN@!ZH[U::[IT 
@^!=]L=K=FD85VKUE&<X,MH;)MST__,YA?8:3+VZQ;>@ 
@8:I!K'D6;WS<E!.HJ!#2AY5+RS+?^H?QM(&:6[7W86P 
@9'ZSCVB_6Z?@CQ 4&VIE$/1"*-M.ZATS!J4B^_PG1H$ 
@!*BO(M%8=6)I'A%D&:YP08,-N.O7ENP_#_9DV-!^$0H 
@4V U H("$QUIT)HADXENIYR&3^4?S0U%3:IU#31,$;X 
@GZC0V^2"EJ1Q\K,@3=B$!L5Z.V[)RV;N>U@_#)*M$J$ 
@['Q^O?4"IE&TT@.M.G_(63.=KZ0WY7>ZU=9& Y.&CV4 
@3^NMGW6:0L*>[;36\P5N^$#8V57Q1L"./7,NO]<+_.4 
@?:0W>Y^_=V52ARMJAU)XI1N/+E&6:_$,:[<)9D+&_A$ 
@\:5?HY<-[4%2T((7^#N/G^*]M(3-#*:M^$+GU\;Q-(X 
@<,:J5U.>E0(R>.8._H"90HK4 VQ2&F.U+H8N=D'],.$ 
@'$ZQF)I/Z6_CRW<[C<L]Q.TU_(W?R6U3^D(N1HOO4K@ 
@M$,_9^3HM\$VYGS,4;TX@#$\M3K!$WE??3>,U(->6?8 
@"-!S%,2(&/.3D3$.VMSN^!%J0D@K.:<\ S;6-#J=7+( 
@#1LXXYD!A%-4\EBA+G\TR+<X'8[EM)TMN@PL18AY"RL 
@[YP<W,\R%"K3HN];P^RIN0W0X@\]""PV2%]Z#&XD1;, 
@;XSYU:3VD/BZ9]C<96.1[8!7LI$AE]&DCMAY=?L7;#D 
@#\)*YP [WELN+,I:8S@URZB_@@LR53)X@MU\!-,+/4\ 
@K/X/?>5)&EF4J6I NC#?:W0E79\L6<;0.Q\/VM1W2\0 
@'0VYL^(AW"*NV567/7M4FX MC#-:3(^#Y)R7S,05Z-X 
@:NWLS.]<:$<@NQ2+N[<%9,:[\#N_=3_- TH>1A%IJ/  
@V=<_Q_R2H/V'X=/8B[-LETK]K0-LD$/$/+U*=;52L[\ 
@BIZBX<IN:8UYBN)7:I[=_:$8 \7$^FD,\F@6.>6Q$8\ 
@N?+;-[]D3&]UOU+>#&F)K@$?W]Q[<F2Y$SN_3)WB]XL 
@D?J/T!LLKFXG-<LC6:*("*@;(T0+0WKB%CIK"090[#D 
@.80 9@#6$Q#,;F>]6WUQ/V9G(X<,7)7/]SC4W!DB0+X 
@+(CV<J3^]>Q:A!X";%EE% X_,)J0 OYQXKJ@ZZ^;_E8 
@"XOX<G[^!9N"9!$7A)=ZZ[VGAZ:DC=[34X1?<,=S8#< 
@61'X.Y)K?[3YFO%WS,N^O0?9_75T6]XL,>3*_JK,#W, 
@B05D]VGMIGB"4.%S<TL@FUD7CZR$I<\'OAEDD,V2;W8 
@+))NM1)>DAZ$4]&#E]O2X+68!NQ@UANK"U==EC:!3A\ 
@[$$=&B@-,FAL"#[\H9=&$UKM032EPK4;+55[L  [BS8 
@("(.<H*NFJH]^U6*H [D5Z:07#HY/V?]EH27\@^UY$( 
@^7VW? RQ_V5J"(^^..@?^;<J<ZO&\T)SQ+TR-<GSHC0 
@U^P92I*@^4&>?P<_'H<V\16;&.*#1 \K+\-QN@+8^+  
@NB\ Z4!)@HA-BG2/G3&XK90=DO"]'*ES98>[NF"R-'4 
@SP 8,KTRA3%F?GY->V" 96=1#GK)G;G#7_20'^7ZNF( 
@$U);8)%:##PO0D;CJ)ME*L))H\Y1G_[A%_10<5TY]&( 
@/DB\*,!I#%L5'F$0AK\OH_K_6"7&M%=/W4S&RF2L8>( 
@Y(2,CMQ_^JR$JFQ)2^8_0:9LA%+[1!])5\ K$-1I^&@ 
@9<,Y=@^*"^PE50B;EWQ,\CMNE#';-]N<J@0SRO!^%C  
@I*O,YDB'[Y:U;QT!0S*Q-S-#@2 N(ZT8'D'ORIXKJV  
@I4ETMN"1AM\0<'K/[J,T2TO?>WCMUZ$;>+5D0!+1L'\ 
@7D5 ZCA!]=<N@N3RR9TDY+T!X^(G'M.,L?IZ1:M1/(0 
@\G&I*=.YG7I%J#LG^+Z='@,IT7R1>\A9\HU;+@/[)5@ 
@N3=_^7#J[;_ 7Z8"RZZ)J%"K/S?1XF>&1T.0+CTFLF\ 
@XKF/"P%8K(=P4OFQT7.-+5YL3:=5@OD QM=FF";T<@T 
@T]@,RFN=#MJ'DGCIALE'([]UR;"D");2[T_]>! &9KD 
@NW&=QVJPO&CN[L&KKP6K1!15RTC\!"_M;LY^=+.:#PP 
@X,'+H9DB78WU>2&Z@WVV@%>[BCL:K0V5F%H\6H'/7CT 
@6ZXZC52B-0EC(05J+.5C2T?ZSI7./T_?4%?%E@+\4GT 
@A ED,"[2*R%R4[U6-+?L1N')==:W_&K?;5>M+[TV%88 
@]T<:,! M^U+5HT:&-^TA;#F0M4$9C>OYX;<YI3)/%R, 
@:R.?L'3>S/ Y10L*&NJJCLO]\WJL$/HHQY!DFR^"E$, 
@(0PVF%)!L7"::0WR"=DU"Q129_SI6-<!#B7[SCY_J;4 
@QZ!R<M!:*KG//KTL1Z$.MQLH7AS+;'*;-Z*4%/Y90AT 
@YC"*M_21A%=%.4=^/6_1C7C!8EB#]Q3$[I6H8=/A^;D 
@1=054TZ;)_?78X9D@4!Y)ENS.F$-*JLG)+C%#AROJLP 
@7#AC"$>#$3; +B$JI$4+E#\M@I63"W_%3@#4&CC==3( 
@'ZPQZVPU6 8;\*G"Q3^-IA.]#[U:U2C*J1*"23(YMT( 
@YX%6X\QPUU2MY47BQJ2,1NFXTQ2I&5-P..D_+97C29  
@^5<E/-/^VSDMLT[W3[4=$PLC+%UA$C,34@9&QM)0OH@ 
@.J2,O+C^7I*>$!Q?3#.^62=3H"Y_-#[M_Y4E5^YB$DX 
@,/%;;O^$@ _T?-]:"E&E=PVWX2J76YZYI Q6;%5NSH< 
@X(EP<+0-D:U83Y/V1A-N,N:\V@[@]]26C:;395\^NC< 
@^^&K[&J>'0;HS AC>)X^88PU: $.7X@XWJO%KW$S96H 
@AQ3\-7+'&XK[89CJAC.1@1(5'TS#[ 1&T:[NK^UG[#P 
@L4I=Y574_OD[ME'+NF-]^%*!<X*J#MPG?(F5 #6Y1$< 
@E!+]8461^X:%?O4W]&@E#W7GWQ2&).]7H%Y#>,XO<UD 
@3CU$OJ&\3'\FJI!B\F$]]CK:1T!G2LNYO'@)1F:%GT< 
@=H!VR03P04GVJ:3<#]\KZRZ2)O_7@W#*$[6S[<5AW"  
@YWHFFSE6/U9;G+.^AFJC&M]2+N@9\ B!SBY3T*+_X'\ 
@9L\!/YGZWBG*8^,.1<],9E.[A7=![U-H>4E@9 )@=L@ 
@'HT7VZ="#'8TN[5XPVRX"CC:ZE">=0<+<IB].6XIROD 
@?#V"E\F!:"U*(J=U8 P1,#?$4]J)O-"*%)SU9.W3V\@ 
@S]*)%;OTQ)X%%V::>ET?'R5L'3X'[".[<3WT=*FV>D( 
@YI->1#X)YM&UU[5-<&^RUA+=[BHML0\;<*%5O:CM"EH 
@V#.):B7%243UIZZ^L@U;&PY3LI^5SC+%.-.UX:M$P3$ 
@%,/:<& #_]XW>H>Z)C$(>F>%Z2VJLER_'BN=. 47_Z$ 
@#=V-K)/BRV0 0,[B. W6%?Q*0XBJK4?[==GV79.QQ,L 
@#6Y+U#VFNAG$K*!48L5&IC_0\\_+<C T1,O #IJJGTP 
@97#C#9ICS:\;.O<2'LTVHPC[58HI:])5N$LL;V,WG;D 
@**,)D[4I[^.RT%(LZ10V4?.!1%C&X;JH?D]@+SE^H4X 
@TM6Q=N;C;M%))M70P<(5(9JK_6WL0!LLJ1/!_3[].@8 
@"&SNG3ZR5@@3&V"\N_G?:\9(.]7=U%PZU\M.T'SI3C$ 
@O% 1PDT29P53O24BO'CD#E_B>EO;[UI<U":';E9H5$0 
@3J&A@/!N/^E?X244/AEK;>3ZB_@8],PN;&7<-_I(:V\ 
@E-VUQ"^%]LQEH\D$&)8N19:M<Q5@)=2C._IQZ4+/W2$ 
@P2QPVDW6I$%\:4$[\\RTE(.\1\BPCW^^,"'A[RA!N24 
@IE#W$>F&05KOO1],,WA*Y!1FA!HL(@\CQ&>NBO8I&\4 
@/(:SCQ<G11O=+O(BZ>QZ'R'HCLTZ4@]3#1,'I(;[5XH 
@N:J>+W*KAQ:H%1Z^]>OD'<J-%HUL0Y 7JZ.3#MP %7H 
@'/,?):[VF^]Y78>(1<TN9$$&]ZKQ22JNS*J7%'.[*:@ 
@O4#PXI";%>SJ-'MQ-S#\\.<14O+D8#\B.ZJ;Y-\QIY, 
@QO(+8)CLTW>Y1C)\8A3;4/$=>GI^4XS<7X>O]%HV /< 
@@$ 8<V2]P'U#';0>NEEPUNNIR_&3U\U[X\IW-*';:\4 
@(_Q<DF A#1I^"C\$#%Q<:XS@.)W#W_L)'M[M*W6S8A4 
@(K+7+0IK#9KR";-7@R)];5 2,P=:6(H?"=_\<WL$C0L 
@\I:>-[3E@O_6/R#/0MK76TR@D*0I4'# ZJ<^:H0*GZ( 
@J#**5ZUUT>SWBM\F$M@-'Y#D=X;M8V1O2<__F_=:2&\ 
@C_1V!Z;9^^2+.QN*?N8K([L$.E1.[,]FMEX#7?;#+)  
@C5&R3*=ZUM*<CR%LI+M%^D%A2&&]CBSR \XE,/]Z&<( 
@;"D$1\.YQ+[]"[.N'[OE04!&J%O9<Q=V\OY)(Z.H&^L 
@E:.4;U\03#2/F=!5%:CKHR:KC7+LO\)>Y>W "X2QNZ0 
@62/WSW$&-K1AG;J?9FRR5S)A.HMB)*3+V]I;[D8]7R, 
@TZ%"K](. QG\I@[\#/)10 S1U8P\UF18>;I,C >)J*4 
@!.2Z9C?"2!O9JSEF ?_H.!U+Z@3(SV4AE5'6C,E4)*D 
@FI?^4R40Q2)20<X+OX8"Y6FA @X-\YGW\>W!ZH('MZP 
@F"QWP(+GBV%G&6QA8V=-3>HOV.#8C;D0!4U+^?ZX"50 
@Z27X\?=O6^>>"X&\I(<]E;^JN.-FAZ2M,OK]+RZ=, , 
@^B<!?'TND3OLRWG/"8G31ADQ>#A%6>P]=:!?(HQ=#_T 
@6H>++VVO4(O9RI/?T;, "$[V?\>BKT/D$+31&QZJAS( 
@[*C*:>575RW"A'1&_%M5"<L_0>I#"CG6W&=UD[[>G[4 
@4IAP&T:5 >]J.(%Y.AYGPKF&F]($N ,6 >RH02GW3W< 
@KL<81>[A9(O&]OA?<EO&8V,W*>(ZWUR]*^Z5S,^K\.T 
@6#6V;,$)D1Y\$Q0]5=WK&)B%C'HO./I7DLB7F=8"63< 
@#M68Z99@*R-X,4M6!C>A6/CP,MQZZ<52$[# ,;#_BI@ 
@\BG$-Y7:O0?FV0#5Y _SX0PWJWU?;+PBT?!SDE7<TU4 
@C1U"48 "92GM>0U !)M*_U0&=R1:%PS>IW]C]XULTQ0 
@^HW(553_1S6U_N]X&5[PR6;3B2;P,[MN)F8P5@<Q/^$ 
@B@ZW8"<7<F7/T,!\N@?_-=3 0+&WU+P&L]GVWM"/(<@ 
@&;])KV=:W)D)OP?!!1L927B!Q 'L'T$A_-](5="\IBP 
@^1]:CQ.W [Y^=P^#PECUYRNQ!?;0CJ:@MR?P=E3*V,H 
@8LQ6 .MMIB#F;1;W*1G.IBW%?DT#'+0#.=2N0.T\C", 
@1Y),<PPNS*ZL-,=.F>/*]3"+GSH78+%D.YKYS76&V&D 
@0F,!.375 '4NE+?!W!LP7&VA?A4!A^8?V]A\ZI(!27\ 
@3W@K[X3!T;-44M3>>J\P[@N^YLCZ*T*/Z1.V3+ZYW<( 
@H,)-@$A'Y$R::4?43VVXV(:3I!^#7@\(:KGEQDP.D[X 
@_S_Z/(]T^JN *:Z\_TTJ[=7U<RCSD6 W',*^Q^*!Q*\ 
@Q$(#-HC6]*E=0V;!-R!!QK4*[E+M5*WS"R/ 3RJD -, 
@4NWG&,W=7R=L??MR.=26CPKHR0O)5_H.2UFP%P4/C)T 
@O!<D:?H62EJ81VXOM48.,RWKH?50;5'TY)*G<*@F)<8 
@<%<.UG*AE9^;KL;T+<R5RO-@@#R0E6C4:$09R6RVU,P 
@7T[RH0#'(+UN^YY%&YS"J;E\PO 8:;'6OO< 16?+=D  
@8HTWI.&QX<E+5%1S UE"J[L<-T3N2BP$?;8W-HJ>2<L 
@H-_=-8@U;+E? R<H\GZ697GY(1XVV=!N>SWR/K^QBE$ 
@C$SE982+7_[47ZAAI^F^#&0KP:[$>H?-ZG518&>423< 
@0L!>9L&\N5.:*'DEM%];+PD\FT6/'4H8^[+7]3]+\T4 
@$I]CIRI5"_I,?!@_YYJL['084<0VW L';=D32_+Y<0$ 
@)G-U*D;E9WG#?\B7>4GF 9!:$!*0\ZON,NPN8"H$K5T 
@D$H="A:0)CY@"H%P1.PI(5\_\8"^4.=01V&F8FE6)0L 
@2>N-Z*6]FJ-Q&"@5H&],4BB7XLW?'W8^O-"4+41/,TH 
@8!N$%Z">:$<5IIG/H;RT73B7#TD@ER/LR92F=Z)ZI.X 
@CF].68"AU1EVR-C\\3ZOCQ%W2F8SY- SE\9/7R]26G, 
@\F3/*)N;H_#Z=+*1\Y=!?N1TIR459F56T3W@&+Y!U=0 
@M GKJ\9]-A#2'MV>2J&V56TNYAJI7T+&)N\#X$Y98*0 
@KXKRB.I.=18Q%573A98PE2#;;/IP#-,2>$SEO(JLJZ@ 
@I6Z?R1MT[&R84IW;&(JAKQD59&IO+WKM+JA8MXTS6/8 
@J>D&D>0SF;''I8GO2%9FCM<H*P]9>-%8<M?^]E226DT 
@M)8H>NV*Y+)$1S!-M)K9KMWU^H3NCTEP*)ZIE+Z9!<4 
@LT$&_<,(ED?+S,A#Z4"Q>X:Y]KS@OW4;/228]E"?DR0 
@2,,;*@M_TBZ&1.%/;B[^G: )^CEJ(&]@4S?+Z78>O'T 
@RH5LLR&=_6G<YP/X!.H5BH6FI MA3_,]?]'[R1S_,R8 
@Z$%Q@ZJ9= [JQ%$$'-A#V2XTIZ0P6A(-F29K*#H;07$ 
@ER6[?^ORWA,X"QES@L<OHT7*=6+LT]C0X KAA@]S\YH 
@0]I 3*D$_AY; '&,NN<EL]PI/-\1"@\=U,HC(;-I-GT 
@I"TFO86E:*U0$^)%B>*9S4SQ]"=:=EYEXVF&K]=JJ H 
@[\@#;QRD4*AT8D/WQFZ3(MW*.5T5%A?C). RU_X+C,L 
@8W<@'"'-==7D6 ]B_#UD!3YL+B(T,G@8^_;T9XN$8@\ 
@LX+34HUS)\=B^+L-<D2!$S-_ )X"..L:X<@[Q*[6$+, 
@-;X5MN/1[<DS:M!EZV'4?3(M)UWKY&/7F<-G1(JIC@D 
@1S. QIS%/\H.&G;N,M'Q6$]SQR/%D1,%+10>HBPI>0H 
@HQ04]B750P&+KAP-KL!\(6NL?2R&%LX @F.=LC ^^W@ 
@R+J^F$ 'HFZK?H0/3AV4QFT&Q=U!]>V:'8--PY9Y-?P 
@B@$(68-ZGG6#MC)N0EI)(0VYQ"91VG:<*'P>9-OWN*@ 
@32*1$307>WB&G^]ZG,)-4T'V7RWK^<UQ-FKP!L,P0?0 
@5/XI<6@LRU\6X'WM?$(N!DO"FX0K*Q$FJBK.,P(FLLX 
@R8]AVDYYE@7VB=>6)?@(%435_C<PQ);3W<O%&:5R$XP 
@\)K^_J+JJ['^1AMZFG*XYI/F(,2R]56+!%]WGY/1VA\ 
@_6%?*J=:A\^7=EA5:LX0O\\I7I=:6^GL;1!"R$M.7Q, 
@V:I472 .LB8-R=.!Q8&;=)<) W+21C)$:+7VB,/'UGD 
@Z7,]?7FF8CP0K8GY:1FWYFK%K9*4:0.E\$U<[%*A&[( 
@0.BOKVNPBV5((JRT9K.Y*Z%PM^3];%4N<$WE6H_;>N8 
@O_C%Q/I;P[U>^ .1."*=-.55$?_6M,.S K$;B/_^; 8 
@C^O1T["9!)9?/;&!!5%$SFKAYE3D/H4MS6?-.$;]S00 
@\J8P%K,ITCX]+08<I_L25XB,]<7@X2-:P@6.VE/I7UX 
@K11EZ=00':XZV%I)FD*\!C^8Y/62NA[%)&$/YI-8W\\ 
@J##LK#J:O5.L&N,=!E,:2Q.2!<BB=40&43EE'/,1IEL 
@B;K;';R<_2F29<:W82\FL3D+AE IUZD?GUN&QL-3V^D 
@_N;$D+N+LI6*@VFWX$R6/8 _D+&H"]R9J^=G(^CHU]T 
@_48OU&-E_'#;'92+-LHZ6=T<M%AK$F>S%GSN>KDJ=L@ 
@><MOEQ*15$>;03T$_^BADL6P2T)_UQ1A$MK"NYJ<V2< 
@"Q(APEY'/_T7J,+:B,ND?U5U"P#$YP)OW<9Y,;70: < 
@% # @M/XIM*/!?>I:W)U(N+05#Y4FK+7U/* BL6J?7H 
@G%8.VX=2'R1Q%4.H]]'9'L.XJ?3.5,-J."%LONF#$<0 
@6]V;RANRR_'*U'%E<>Q[ /7K9KZ+M F9:)!!E:=Y!P0 
@>FC< 2*F>O1F/:9D!M%=7ZD6MWZO,Q.]^.(Q1"@7#-  
@0<.'GKT$3!OHE+3/!_02S!]O_$(QGY6^ MR6! 9%C&, 
@A;[.HO0L11/!7=]Y\OE0.B66$*":#YE<%*E\*_ME? D 
@6KD$#"[QK_&+P'31Y@N/:I6MB?$8/B_Z2!PPNM":D(8 
@NO.XW3I!T6_=SA#5"ZW 'UR/E6P7SJ_O"Y,MM20F0!< 
@J5B!V=NG$8CL)&J[5RPQW?( 4]/8VJ-/PG,J?(KX-BD 
@W(R:RQ/TGQ F6=<P^SHSQ<" &<S:C':.;S7_9'.CG6@ 
@\LHQJSA%PSXLJN&O6%<+7_H=F>_-T&+2[8??N!Z+6V4 
@RW!^]R:G*.MQ4=LK #!)=!:G7'%/AP4@<^.<C;16)GH 
@2X8(W7&E)!R+T++B8SZ3,\8H B";H34]R4[(_[>G"<T 
@-:UK>%IQ2,@(7Y*C"@'![L8986F0YB$B00!FM'U_Z"  
@I%I10NAI@'LRG!,PB!!5F&CF,](62O2Y#[0>N43$IUX 
@ JY)735"P5WOT=#6&?U'?3>SWMMZYC<5O9!5\YWOP!  
@8G#:9GE3R8QTHA84^+;,CDWT#Y??CW,J%'W !+@= BT 
@</ -DC>/J3H6 ?>U$";SA2YL6J:-SB/M&$/#( P9-D  
@4P>;>/O1DY]F$KR3Y3:1B38/=Z?3O&;(+(,M<*S'(%$ 
@(,#,="9Q"P&J:BAW%Z1',7F+!,D\.X/ 8IP@:0^Z(DP 
@#TP/ZTM* 'B'D+_1L\ < D5ZW&@\ZUPM;6L>O,ZU2[D 
@#!Z"L'55N^) ;T(S &BKI^W_P"*0/?CE#8@!G6 092L 
@1581S#.Z8%K!XH >BZ0&?ANJ-[C!V'LU RO[+TTMG+( 
@,&LLOY?9TQ;+>&J"8IYP]+=VV8HESF'$9^9W=3R7<J@ 
@JP]4*(=<'/TD+MS$3^-)!@S7*NEY!JJ7"\YQLJ$I^"D 
@C(4R5VR E]2-6*RW@!Y* <#FTZF%AXG2&&1'X$DG)L  
@\M _87G3H G8Y QJ"D]<K%(^B\5_%['Y55T6$F[5Y4D 
@$+O%4(.^-GJ3';*/(MO[EJCW>6$ R#"Y-H5@:HY2NO, 
@[D<S'X&%U I_![))$'D*$BL6Z(ILHU&.S(,9RCH+K24 
@7IJT^&_#COF[-R@N(7. WQB78IPPB3/VXJY_+S*3+:, 
@TX:78R7^='</RU4@0+3IB6"KK9/VPLFVA5HT[<)V9MT 
@<"COI=/'\DHP2%4DIX=QY,K>_LNW8( S52D)($ZQB@L 
@E ,KA[.A[1MQ[D)+S@^A?&2O![0%$OCRPS8Z R:?B_X 
@7U^:=*1S_IGP0R"YMZGL(6[S%%/N<MEPMK=,U)Z2>2\ 
@ $.M1]2ESHLD6543;!:W ^)X"&B0YE+H.\,0->CRL=, 
@2+M1QO Z4,[6S^GYG+)XCN.)WM "$WIX(ODF&JJC:C@ 
@G]DC;J"&>Q?WRO&7J=L,\L@6PF?/T9PT=8T#W4<2PD0 
@_ R]-L)^31B1%'DO6WLP&#A*67I=*#)B:YUL[>VP4"P 
@(H+=%]7 +F 6S#"5(P\8&5%J"_4]ZB0 </;M= >5;Q( 
@=E\!RXBVZ*'(0#<+\9#H<>8]"W1BZ,*9XK\53!"^XOP 
@(K<K>D92;U)1>C6D,2,#)MC,&G<AE)PP^Y*PRKE'\6T 
@0B]$:TFJ") A*^9-0]0#"#E//M_?@NR \C%2DS:Y,6@ 
@@5'+8_JGXA^O^>P<N8KA_5FPM/1AAJ&1L=W9^K;UCF( 
@V86F 413,;)1<RVNE"A;;F!4)2P$A*/7H'WP/(VY>^T 
@'.$*-JBI:&V.&!#-D1UV/@Y3N6Z&BV3XJ4AQVIQ]S"< 
@:]:ISFNL0L/%Y=U"O[)$?^_1]\[^Y%7@+3:M:@'LT0P 
@0YZVU^(YHF9/(8N8J,ETZW_61>VP]H4#H!JD''<TC;P 
@:'5$5B_K,WK7RA0&W%BMGF+'8%W$K+XLNOL^\,\<8%D 
@DC?8]_5#K>5UR"8'RLF/%VC\!?*,]!R*7Y6[TBE0U4H 
@;QG=\,#Z5R"$AFD:;ESW>J6]]ZYK86U!X; %U<^Y#,X 
@9K&W)''?C-PM%_)3BK??'((7];4U1<$5#X*,XO&SS;H 
@!'42U,R5K!B-T4SL^PJSL31_)*[H;*[>"4O8C_H,7%4 
@!/+*Q%#*-BM2#QM\\;QH2O'&8+,U 2NA1$_BK7;)^<0 
@#W (I,]0[,:]31 &: \U=H;VYI\,S_K30&3$_72Z-ZT 
@X;CM\EX@=B4Q",XGYTV0>FK3"4T>YF0P&9+@F>^U@&< 
@VK,#9=/5:9&9"?VI3 MEUGVI3E9(&+N<>K,ND61*;?, 
@%S;9D@^6/B7'BU[A,V;]L#[I!,BO:FX_ZB*O%7'(A*X 
@,D4A;OQ:E.O-1.2ON9I7+DB#>'ARR7O'QDIJD6U!.3T 
@Q[%9,$%.Z;$V5/]!]-:6B%F6FI-)L7S)WY\AQ:\1.VP 
@FI%VF(K3R9))JH26IO.0%8,8?6$'=/P[ +H<O#^VPRL 
@>86&?UATX<PL;1ML]K(<W7QE=+=IARZ$2 &NVA@T&>< 
@C*5_VO**O>?O3%>&?TFZ &2U,/\='6#(M^31M8627@@ 
@F45,+YM$89@-TL>=XT_;A_]/3]Z=  \D#9?N5ZX$N%( 
@M=Z^%T/PZ\"NOIY]]%; Y2(KL3R@)2W@:'Z_3Q@:.]X 
@^OMZ$L1.)];1=/,Z.G9,DKF!6:R'+Q15)QD?!7RD: T 
@[\L@5'>8727F2/%.*SSXH,OD(EXXH+=PYMREG3H)]+( 
@&EU7(-G[23+=!4 6/A<BE, BUAGKGZP5C$+;76Q J,T 
@3@37/J3>A"L\8I' BU$=.4#-33"OCUA)Y&YLU%L"/(4 
@->"+?DU#5'S6Q^N#Z7<6)\)NP)O/)A+H4<F[MF62U/$ 
@%-TYA0><5 &6TV.V>YE,UZ#6FA^O1RFQEL%*)+(2XT( 
@O6-K>P1=ZOJ0QNK%(O#^(F2,*TVC7Q!A:E4U;;C\+R0 
@/V8";5I9\'-K#8 F-O<K:FX8>2YHB^A1WM&D88TD"?@ 
@>@M\L;H0_%6:](@8 $H<JBX FC+PV*XW0*^*2+13+HD 
@K">@KFG*:?&&9>T*8)_Z+J6U;6N;6?JP157RA$5O]<L 
@CWPBR;SE^<BGG0/X IV59GP:.[6$N3\[[ &"(CHM_T8 
@)3OQ,U4R#T<.,L?_@G]W% "L92,%:6X6]3.9J[=J7+T 
@,KMKQU[\RE!$"I+\+IM!V/5/W !3MQ]$R[<5[Z,L5)T 
@54.CM4/SA0%\_+\=N.Z/[.,%P]'G4!-F 29;%!^?@8( 
@ *:!C[K?9'AUH"IDIP%_/IG_1K:)8]GK95,ZDD:KXTL 
@\NB\Y'<1!:?#_LTX]#VG395#Z)-5MJ3%S--"F[XK#7D 
@OPA7%6D[;*BU/C\S23X"<;V!S"%8APV(1NVR<N6G+38 
@VA0Y08P!Z-W!#VAP-+MCG@'N,2#>F:><21,>])R%T"( 
@5K% Z]5S8&#504"1%3KS]M@6B4]-5DXHL!Z>*8R H , 
@TT!)^<NK3;.T_P $YC_<\P_ZD+O59&1$N&S4"*/]&-L 
@06"M*BQ0[P":;!T?FYYU3I3H4F]SOZN*NYH6TG^G,)  
@O4.F4EH6"5=90=Y.N!]@R- ):;[Z%S^'7#G"P"KCL'H 
@V9F>K/:(5 J2JP]E58IW/O+?$DQAAT<.FJ]W7*>]80L 
@^(JA8$X@VYVU[FCP27RMU,\?4<$^$02>X!)KB#L+%L$ 
@ 8T1X#XT0^2-K M#9C3\6S%Q1ET0Q10IQG1!3E$FY4L 
@II*LGXO?G7=)Z7"9Q8*Z="EP5T&RTG3ZSR8G)0KJ_-@ 
@:PDW )8=D4Q'CH6:6V%1*=$@QZG^)$ N]A$6@0S ?S\ 
@)?O;GS.RJ':JN24QT3I7.BH,:0L5M$[,!2&:!_XDB#  
@B8Z!3N9H/J"K\_$L6?.9>N4N1!4P_.%FE1*4-- #A]\ 
@5)WNU %;#0)T1\LUC\WV 2R0=/X7LDMPB_,#"0<V4<H 
@($4$34WUH3,;_W\LP=.D>5WA2A\\^3;8]CO;\FD O20 
@Q] _D1#-4+(5V>O(2L LV$6G6XB]328XUYX*M(Z;!#4 
@N<![X:5[V"^6HP=2 .)1J[H*9E"MP[<7124PZQQ99?$ 
@&D"Y2G:WT?_!.@=WMUV89E592OK%25-?3D4 Z6Y")X0 
@Q.5KN99+ @_H _@-NN\."W%3PA__$8H$!7, \@!L&!$ 
@@"(R22)N59VZ%NSG%D3SQ"'-Y[*C(KHZMULC^7*ML94 
@?1=U8QV!.I92#U[ -=;ZW-:,(&BE&)%"L&A\WM==BP( 
@63_@R<$L*E_<A4 %[DN.^(XC)!_(!0 FU!9U[BZ<F%X 
@-0".S6&VZ\".]14PP]>X3-?^7M#"G& R,_^43HFH] $ 
@N[ARKA9',?:THU$8[=(,+%;R\5I%P2O),6=Q<ILVD#X 
@P+\^\%!<U+">,'RY;>=<AT>@,9@EVZ+H9)OBU<L2(5T 
@U]LU.Z[0';+U^1%>8,*C\Z%M1C:F6''\VL'JQN9_+3@ 
@H&S93U$1WD^.W2>(UO(X!$^[+PB 8\RH+"[K.-9L:TX 
@(Q@ $'"%Q9I9*.^ B)5LVF=,9@ST2.0G$P"L6C 8!VD 
@+>V\"A'ECL(@(Q131!\XJZ9R>[9A^F-I^N;7J:0*2]T 
@[<1GU $[F9+_FY+G"K,-$=A=Q%DS;;H:)7'?<G7>-OX 
@I?;1=>4D)^Z0;-Q+N:M, (=X1>YC\S$8F0#"M3.#\\  
@<WT862#8C8MJAST2^8JF9C:TE&MNSQXE,]X&PVMKGSL 
@3@RSS6'RU D@)"AH%^01*%GBFQE@4H_F!;*2V3VS8'D 
@!]>9I%6+L9$=)TV(-0[(^QO,BLI>&>J8,^XU)CAA!N4 
@4)LOT^[&+&<2M/Q:\1E4=BO2H"12^)Y$MZU6R+U<W6( 
@4UC9U<[(#JCT+ X*>1JQU6V2460HO\4*,\FK'[-(I@P 
@92S2RCYSB[W2! =H PV./@T]ZL6*:R0J])'4?BF:D8H 
@I(4M6OJ]@@?0K/7:"\V:7H'U;KE.Z78$)Y#INR)P(,8 
@#JJ+"&)O!S[+4!83,A\C;K0%C&2V<A)HOQ>>4BP3O'8 
@; :&%[:7B,&N":N$UTVM$3.D^&^ER!!-2J,V46#'IX4 
@R>5?)MZJ('+0B2LX@FHMVKI'^@!IIE*2T1$[JA1<YOX 
@(5&MMRE+2,046!0O=Z:#I:9Q'"52-*8"RCQ4Y3\\#B$ 
@#JUO!FO;MN8AEL] *<JP=%Y]#T!I7$T]->*@5W"U(\< 
@J_%7J%I/Q30M2IB]#3=7UN&&">#J,RB6$?U;^\265C  
@XQL5109J1U&? <J$A-G<.,T_!VX0 L$-QH<6J9QET>( 
@NW=)F%6<$:;MT&G#\Z3%VEJZ7SHX>H'!ZDAS-AGM[/T 
@!W='>+=46BCUXLLP[6@Y??KSW"@+@=_G>:-2S ?4;FL 
@>&WKH%.MQ(A)/(K#DYNV#+ 4&5L?[>P<KHHT2 ?,PCX 
@412;U(P/HXA2\W)A)!&0E0RA=Z8<,O/V=JZ^M6JKH2P 
@L)J.W$0"5-I6,'<W9^QEF; )E4V'Q&X=#/SZE+7AUA$ 
@1%,OYWV$LVQ]9$0(-G:TMX!<E$D&^S,O"_?,ZX3"Q*$ 
@=<!MZ!(IMT=IJ\7@G%ROZCC8)A+( R$I700;KK) ?1\ 
@Z+J5J[!E/HB([7AXX@'%D+^</'UG\,UO-;-WANOD_), 
@V74'N&Q,?>]@)9-"R!(VQB%%.Y/"Q[K.M /QH@F6U5( 
@8\6TZ)#M%JL7-IZVAHH6G%'!XB3A@AZ!)YO9$+%$[S, 
@?$+_/1'E9KC_ V@Q[_LP,O?@!ND&LL,N \MV.:'WDX4 
@&%$'[S6D-+I0\C468.(6>$Z:8D1\,P4N$4RT@JW.T0D 
@S/ICY?2HT:=//Y5> ZQ?$S%=P;+7$=I;Q!VWFM0,2MX 
@ABUU>H(H=*?P!35HP/FK#KB9#)@>T_D?JR!4>OKT)9X 
@U"Y5Z>=[3"A!YA5+(#+:P^<U*3+8RN]"1U B^6:HAD4 
@F"766NC[85SMU'/5)EX=6 NEZ5#\+4$+ R@-8KH;(_H 
@#K)&5K*5._IS^&[G3I!2ENXMP(U]Z=B3,#57 <0)G2, 
@A8]TR+.(+C,T;(E]-?,,SMUP'^-V$0_=EV-8:1R?L6L 
@=+O.HQL5,>IC],""&X#I]ASJM[X]M@"CAH0USP4FC%8 
@FVIM[&/RQ?1[4=$1-VMHT)[-TW1GBOZADU$ %"!-BJ( 
@%1O27I+56L\QJDIV\9'6OPY<O.D (%'8KJA ($"U;-( 
@LMB'>] B:V:Z09J+40$D*(1?/^9*(BFR"_SLTE&&/NL 
@UJ*Y\"KCG04%^*97]1K4ZUCXH*\3K@]:R206-7[2Q^$ 
@H=EO]$DPD,^_)$6Y%6F1K[C&01WSCV9,\*MZ82_A:3, 
@LWB6$W[DQ6AZ;3BN'M\_<,!3KVM.#@]P2C!RJCL\&9L 
@I'<)"%7R!:FP"7]::- &%$?/&2CU-7)C34^&N4K<K3L 
@)%^=QUS&DFUHS#"74;>OGD=-3*#/A>CG](WDC>#!N_0 
@+\,GHPX$]"6_7$.NU($R=,K_)HRXLBL$?:MN&C1/,90 
@SNC]O_/*,ZH[08/#X1*(+&D&;V< %Z*GB%DD.<7-=DT 
@,"%[%AT=$PXF075N=]T1T@B:K#2R*>D0>^/5%SMX_.\ 
@H1HRW:U%9$Q6UTUL0SM%-"+GF8%"-S>03$G.-Q E:N\ 
@J^5CV,0V7W7AN];5^A26M&Y_G$XI&D\:ESV,2Z<600X 
@C6)_0BK;Z%$&O[T"UA9('TLW(VM S>!41^L(9GENX9H 
@B4SCPD\ *H3$F/[LAK/PMJ++=;MCW-GH7N1&WX'Q,54 
@RGLNE8!06#\*BEOLQ"2)EQQ6IUY=,T(A^?Q8S46^S$T 
@W8QKZ!OT8#"V':0!1'O+^K5DSEFB=Y*N6D"J#C#2SHD 
@[T< ,4G[N=]%B>_)45M!SHQLM,Z6;D%--#"5*IYXZNT 
@@.^TVQEX:&/ $.Y?/9_EO_%SEP$W1=>_Z?7("*Q B30 
@@%+)MH6SF/I;#@K!Z!)@%KL;I,I.,3*8!3 G'V<J% H 
@09;0R4%S'EA2**ZJ:7'T0I;XIFJ/-#:E#EAV;)2W55< 
@'483*M>ZMC@QP.-X\[\*!M9,O$?KUD4#@3%U8ZXJ9H< 
@%>,Q/"<!Y^5!5SIRXIA:\WIW<9=F1 9=]^D#UUGWQ#H 
@]%,F\]3O)K;CCUA%70LF;\'&3SP,ZXJ"6/4UP'Q6#I, 
@MU+0&*GE54TYC<1-PS4V$7^BW&W9:69R"Y5\,8M=)@, 
@&V+M?]+ ]89!878TCGN>4VBJ/!EQ7$?0TA1D<%\*O%0 
@ZCT*^<_3.I+T2(NL6PDB>.C/C(KQ(QH!=P0R[=](-1H 
@)0L0OIX.J8+?Y>E)F\+G7-03;1=VXVFPW@ JVC/1]4< 
@(/B^?\GJL98YLL_^!AJX7TYXHR3)3.F';SUM>IZ$"ML 
@'<HX,3V-*ZG0%CT#0+7?>%<CLV_9JK7JW%)O7!M7(3P 
@T8&-@H&5P8KD#&PD^XIY.IKB8.M9KI%4%U=ZKR[[AA  
@#8ZLF3)^@X<HG0CD.V%>%XZ5QKGEU7%_!&<!:A0*N+4 
@#I8Y40G"=@ 9P^(5)LF(77V#:QC0<;4%!X>N-2$0X@D 
@@CXXK+ODA-(Q%@Z_(6B?*.[SQ1RM1<<'QV02'#'1Z), 
@8]GLQ<2EZEI7;N4+)L@+KT*W7#&J^4TNS0F=X5C0AFP 
@XG6^@P:S5_80"!)\9A,]#&FO:W7.VKTXR*OD$7A/4S0 
@OCQQWW0I??IPA-*IG5G51X+JWF7,2%=0R4>!L2<Z\B< 
@4C=;LFT^V5AT6UH5E:&U'GK\W*)))"E182BE?*'CZ<4 
@][>.:D510]U^@4BH4MAE=$AF!?@,T^#Z9VG?F*<U[Q0 
@5M8!;KA\HNJR>U?3 :NTF?WA,OR/@#X$N$"JQ=Q\#^L 
@J9'BP[0MD\L]3MDS=]Q)[H42<2*,Z"UIQ_Y\J"(**=, 
@-F'5R-M2$"T_U0X#4JD'.W,CF%(_!S=2LO5TARF@]PP 
@XE.8,C4;$[WP5$/X/B^?T<(OHTZ&3_Q49"OON$6@W+@ 
@$^^C*1^8&@!2#8F(H:NQJ_UU<2$(\_V()RU3- #3TDL 
@-O<[?DBE[/2R@=8K6 VY[0+$0LE:PAJW^VL</C.\6!T 
@#/R"%R2+1$J'580Z>08;S'M$AM>#OMR.)59[.C:SX5X 
@]*Y]'3%_W301LQ-S6^E"2+C4AC%B#M)L" &RTIDW_[4 
@KR3;Y5L54,SY<.;H5;I,?M!U^H!FPYU0[.1:")4*"S( 
@DKY>/#\ASJPU;"IZ2?5)ZU<"ZLLYFG6-R?D'@8(/([\ 
@'Z$<22 "D2KNL"_5!-+[9GS6X'GKMZ_%PY:9A*;&;E  
@')GLW<"/(9?P:7-X>EW'/.%YRXYQIZ<5%@6-O!UJM70 
@1B<1,9CZ,<U!50$KT%G?/W+#C+HWPHXHC/F8F:GWX%H 
@A2"&'C1K]QQVU0 "\4N)VCMK8]IG0C7V/CP.Y4%>=P\ 
@P>BY+-J<Y-'TO.G@#\HHQA)*^ BB?*G* B+2LP=BN*L 
@E2$&2FXDS !T]AS:82VY:,V=^N7?@.9=G%736U3"XR$ 
@GTU-#FEC:^K]5E#.":Q/ZI%2J GD2[C":W88,:/1JMH 
@/+/FTQ7DZ74R>^7FP=@E$7$M:_!">.=7XOHU^+YY&^@ 
@3A&I:"E-F^OM=M0"F>!UZ=X.(+MELSHM'P=.H%7V^<H 
@"=JZ//W(^4ETHYHQ5LT%W:]L0<C48U;SV$E)A.*/RP< 
@NS5DP53:]L*6J%?!5RN;;;R#YT63.0Z*WFP>+-ZN5-  
@!-!!)&I%'='IC>T6B>(ACCXDM9)3""RRC3@<P36%JTT 
@A!VWLC>-YA'N)[#/#PUR8;ZXGQZ>#A8#Q8D:EB0Y:A0 
@(<==?V6VHW );35W3/U--M/L2+&Q5FQL_'.-0?7LKHH 
@RR' 8<IEM% Y''Y^QHS_;OA^:X*/*3%98_"L^EZ\J9H 
@(#S^A2#7J4%YC\CCW V>AG)%ZNP-X'3>TEY";(#8R38 
@K&+']CA%AO=B=#8_'<L<""01/W)5'N<ER+X-M72Z,;@ 
@'5_6/6T;RT&F5;PB-_O[N9)Q;<^<?ZV2-=TONQOVNR4 
@WE<-?YB?Q[]B9Y$++LS0''7^MGZ(Y!1E&6+LZ4T('9@ 
@N,55Y0 _9H9D'!V)Q"R<==3O'17"0>O;=I*' <19!1P 
@KRUY8^61+^8/%J5_6K.:[;%8TI\OQ5R%^=?T:5OC)*D 
@-Y'0/GT4@.V(1C;WY_TGRQ6"YL./X@4(9"%[&F,)0I\ 
@M@LX<ZL&2+TULMB:=QW'(*M#$T0B[A'W?WD.BBUT$Z< 
@+P<+3[]F?63G"M4HJ7MNO&!TZ.D;]+5;,I6:BIZT5RP 
@/L=HVF\-@F&.%,SH]@^(VMW);&\.S-2Z%"A+2%>7Q9  
@,E#ZUD5377_\*<F'=T>&.)4S9@^W<O=T])Y#%>A10EL 
@CZ\]([GP?L!N)-8W>#=L'(,*(#!Z+-+E:[0UG]8T(\\ 
@ANF\L1P$">K#]=1]AJW-/'^E@J908 ./&X$C23(H'2$ 
@@%Z:XJ<SF#0,NSD:W$S5TJJYXK@K.L:V*PO[&X E&6X 
@JM&7=X4*N ?)_12(V?M?G\6=LF[YI?[_[<FTZ<>9,X8 
@[*6J2\OY6](@QZ:J8GD3KG**)>:,Q+B#14Z=\8:^(1  
@]XIU9KS_&JO4>O$/[<G4::P\3\EI7@1M,B7.K=$T2#X 
@%&Z?\JFYVW7._0/-EE?,:4Y!,7)CD\R"BE.^!F$YS!0 
@M7WO_ &G( R1<+S#@ZF<6UG(;A^8D@DIH4U:+OLPNU8 
@*4W$*#  ]V@]=5/+H1+"!P#%_>L[)]'L%[9;!4)BT44 
@K]>)H)H3R"V!UYZ>6)I+IOELU"IYGHEZER_HWN/EV_P 
@4Z2OCJZ>5A5:<XX<65G,+)T:(5^>B$)T-GO#BC!S2EL 
@E[_6=R<$]&VOD/R3D-?0H=OA:;C]A5_R0L1TH>Z"70H 
@4B7B" 'D.3C#V\T_9:KR#SK#&0_1SD0;51[Y')[1]0P 
@FYG::Q9!(PH]4P=((V6HFT']KZ+[;15 '_?\8_S$;<X 
@-V*3-JDN'>.723*7@^J,A\%>^S&6(MG,[OOO[J*$'08 
@6+<RE.)0!7REQNRLJOIX"Y$9PUP_K+ENK_Y\+I:G1&\ 
@/Y0#<7XKJ<P26ST?_AA""O?-QG.[2AU@8D"/14_6Z.@ 
@EI7AQT*S1$,O1K83$(/1T-*,W+1F\%;Z'L7=/P/"<=0 
@PMJ4[0V\+=^JO+JF$.]O'%MK ]: ^0J)8?)1 CL"J08 
@5'QF@OHS'*T4"0H]6G%*&N$CO$1ND".BIE?R3<\#X0P 
@A*59O)7=R[S%3:J95^.*ZK<B *^<V&<Y]PV?\VRM028 
@7F)PB5P<<U,"STK*N3<KE;1%+.7"_.E[VQ7\ZB&,!T\ 
@(=AT?)M9 /9DI)<:<W,!7+6NO"3^V 7?J0LO&E*+9IP 
@M>M@'H?VAW$]H? MY%9V<E&(2GPO]7S+[H&%^6(@ G, 
@V?F.V?#D[S$@;2M,LA.16PRN>4$;#(0[,: ;T0Q2!SX 
@V$2;V 3MF_FCH7URS:?F&R@A?5:^D[R56W,-<FM'WW0 
@?PA5#[H6E))8DGR:Y7PT3V6[Q$D%+Y;_H7]/.(MH"AD 
@ENK_=QMK:=_HT*[*;)$E8YB4J([E0#9P,CG9"/.,/@@ 
@5Q@WY<\.^@ YA4\XTEEV8N8ZRA), )-H@1\_&>R"/%D 
@^L[&P%OCDQ/AA&.EV.FORP4_[K2F*3^1[MTU7"]&: $ 
@VK/T[%EFZ5Y4;[P2_ABU\7[!KC#Q"9/D<>AI.\TMVW, 
@J F<Q1@?2Y>DH6B[2^>FIH*/*@"QBU4!P36R!HW4F8  
@M D\/X(1[Z]Q^!ZEW8J)CG)2)!9ME"&F.$4(BBC\SW@ 
@')L@[V(IG6.8R*C\<F6F0\BRQ^3FA@<W:OD4"\26Z-D 
@=$PP(>HD8T_AJ+!!A\G&T563FR:0OC#7+K]:HNH*[N8 
@\K.]53U'B[_B(VUH\HA,<.W0_*&WQ95Z?/X7OJ*6G2H 
@IV0C'WQ*5L!@!BI J-\VS7JCO@9Z+OM(U*7__@!L*0\ 
@$OB9>J(X6%%H]J-$F#L+,4WV(MBCEUD$U<*]$ ![H+  
@LVTPT2:/R<?"_N[R;O0L6N;Y#98.DE]//2&$\@TA91\ 
@R902>*L',.84DN$88BA+63Q)4OT;.0CPZ=]F*V#AH=@ 
@0HJKE-GIEOVXW,V-N6>AQE3$^R$FRYUZ*-U&=LI[][$ 
@2\TN)+$97_N^PT *-Q6I>\&J6.<,"\A&MA,G%C^Z)PP 
@V+]QT!)I:SM/^[&_909YNNG#ZG\.KCNQDGO2!Q,7TPT 
@HX<H=FS[MB8!EK1,Q\>^Z0'7YN>)9>^^\UP>&]=6<'( 
@L@'<I]U_6U/WEKW$\^'Y6J6_Y+"=4'14*V=A6J=YH3< 
@9K6=:/?=*:W[F+*Q9MNL:@D](SG&1NS31B*+ZR)]]PL 
@TN< U0N@7VJNDQ\"$2CY1]/G25>HND1FG<AIH7$=!VP 
@Q[C'<LKSW=^$7HPA?HB3V4PJHUWL;,\;'5T*X&B05CD 
@ \B#3+M&3'XC8J:1#5T_6MRGB %P!:Y^;T3E8F=$LK$ 
@]BA5"?PX+[RXGW5RGNP+1[GG%GFVB ^1WK(]L ]P_QX 
@E=<>PM1]TF4EX\&^,U1AEOIS7!U0SUH#P+J/ ?CN&?( 
@P4O=S#G@*F[>#$.?P4 YSR :.^C=:J1\A9J8LQN<LY8 
@6QH!U2LQ!=HR^N.B>)K(5@RFP$17<-MWQ@.@4!,?,M, 
@%;*/LS :NTQR7^,\KC9&Y6%K2#7WPRI2. G3\.?>R48 
@T>K4%3:$\O$R$!@>Y'Y(S&K^-'W_IV.N%-H3#-[@%YT 
@CX323GL1[-;1=SN$%47%= #91.%_@S*JL*81W0KI:28 
@X5% 6&N'T<F9<QJ343;X%F6FH2\'U?$Z<[\JKTY:-^, 
@E)\$%XBBT;1K"YP)?%6J,C2E*<QTV5D*YE<@1=2Z53( 
@I]X&UFQ^ =9:]=:SM;(55TD@4" GV+T859;@A*?Y\/L 
@[^R*V%=U1A_7,KK@$NZ/)TO$VRHYNMP+6CUQZ#=2"QT 
@D.X?='H*:M.^S-?JA*LXTY8G R[Q!I@^\0P8.G(6T*  
@?2QY&DX.NU6L-6KPC%>1[!5"7@XB1>POA](U23]ADL8 
@@.5IY^\,)#V4%WTP5:_$^2RV$_A^!AW;K][Q!)]%!*L 
@1VN YW#3WE-LW(-PWA,$E:9%^+WUYIR T 74QP4FRC0 
@TJELPA):!2P_C(/MT7L7=:^!4H'SX-^.4&MLE:8@Z$( 
@;5!WJ"D[);44""A69@5[/?NI3>H3RX.@7]=['9TGZ98 
@> W[@WH3;6V>5>3EZP:2GWNH!9K\@=9;'YOC*Z>]]QH 
@]>BW<EDTVYS.AE8&@!DO_F8$'22"'5JO%]HP?[T ]:H 
@CCJFX_,LJ70/=>&P&+@O)1QLG$7ROM,_'-7D0<)K@QP 
@TYVE5\&S2ZWR"O?L!+IQ8O%_B>BL5E%-*()DP<QG\IT 
@ ,X@--6_0'C B\NFU;;S2(&2(H2FUD)G22^A/!LIZ&$ 
@ /\I?5)[ZD<%3,C1_O^F67S4TWVI<0JZXZG=-$+6K0X 
@1,MA%G_40_B [JQMQN3$!9'S3/\]_2D3=\W4E<Q8]#0 
@1;BG \Z-NG*[O1,XJVIGDEX56SY\HVNB/PE..C>VO!T 
@_/ID;VI/3NB)X=K*NZ9Y 21@Y1$D:4^_^!0?=R'-4*\ 
@@P$ (&D(L5B$OGI%7$6H.OSM[44,&L4UA2/^2GAX1KX 
@JMMO'8PB5RXC<@,RQ=XS+PY7D:SI.6E2:@@2PC1?RJ$ 
@PNE:8AI"7.UTT5[NCDTN0$MD!>2($-M'3B$4RV@"(WX 
@5-':&^TG67T1+-4I[W,;0NPPYOLJY::#IZG-X'_^/]L 
@GJVC2M,-*U[$PS=C,W,=DY]#: I3D((A4<U%IZ714\D 
@S_BJ4P*JM-LX,/4*-C;7^5=**C2Z5<L=1P;(9E&C7>\ 
@+AF@,]L$ ;UCHZ-LA(^"_AW8'^]XSKUITRS!<,V$$>4 
@?KNW$T-\(!$OP>&%J"!S<I$*EC,WB&1>Q<B>?23+2;< 
@(!D&,Q1$=TH=CI>N'YB+JH7#7<F&/]P/$U909%I][H( 
@/D<=QD&#_L!+-?+(Q?B)I+]_S7R'Y7OG%/R5688>BR\ 
@U*.Z%T>1F! L-JFWC#%]\?U0'<NXAIQ:9=.!YQ*1Q,L 
0@,C'FF0,M>'H(2]$1"?)-0  
`pragma protect end_protected
