// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
A2IFWrU+gXmjruyqq98RoviLvHzGqx3ZWm+FRNz8mO0Fqv8VX04uaQExXei9r/AL
x2AXXpxjfCfJE4Gj+Tob8vJBAtk5vjR6GeSErkQDgyQDay8DekbW7KoiVrNtLDsg
s0tce6MejNHOfyy3RGo7Ey1EdfMV77vkGP130ZFTPz8cs98veMj4Kg==
//pragma protect end_key_block
//pragma protect digest_block
W9i1024wX6+BJBb7Hpe00sXmSIc=
//pragma protect end_digest_block
//pragma protect data_block
FjFpjK8oa7vDu08kWF+JBPWunKOwB9UJFZYOGKMmQwm44gqOs65zBHBQ0rL45GCT
I7u56hDPpz7Ph8HYrQQJ8ERjdra5ubW4EpqXLYC1T6rDqubv0pzsStlWviDHwXdg
JRJmH3l/MWe0bzSLbevcIzYVJX1rTHYSkUySldQGxp/MxZmLZx78XaHgKPj7WrkE
FmekgYhJCAhgnJUfdZ7kVHmDwSx0Mr0l192WL68l5OOeV4mk7iNP43g5W8z1YsUm
dz+aLr8rVHzXiPtvZdbxhpj2QTjozhE1NMTOQPFOFXsmev3Gwn5wyfglkk7cs+vK
BdxT45EBcY9PYlzPVxJiytF5IChGKGaXXBJfmGNo8V+rJnPm+UxSgZ63tE3XaolT
CtcsbpNV362j/+q3BtQOeQuittQAkyGpsGCDaBNDPQ5hTehZ1eQYKHMvmQ/JjecZ
OhBhrsidDJN0ziboBkjmDBCu9vXyU3ja/LSCMu/k03M50/sSjtLL90fqeLfmblQD
KdQOaA5L72y83lSyYTVl7cWEHGhPpGZic048VvUDC45mlNM2wXxMh5dAXcjTUriw
ycmAxDybteUKQ4ZWP7KX7svhq7LDNnrIuhLdXH2iSedKL9ODlj4v5s2zGYj81MoM
DKZ++osl+O5A5sO68e/9p/3jE0tx1j//mRvWrVhkBSWifmD0Q0hkE+SAZ8t0DrU1
WETcAEyr9TGodZGAewnIE6vNLqVzANysF6G9seeEchvNmyoqVLtVEL0hIBo05igB
lxa6yDa/J9Otg2iWU0ZUpTpvYirkLrnBYWGeQP642NF8DEjit0CESS8x9KAQ9Q5O
5G/ghD0G++kAjfC+UTPlrOjfrsSz3YtoFEpaQfARZsdAe1DSxG88kFx2YgnVqTIm
jJ2hyTh9ufRrIQFHVlu6q4GNkuEVBlSCJC1YdtwZ4PShMwg57e/w8sbfNa0RCVvh
KLGOkHyrhgqdRTrotDFSO2CNpa/OhjuTDelO3KUxELhCBqk0Hkf5VGeANHMvGBlG
10XiFbv5rWZ674Yb9GilEoC1FSlMB4gOLNPka/rp+7dfFJrgeloFRGH2Acukcv+l
csN4MCZ369FHd1ro6ssYO+U2cY+l5S/PBhr+eADT4G0dkZG9OA7qfxrmI3bNAeyL
hi8y/9oNwtXCPXmUx/nGqAVMC1236Bn9ZYBAxrd20rI1MYa69x8c15bTWWyCwPVF
UpzOYdxtj4vVHhkq++YEX+/volD0z4y64mvajFTkV4H+TZ0tpII3rEWVOSSQy2QK
zT4xZWKkT5mZEUnk8otatInL07I45UpxQf9TFcftCqzPlK1ju7RjSuCfS6xZc22f
sQYcYrMenRQCzh19+hKwodcDe6/bIzDx4jWLNAh0Oi2r3IPwCusRrHvUW/u5Wjme
zVaxnSsGt9lYxBwjiNpgLfL26OvOtwsfH1LdYx5/sRRQE0VjWyjfHou6YM/wYCIW
lSWZXL0A81AlNTJ8QYeJyA8N1hgGEKyt+Q4xkfoACQWwgZBNQWkpReWC7NlBVevE
tnP7DfP7lkxRmRhbZ6FA2WM3swMQOotHEbugV/zWHmRqjeX4lS7RoKFw4y3vRkRZ
GT+LPTnODq4ItVHessxRqJ7tbQmIAMjxquoyQ0zcY69YYHkDzHpwPOh8dtmGMito
xlNAlcOcx3FsspAdaHYzQHbCNM/AY0vXn6R/M7DVvJe15YM+F9IAtHyvLG54Mxtk
nGn/Gb1uR0d/+32LfhFf+d3Tuhvl9Kk7j/9SJzxZTic8cX+nrq6/BYOCJW0aPEZ0
joJo491REeC4+hiJsLajMY7ZurYqKRlbgYsebzjQ9FMMsAi+J11kgry8l8QgPwvT
xAHZxs/h3WMmSs6U9lyzhffUXnXDJA9jyO9wIQiwQOD79lUbOS9nKJoMI89JrMCW
jqRVWACOBRBQMyxXqLyPDX0Y0y52L7BNC9okl/Y4YApHgU4hLTW74S2t4Cef6ILk
WTaC3WonJM0CesCE7keoX4oLB+wjiqy3z5TBnbCDyDp/oMMLmFT/bkUkJ6dQ9wpf
TUOlZlysqbrrpTX7l2oBv6As09sFcg6JeSbkJzT73OiflnXz8BzDcrEBxSxgxRuk
Gti+EzTuyzOJ/eZTx4wQ+IxBeWDI/Le5FiaPcuKvXuVFmMgNmobqORQBkgr9rsE9
qUww6bY2oxoUN7FiomEI8ICpiWadfLOJsO1XwWh/Q/y0NBVMmtNp2l/cMo8u1mV4
kJz+R7nQ1kgjeLvDSkpUndzftcXlLWvw1xGzf0XyY4evNRsJW3SM6P414UKGcNpm
J7ffe5n/C60eYsUpWJCW2bo0QZdC2lGUn3muAZKUYwPNc6XUGl9VsDpUtZUxkwTl
12WBO+rS9jfsAMD6tK6ghbBwoNZCNqUKwDn7TDp/NsUYQ8/pyR8VZ6xuo3448rMJ
s+APHhSSpGVkNg9bG0y57AElLBtldPPSBdMylRg24JjczYw//vifi2pzhovEUiBf
3X0CzJ1sG42SL16PdqnaR6Bjc+XnwdTrRAQNuOnFRpVcUXeJUU+4ogsn8B38Cn6L
gzjUN3UklZJEKaMDUaQoTAwNEHyslozuZtPo99dcQ5ka/g9Qp1/iFTy8kVi3qUQD
SHmedAaABaMOzS2sUQtFvzJB/FDdal8QJMfATG9S8owm9kvrgCfA/KreYt/5roor
lP0//aKd7GIAYDcBTBel7Pvx4zwefPsNr6S7BJmEY7tV/+P2dYOeEe7Wl0ExwMcl
k7INyh+Ih4hLvwR7Vos/8cGIPMZxUfMPUVVzVh3ky7orP+f/lpmQOUMkc8VJqWS0
jtlSRwryFu6VcH8hQ4/5MoFz0FqJLMNYXUmVpdFaaCdrxvRn9TfRK2TjUaS7ASlW
rMd3tGX/NPCek/n/CLR4dFPePNRdB3rjOolTnLqerXyFyaxKn/egX7jzXvhcZ6Bh
ivnzJPqVCN4ZmJQFsSEBpSGHvgX1RYewT+scr49SkOlgY1u/l2E/nvg1j53WhDM6
LfZDU1huj9WBoygX/BjSI8iDLR8U197uzRIkNEGc30kou/i/Qcs0wNyZbTT6nWSv
4wTcq89YI63ssttK+PVDuBeMsVdHU8fVlm69cG0TKUvG8nAvsk+58p1F7GMolQ0t
1MR+e/SWWPDUu5uPGTDkn51E2DZmMBy52puge9UOfQtwSJvXDWlhQr8xp+TclOcz
lQMoK7lYNsleaON3pEvDuzLnprFNqCK0S1Mebi4S60FhFCzkcVVSZLDYiMibY/Zd
pqtQb9iaoEAdmus2oSuvMYmnRbz8vbe0Du9yA3/V6zBnT4ZHWcb99lQRqu/a+7Ij
eam6JVS5aK3XW46/XnHRtiJFXYz0UD5sALSjBvn+pTMpozYRRz1MB49Z6Xspb2JM
B5GCPs1leTiUSm2YBLEWadKVKk5psagDzreCVG7xCbM5TxdgqxCWB0s3i/EpgoSc
BDjAEDBpvidOrsi1lqudXQk9ZtFvqLI/UKeXnD9zu43zWcFSw4n11ul1acfS1AP5
d79AIbhzc+svYXtzijmrqsh92J7lN2bCIX7QQ71J6xAfT904yKEgtM5LyqtxaS1q
pNuNbL9ie4D/0rtxP4sKEYAmar2ueLun2dm3RjScjFZd4nXRJPlPtQ0+Hl1HlNxk
cJsR6NDsvc9Jiw7t1Ks9aofA7AF+WMmaKD4ozqaq7M2eByrq/Ve9o62qD4jCs6+f
Wl0SkhhI5Uu0cv5G1jB73H1G65KrIDBNqZjUlAP+hHob2agLUhirhR58wCs/QtK4
2I/RvHjt0m9jzUlKfSOOHjfyMHloz0r3EvJwFALXDbZqlJGqSOqYKihuu2SBW3j5
GiMWmlCSqk2J+YgGLCIgLJz7mHihDtyBIzrSU+u9+9uuI8UWN2ZHbjXm4TID375N
Frmj72rVXiqsbpNAxUpyz82GPLeEt07EL9RX75G/rdOfVXuLXpBUqfzqE5kS2SnV
CSjaTYLlHctjoLp4HmDN1seY9uLFjKEO/d6K2UG5d5vwUblp8pZ6JM9+CPapqeMJ
tjNlUOhTdvtyHwaDzgfWG4UVOIJaKd97HTrBwH504yjtxN6aC0MMVorNv+03DFdh
Se+XK1ic9bfO9sMTmS0lDQa55bkNxT755eSvi9ocVEwdxCv+iHO24rs9IGAWSIc/
28ai5ea0aQcWNcqXf4gNUhHcgdxuILjvc6pAYfK37aQi4+kMVLIotxD2rjtk2Mae
S/GXUQcjNskapxO+rjBRKJux+Y1ydgQJVfpux2gYV/FAed8qQhW9ynSEwmkjvzPV
Mk2WKF/d6DcLr3Nt4676NJp6bSL3o/Ha7wG7xaxWlloCWewsIhO4rjgJI/QLRsdt
aTwJqK3wjVVc9gIP1p6yOgMunwAxUvPinrSsAfkA141ZyOnU43fTJC0+eZmvo4WN
/rFNb/Dbjua8whKR+z/HHwaxssUUglhMspIHQbNLxIewC1iWg4FOIARQCf216qnS
5tjsZjeNFyq6XArtOvR1UStfAJ/tvcuzIqpe8wPB6cGFCe0yn6YD7qrL8btg6inP
ycvuW2Cw3q/veKAyqG0Dju9hj5RrvP9dx8s0zSws+Sk/fbNrZqpApa/l0HXWgj9/
IThY5+8Q46a0DAwtQ5Z4QCP+rn73xW7gkKK8Oq9kac6gb2lPLh/HjGr4hzcdFtMq
ksubXZ+73ZWe6jvpzPXlF1LjGxVkOwHXaUOT92OPDNNV9LAxMqvi+i8l40AQlL0X
ssSseEIHyGIhV3y54gtx6o6ogIfFcmd5puwJC10cwb+DpdbmpO2VawLMheQmg9Dy
GKRZ/MQ4rMch3s/Rh4KC8EZWkj2oTDR7kWTcBzywdqBFfz1ryJDtscubvmydVsWZ
erh0FBzh/E2YpXNvom+6R5Lwccm3Dbi/bx9HIhkk3v1vy+xVGisZX7HbQqbM/jc2
NBqqWMld8Xhq7kHjMjBfWIhypGGB0GHxrBSqazH7w4iGmZ+Tn93XxJfa7JsHEz9A
AOWvIpSlGJvTEJy84DsMzQtwr7e6BoX6ucMhkDyjn7m+oavoqgV0bPaVNiVFtwtO
zWkv30NFW0mdQUASQmsZ0lSAh2qUTsQEKemOMG8Azw4Lz9nPl8/qV3pTlws1CpQF
yNEOONl4xNuQMSzC/yB4Zxs7L02NBYXSWufp8AFzz9zFqbeXucE2UH13lhayZEDu
/o5u3O74G4J07U6INb76Vn0edBK3kzkzkh4hWLJFjMyIdx8X3ful2/tOaxnpYagw
pEZcgxry6Qdf2dJqyh3XnIchaWTlSK9moMn8KzESQku4qkZGaYLeMDbNBg37LRpY
eSf8epKaPEu9ZGjEJ5pfO2KiFQbv8/P5bv8FCHUuyeOircUlyGyxFYJ+LR+N7h29
CvwLrvuF5gbrUA49I3d/Vyue3hCkLI2jgr6luzu29ygv751hpjGFpxgUewpQsr85
Cztt46r0tIS9aELwW+wsvaEvK8I2Bpeht5cpuiVvnSFztZc55Al4B7wEklG8rC2w
KRBa7FoOiJiWEhEjqz/Ezd+cPb291LgtpiLnXbKzpjrp8QEb+oHaflMrkRWtTZSr
dqSKhv236bM8mssLWyLvMslF6VtXqup7wSJ5oZXJoLZtQUIV+e4uX1i2X2sXyjMx
pb1dNgiSjEfo6WZT3KZxnoe3a03V3BudKR9ou19wXZyk9Mhkry/yY3KC0P5dSBVQ
5pikTOL9zyVwhvIoZzKSA07fV8K0tr9wPuPXIrSFt8yB4SXSoWK3kg3NLmzqHPqd
79RN+UwRMHO7K/tNDRnwKZ4ryn18fS+m8+veK21tSj2CjJY1hOY33KuF8LsM5MKh
ZJgZYnEDqs6akQtfII1G29WFmAZ1g7UpPCwDEXxPnvQKeXAay+302R/EtjLQSQ4X
xi5VhAoFbZxXGOIjroZqLtCCeWPIsqgOnoqVPvSV6rAsWp3+PVDVsMk/9nG1jKr9
iYKeXCI8rkeeYG3tWdEpEH07FQDkXAiwUAcQOwknVfKXEMigVcPxjJnod1YGrIw8
A+GSITqNNb7YxF2C6X4aapFlw8bMycZbIAMEvUxM+sZqIRnzA/bb/VIjMnlcGu+q
uMZL9iZGgGQDrJs5ZD5G5Xi+y0knB8K4At0cCk4GqF1cGkhRJYPUFba/1O9sFxjt
N/3q3J0Y11CaA8jVmFfluuPQwhZFxtlx5Lhcbp0exJae3VEgDTx2MJNlXdtEXNL7
K4HaOqc0I3Hw3EEwFe9g4wzSewsXFzUn3HQfYPtk32KXIbv3UmGzvVQ2k5UHuo4t
/uS9YzO7eejNOa9qjLj/hK7/d3AhuQHVs1B6BUWxCRr8o99XP1jNYJyWoRWeFsiz
6INu8YYFPTzkqujygkNXf1FQz9ASDDUzoWzuPbWJBS77mfAhH2Ge+GqC6mBEc5Uc
6uh1o1p8TyfpRjwxCQZElm+ufS2Tam2VPGJnwnsVfb6Y4ZrcjVcMvLIFSdZVYerz
Rns2WYSBYY71OccnF0dMXRmpSkQwxtDRymvxCQ7zlaIpqMKpcS/Z/L8AtY37W4iB
50NS0PAOBBaQefR+QinAxhNorOS8TwRrzaEWFS/bmRa3mpHW+L9vjU9H2AmgMqOo
vnQgoyTMBPUKbQyXcN53DBVSoBHzQ/eo+E4EUz3K6k0QtvT72G5FCdIGIkFEj4Hh
pIl9y0Okirf2sr5bBs8Qhai/j1nrE8eF7lE7jTiqx/Hw9TD4/5XPExqliS9+aZ/r
lXU6nQiC/7Vv8DKt74d9W/TbnwigdpdSr++v9QBeyAMFVFS9Zg6vHivwoUMc2R75
vXnwUpQX91AeQcIos5YMxvhPrEGVl/PFwH88UOx1Nl+VnTPB23xLQCNjMa7tlf3j
mpK3imvMfc92wF2Xe9L0jHI/j45vDqed/RB8OPrytZnZ4b6K9GgF14PG/aZ5v4Cs
w0iD1iNAFh4mwKHOMPWt2MVfBDs4iYepT/2UT6nB/67zNXptEDWkUyUA8w0TdNfB
kUewLDSvqG7LN4M/bKuaqxLPAJnyQMJyBCgrFdVmsSqb9U6ybanXnQyv2Soc+uya
ZFp8mnRH/2MlWR6LHkDK2UI0dgsSC48TZXqf/oVIKMTwFUxTHd6apyYiiGn+z2Rg
kJYGIrdoBc28R6ZJJgiEeX1EjizE5tJEIFI27W0FL1pnH7gmTO7IoQnxBnKYeAMz
r8WLRPDX0GrMvYtjO/VLUwvLO59TKkyLiwZSuDBtVCEgFxxKvenAs7zQBImSulTK
7lScrx3f4xNRkTfIulsPf8XA+YGSHxUDXEO+uxe3FWpXJ9IPSqCBS07CqzwRdwhl
3Oh3vqlEyIPngzFWoxrgVHDvtMzNGGLUA0jknKQjTsIwvnQMfcln95Uyj0x0Bxvb
9vExr2zPGNVjmrnYKmJiP1NGBJzvJFLxS2I0PCm3GWpw955wydXp9ryCP109uUbi
n0baoryy7InFQyd26GbZrOpJ3ZSJ6Rq+/nLZ5q9MaB93ExF1B96+yiDYjG8n09px
1DkCJaZdy2ooVh7MfqXfw5dV0Xm80NHs8smgMEf/ah8wbCMMu2ulqLsukn3V3YAV
R2z0VhRhgYo5aLOe42D9PeAn/7PtAXGgH/4i0TB4Mir8ya8/MJlZFuXh/QN9zXsQ
R+fIabx9b08wEE/9VJUIUdAdHI4xYPHOsQJpiH//Lp0nqUOitiX6cd39rWhlyq8g
XfQwADr6XBbUMAqgV6zOJeUiDrYd+uNj+3G5g6A35rNRhBah9+MJ/KNLS5wF33WR
Puf1pToi1q7t1X39mCJduF8e1ym1Xl8yVnCawZj7TLvbEB4fWsOcx1Xl2Ka+pYLF
6GL9E/qYJrIbYUplIA5WMFr0YukUw/HTc9MwbPCgWSHaBionPI0Cvu9QTOwcyqA6
suBo16Fe4H9+2tWbsq76n7qYQ/3cqhhmdxKFVZyzqkvV5P6ZfrLd430rEoJYq73A
u0i87mdzkebPMMvPdoS59e51R4yFT/vf9l1bN4I3h7/T8PU7MllnkVACr3hfv8pX
FQghHajicv6yTTPUZradW8NEufCbJZPAKyWFKokeChwsxhY4LlHSKYDx7wFZ5fdy
CbZVDPrs5d7Y1beM+YJMip2FwHc0TJ9/2BA7KfuJ0IkWBm47pCDlRlHEj8f/nkeN
XufS67rHqdnCqZihMI4bFzTAcFmx3DD+P7yLAbX9a+XpN9HUrFtQKWCrfykFxcFX
SgXsO6PzhXeFRpBvM34SrPSdWzyyy/3NL26fzOh0/PzWi/6vB9tZa7m87ZtR1Y1r
hYJEUfpoJrzL5wyQhEUGFJLSOI+a82bEF3KZGJbpV+E3dNrUk3LOA/u+rpGZpZS/
mcLN+qLCUKquMd+rugziQ3tLIqV1PRP+F0zl7kiT6TiqglelFcxKr5S9Cxvmb+io
JZttbj/yHBkwA8HhcPC5WBFDsn7NW1X8G/iYG2VH5wHaccmjBFwEASbY0Bqgk0It
B8vwgEFMEhjbz5g41pU5OBPEfhw/Lu6WVvqXn8DZFjGd9KczNpAZM1Vuw/24m9WF
2soPHjgQ2Fan2SjAxmwQJbhjhQWjD5vzDe798N/CFJVf6m+ovQO4GEnueyUORxz9
Y84KNtqZtfZZPFE7uT7CItNDuzqQNl2Ao7GKkRunCst8xxDIS9tSHL7NmKIRVXF/
OtkWue+Iew8sLOF2MlS/ReUMPO16W7wHmg5jz0FCgaDOu93hiklek39QXgFE/Iiu
jFNih6l7u6e+aPbEDrvh/hvME0r2S3Nig5L6bXKWgAZ7rbEg2XzuZTIr191tcCjw
VrArftNSBmwK+jhuRPUhGV3gKoDnFtWpqaCi6NnPMVBfwTZcO4s3586CiOilyOnP
QktzKhVP1j29Cs7lJ0ipAIRMVaTzLIiXNdNzHWE9gqLk3A/6AKoUm1Vs1DKIuH0y
TvCdww0jEBr4ZtA/9R5ApURHRrRdI3g27RjN379Zs0GR7wpGtS1cuZacHyaMO0Hi
RZ7SdQcquo2y7V9M7Rps806slJIGCMvrIlwxjz9XkPi+at2ZG35w1FWhRi+UFQ6v
GujaGIWSk5pgzzaxiQ0Asmnwsn1p6PiDNWxXytRJcfn+dyuItBnA8XErPpphklsj
xuHT+fawhOt3YQP0G3jaOf+p3UH5L1/Ni7LMDxyxNmrF/JjcjkhAMi23YvnRF4MD
mFMBYWikdpRO25rg5hyFJ5B4jWXnJGH6UPm0KeFi5eRbtAT0J5jpyjk812APV6Xy
BaEef4EaKZEo0Iq1MddNOiBRzZO6wUtqmPpafeNzuv7CkXSJXgopdNLeePnDY26k
hBRihO+UsYWE09Cjl7ITdaWOV9+a5KE3crTyUuvlXbXSmT8yD1O/Qu6Uca2HbAey
Zy4HFKztsjvfqKm69ghoc5IObi2Hb5uXDnDtQ2O0KpX6hfEg1VZAJaRbyE+vFY8V
1lfSqYu13FykexHF+Obx+fq2CbDJzbROuZySx5poXvzgW+eiM9XhuehGYvLL+upS
f1yt0PhXtp0O9GGbgoUE5VfvuYfXe276aQKOVHdafgBqv2XMBcvAFuuXkJn8PR9U
qWtY1/L7vCDFTF1JIs7MTL2nyOC78QLxlC/TQpeVg2IO6azkdNNXUgkka81iChyS
M7/V/1uSDjwVkRDthnblZVihqi40ynSCNzHdUQfymMW6C8gWKqGpt8XUXRCRV5gN
zCJLqrA/rBqw4lbss88NWaXD5YsV2RD+2FP3TDVnkBIWb/VYlKpRjK6pvq4UeOX0
i2n7GjqBNUEU9DjGxsH2Pgyfpb1f56pVYJ4uIwUFqTZH/xkv266VV86u6Tlxk0j9
/cpCq/CWB62v8aaptuAMGX16Y47hiQCqrB1gPCnbLekK9CmwwEmPpOmH7P7OW2LG
0DdDjIXUtl1A25NdYxsfxoodytUgOTMWujtxLc7ehb32aEG5o5EhTZoxrIBP2r6i
peCu+boTEh47bf9raa65I3D/3FtnduXutrMwQKDvJ4sAI85njhbkf8ODSS4rqCrY
6e6BVoS/QmbD3ui3FnS6pbwy+E96cOyuFrZhibeoYZ6J/cdciu0lP1lXDJOl9kgO
u8mT5XAB4Z9rCyZ3PG8Z1qh3LAha8oIr+t6yxClFahK6oZRsIBN3/Drzk3LrnoYI
M++3CAUdF+7DG0l8jFG4EsG1UYm9g5NXBYHJ82MAMrmQtoNj4bpIAEdqqILttSS8
mRTDkGofsxVJtZspsDubUY+POYzRE09d+9ZDuduGWDKmQEtOJLw6e+6Qqg3Ihm54
ww0mIV7FuN7XgoZl5otZp3fUnPf3PrtqQfsThgbKlYyMOcUAM+81hjfsq/6CM296
3OmYcV3BfY3Y08Jx8T9TBSuPoCHy6BN9lNaQuViRh4JzsyR3AqGpVbiGXurbKT60
rbWXRo3Xalfd2Ci7rDq5Ma2E0rDOWHen7Dxj82Qd9AMrIHIL01V8hY1WuAigSdsG
ei3QNrqk9o8YXhGnHU95zf2HTHTdHR7aHg71OXyNXVZzEi692QR6Mhr0h8d4+s9V
foT5+4kBCV0f+QLbbrB6Yv2QNyoAigdkmENkz7bpwCu3c+xd2bgDJvrTz7injN0l
pJMlfnpcIKcke27Evnh+Eh8gwwQoU+g++YDIgI/TOOqCT1AFDCFqXtB4j3K4cqF6
Av/d0q5hRahTPRgSmgI5L6e34Li3bqdH2oYqTBrfQ09eWELnUqU83Fc6GFMy+xiB
UweU8PgqS9Sb2tlTcBOH6PtdRuBeqmrYTCPNH+lVFBSlLq2yrhWoDSqfusO3u1Kl
NLLi3dHI1vDtuKQpoLkmXYsrBXtYb3llMSrXzgiNqQypFWYOwqtVS19dxb+BKbmD
kZP0/HYjQW9Czl6pSmRYWkZ4ah2Q+31Om3ytWR0x5bcK4RU86lWEMoAtJ3ua5yT6
WfRfphLvLdkq+AeqCKKcAU2oMBbaaNlyWZ47BWL30sQiDeqcgi9zR6B44m+VgKnK
h+QRzswPvHmYiRsHoOSAk90Pf+bvT5OFtCQmXPRUuMbUCFTZVIe3TosFSPybJZom
8jiM1aPVefyAF857MOywlOGV5SHfazfgFWLABMqpN42mMxxn5MZhTuSeKf64OZpQ
azxAGgS3KYIicvkVVuSumsVhM0DiywU2Cm8xkOdleUGj/LFjvvjsrcHFJ2SkJy94
iL10OwTTAAKNB53uxsajfghPE3MUU3GyTYa61zktDtoFjjtjoQSKxR6Ug2xzDwci
IliBg268bxcq1VnT0Uo9ynRa/2SlYXfn04ApHnkSXzreN66VAZod5U/9S9m885gr
guFlDm0fCRO34Q5Yc2KYcC7Ft8Rp7JmNRyNTMCDJeuZBj64kImVUD/taRnxZin4s
dpxd8zsQuHIBzyRhIJHFYKrHH0ldgCXVGzOPNFLuEP3/04ZgNRKscxrCxbiPfAww
8HMZ5yk6iJ/TnBKrl93knCJQQ8xqrzpQudVOXsx6lzKb0MSuDu9uDhmA3sUanVx1
OpqO8lXpR19oJX30wZQWA2uN+TSIKm8u07eKEcR0Sbj9d13kfm53Y0r+VU9WYrgN
Iu5arSOrkFlduB7dc5Tb2iWGMTPwnLbUfOfa8PV9Q4aHy3ebyLJAD01ymX2ko0at
yPLckc6irdmtmsGd8gS2+OEOoJFE4yrGmcTI6Y+lPTDMCnCabL7wGESl4qjoSpJU
Rrt4YtBVCto1joRejo2b2LhAVuKfI9bTCFhQG9GJMDQCv0YVuIqRlyCZFQD6ItAz
ZNaM1MJAAIfJ2WjiDuZUWGhr0I5GA/J2Jysnyt9ttI8UBvmzC1JqYnv6FGqHGjbM
+9HQwS927QRVAGP2RluFYpfX7ACRzK5lgSMF1Wmp8j0lmuX+SR8HwdSPLgT4Xoi9
GLd06iQFgs7h5AChLyNoL0fNSt7EhvNAt+0RyLeSl2v5mVnWR6HPRYKvZM+ZPU/S
vT6IKJGBYxfZNGqFkbU6LUqi17ehjcghac1CquPTAkV02R4QJqIcAPGyfe/w1ZlD
zTdhueXeAuujD2iJSkK8EIvFAYFpWjyo5UKUeylMYLOt0lFUQgBXWNdA81h9XkZm
Tf9CsvVjFTAVVTKNAwWMmTRnnL93vQYVk87EiSrMrVHimBx9qf8DINkkyhOBdFrQ
vBJ9hgmfkM1PNeUhYvisqiL1PAVyunAASh1YbtVDSVQveeELByRf+2dkW4RqR7Py
5gk4E2g/amDZsyypUnxkGBIi3jmyQx8oLuAM2/hSv1+s7Me3HX3oKmDgQf3HGWvW
FhL19wdGVYipMc4X3YEpTiOirGj5kB1vZBgnYzsT2ahadUsQmW8AF1f/CSxk/6Ga
wJS8JBIRqnp6ztoX0MkiCmb0eC4I8nKVjlNXJcBxLg4hdxCfcMS2OxsfGG2RVZr3
kdoksXUKxt/yZDSasil2luojkuaCIv3CaXfeatMupYr97ehYmcf1ErZ0hjqZnXWw
dlQDpVO4w7XHPrpfYdptlfVps0bS71ATynsos5I41X8kV9Cctb6rGefoK721uDqd
KjwNAJcyliHzNEexoGa6mArtUEmpOzfSvY1KGlY+NLop+IMcn4pVa4nwUM4kmf0v
EBGs0TaTyURxpvcXBCOrz5z4/reEK03/9072TVShFJV5AhZltUEpxwvMEli8L2FC
a+HdCVq28L22INe6/5cTw/esgDjH84wCCTfNsPqoBRAI72ECpiR3RYwdbMkcP4NA
h+o18ST3A+LEgEFrm2b6kG2VcxSf/l8NzmDBLmWXtDHRAWKJwR0wV4r8qce7xnwV
7sQ6ZIhi0DI3SN4DPMsQXThZ/MzfB3weZTLW/+ZtDveih2aMeknvDP36K2qeWJb7
hMCrGTPTd5K9u24Y1zYjtKoNcoKzQxJy4awtUSyBr15SwppoNvmB7tCbj+N+pOxk
RfkfurDGSDEli4R2Ec5cixVzug1NgRr5C7gwVDTjRfavow5PXI1iGieY9kbCEM+y
0xZ/PvCxTDFo6AR3S5YNCaRjry+b19VWp0vbBlrYI/iRbLouHNKDNJ5x5bvDlDeV
mHJIwkkhsGoq1A16rd8uzQyIWTly/HTZfox0LqfnjUENlSv/90Ci3B+VhmcCcuzO
z823iBfqpK5kn/hwOcz8a4sKDFz6nCiI8SaR/BWJD/lfivdM7tM7VptvJaSti/MX
Kdkv7/APsTL/xrRLDbneKWiGJHiXDbmV1XCztDKcrkOV624GQMuZdHSjo85rzC1u
UNYbbui2kLj1oB0T6boMCBOGvWglnHyNMvwEaWHBKFpPt6LjydwwviLTN+GcrBGz
5oKEisZO3kNtbHR3ubxcwEvek1smdqASdfetnM58uVjmwqaznSRdkH05X+ak/+YO
MmykiA1QazTz45SWFtmapay/wFn2mb+CAVH1GB+H+ew2KEzCKAO09xse7zf7SNoA
lXKTRWjIVJll1A0BJo3YGWIa8JKyZ0Pdtkxep0OEuMFjaA7pQGiWYnWlPDafJTgc
T3Qgc/Mm3cFx6sV68zd1H0RP3P56rp0iR9g/4BnlIFvKcL1ONITFia8rn2i/u65K
JTTc1+WhfBz8kBDMqkFz5El9+D/g0DCu71i1fDn1MCanverQQJkMG4u3nC5RKTIS
bZHNmmDd8Wz+v1RXGnZjzcK536BuoEz3MsiDpnPbFRPyw4Da6nJsYD0oObhGD03n
pfz6UXA9mIutrcE7WgOVyqGQe1F3LgpQvWddrDH3CLyZhr97okyPaCtEcRhEg0Ec
ptYy1Vx4A0hsYVshind8L70iT+D90B9ph11VwRr5yWBaOFDSHAApJQ5e0ub5rwMD
2DMnZiFmsL6OvDZ3pFyizvjT/QjYb/7Emn+2EEqOPVWAypjWmtGUAb1ilObVTIaw
LFmOKhD8asWwcdGwM6xg+1w7xrN+JDOAJEPq/XBbWoT9WOu4kFRlYQoWECbm3xrf
+MDugDgE7aEvhsEUDtRNoJMxhq4JPa2ljq6mIXh0Z02DudfR+PsTR01MzmP8sjtB
SrU9i76SUV938FSisGVuTDuGul7OOnejy/fHYXgwmHap1QoJvqiv6P+eeN3mJC21
puj4aQ/xMdiQRChc9ukEVIZGSYHoQUxpZpcWomqAT/3QP3T+XDswfiZr+AQWBwvO
B0L5HS9zWhxO8PJImYgJqyavBBmafY7JArUvyDX3BQbETddUcdS/RhC5o/N0DhF7
mI/4kPwI/vhV/eKDKid+d2LwF7PeVABrtlqAPHmKdxPDBRUj/IuUNY+7hhArpn3d
YMYdCQMwL8I7R6KLUDdVTWY/V10uH0bnhiffpxLVsCYnjAi7dwfjlOMljpBwgASn
oVztXB0bqEjLPT5qd5J+aILh0F2PfbUq/jHaDFwVWgiPoHD4Zp6PKOVWVbOcrmzc
ECmWgm2gf1XmM72lW9oymc0NWVkII7UAkWmYdaKdfm3mZTVa6A/6V3+T6ROj3SVv
Vbg/evu0Xr2M6NaRHMKL/4e9AjQX8Y8O28MLlB1UPYer6I+fmWxqoeWI6erl3tMm
LzWFfbpgFi+JM14l78YU7vAShg2XoYEDthdiIBGA9a+/lfSwcOkyK2fNoomh7ny2
ZegtOAu6qo3AL52D6Lv8cLG3Zdi8I0j7IJuPnqUEac9Rly0Xj9LNCYh2zzrSgfLe
Ngf5nGpk+t0sISZ7Ty7BelySto5W0jN4QLve++BxFqlC5h4kC9rE5DMvcuyMb33N
b9DdFmawHH3uPS+vDaYewzhj7hn06MF1wAxQ8G5QqpPEZnvd00ZG1Fy0T/OQ96Zz
zflxK9pecRc7KUE0pzJNguEkOy1K1CZVUCyR5pKdERH6vaQ4LJAHWwVl1VXUMvFY
LlcJv7ipHvDAfk9NExJ9KhXyA1FQ6igKQxx8HYXKr5LlsGTMDJ7XWe3bI61aFDya
mW9ylcgKxGWq8qha74HXw/gCqIH6zUQzxabWwjCfgPZdGeuZFfMGyU9e6Le0RCDF
Tssaai0+w0uxxFuaeLxb9A2NzPpoq/+/WeD8cdhB8IqZCdvs7hKthlJGmg2HnICf
Mz9n7e3oABFk2wx5cPnFf/GXkQcM9x3AB9sBIcmZVzfZzUbGNqJDnN1sy4E4RW0f
fOOsz1nSMg2RSloeZgTXf3B3VOQA2i5h2cgOZmdTO55W+NtefBnIayJaJixdcWrx
EbFWwkBktJZJo1yMqoSJyqDK4tjzo+3MWKxfvaZfqZblvMfgWf+oDcsiaE+9N4o3
Nc0mmQTDdjw15IlFzGjt8qEvn+5Ab/XuYe/ucTkvwRs+oXJpXkei1MuzQublrIWR
NsYwJsJEaOuTj8s+W/NjPsC7tYhY6LVcITZq6borNuWeO1tr/XpQvvVdJO3KaCDB
422n5aIFhukZ+2GQu7oNS4UhQzVRS5VtsnXAzurLI66UghUfEyX4fccNmBDRzv+s
qBzZnMDb1UoBdp+Tzak4i3pbZ8c3XOdKZgf/khH7hEw5kaWP3gVRZEb+DFgZBRFj
QAZxRHzWMSSppJehf5CudVIJMr1MCHMdH8u/YweXgKaVLkcrKc4ek/idLYoKhTgJ
L2ge5BsTTDWNhKMQ17QGBC3wrpgAv115023xceOLXdeUSqLOR1gFck0P4Jn3Z5IQ
l3Zdfoms8lZwj6sakxcg8Rg1mxUB8LUiy9tJzKtcwIJKDS9mRZhj8zlo+gxwA054
MzpNbC1B9Yk5HJz75xjLe1RqGoqUQkXvasEsJlHCcIgGKSY7Nyqy6+xuWQiRP9XH
+pNag5rhyyCZQDMPvcClIkgNk4pXtxG6ymDBYlCfWbCQPLgucvwd4f4ESvnulPuJ
IOIYNTK/zg7A7kFdMBHmyDawNH90QeOOXgWw9q+NW/pnTG/DzgTwqREtJlt34gBQ
nfCTXD+bGgBI6CSNQgUX7SoVcHePUaccbENB4p9h3hom3mC0WUeGbBNAjaMpQgxi
0jkvow5YEdmh8aqzQ4Kpuwhw6AZkOZ7yQxS7fmkuv3tVpMLEkBhCUtmigX8VfYPX
HRV1n0q8ffPQutAUNK99J5PpFFru+UcG0YnzXKXxfn+Z/EjwP00+iL6rJBa3s8Vz
g7hthRl1R3W40yfaqQE7JHlwn1GotEpesvNr671V7og+aP6Lycv0xp6Vo6AYoOw1
Y0+aktrlARo9qiPcGQG7wLo420I/zPWu26LUlWt9EKTWhbaH5C4v4IWT2fNmxMs7
omYYATALFbUJRak5oW6TKwo57LATH+DCurekNcvI/W0j9SCd6wVR6NfT0pmnXEiO
wJzNlrTOSZ3/Wsbq+c55GUr0lCo5Lae88mD8bXCvUGSnKnsscUrVFGsbO/+L2Tmw
SE1RNctAQxhXCSs4fVCyODT0ZJcFelzmKJNsPYWANiGeAl/MwKRCczZ/smf4R7Ep
JzGEsG2+owkKZ6wAoxBRkEkEGXjqEiRmpuhahUwRh1bkYLSmV8ZNaMbIzU1SGgxP
2yDHZsZtwmS1lGNrrE5Q0ZQ6ZknoyCgDBKNh16ykLfCmjDV7OXpTzwqR8s1tLJTd
uwojAhhdMqcs2un3+Rt3dJjATHNseeP6JuHLOiZoXJYn+HVDqEAb5b0my84frytR
ABLxyDZx3MrwRw4cF4x0TMVFz9fGSMqaMSUZIIJVFju9cAGCs20Qt5NZvwUDbdEa
3MQVh3i3cbZAvC7SkL0HunAbCjki/UZSrRVjGAb3bgyBD0gFBHEPgJBpvRWyYaRs
4qxGVMWStSZ5yvrkYWFQyerfyS29vUqHmZniLT/hnnFuDZ7cmjmJECX4ThBmsghc
VUcX2RWma0Z9ObgbDU6Gul/1PXGb6LqUU1IwI01EAIxdW/epIQVFsE4Y6s7BL5l5
WJEvN2rha6Xsa6Kdn2nOVo0zMAiMNvEzfFw8XOUMyJ8uiHG/SPEGhtdStfyPv2UT
2MXc6/bGhnyuDOA5q5kwBscYm3sL7jpRPnC8/C0pyg0bHcHhBaTeRiRVcCk+FKOE
ItMY+hpNlYl4XM94JgEm20zuaIymeDLGVS4P6OcTnpJc/zNgvc4Kogs2LYYpVEsp
K3A4u/HStMvBljn7kVZ6AnVR/zcxKYPltysOMPyDo+zL7+rm++RmK6UGXhsXbF3a
rgkzVm4NCelIfN/10ClI/DXGbtcZ8YVYjrPdp/ADoB6uDAgx8A/UwtEYOLQX0E/w
2DundSkIKTmxJhQzAgnRDcCafrf8WsLmpMxdZN31BtXcnH8UIEW9f7sMtLhmzEQJ
OaGv3p+xtAlWHXy1Q0mp8rlZeDcVLmz7U0e5Q3rZGI92+tIToNcRIVO6U8kZGv1k
w+Tt7LOigeNNgLN+9woMNzOBvBj1OEfZjBUSpcQ4ZOSz6EOgjYMBJiU+FJxbPowd
Q3Rf3vZPQ5b/wPyIRJ4gferUFcsxK0dtUkwwu3d0tk1qE+xTVW8Vko2gYeSTVqLW
mJTOIkdJcmwQFYQxj1jRISx3p8Pkpjg45jlk8cdnIR3+2nL4lWF686AwMNEHmggS
WXAWANg8URYz7SIuwAmoRXuH9JEaBpPqmlDLK9x4JtcinuNkVg1eNm9Z3VCW1uK8
Z5PF5znGn9A6qgvpBk+mG/fP1aoxoO2fPjS38xFrb74TKg7gXMO8p1WOI3T2wmPp
KVLDlplCEjhs2K3M6tBKG5VjZW/UsLhE9MiyyGvLDbnBSKbnui6/Gu0cfIKNGWzl
m0AKB0C3UlqO7Wd3tdwYSSRtoBYyt12EQgi0HiD6PI4ZQvCvAqOEOjHl2DuczrCG
FFYvtMmbbHnTFoI8kW5XZ2oku8Lc40S7j3ZdG1VLaN+dRYlVNW7GlZBL7VQXdIMU
NylKF5Qn5gNK55xpT2ASSC/x3PyGdWCwzK2lBkSWF/O/DsNdosYqASw1AsZb8hOU
+UOGoiPlwr3GSm4Oi4dsG3RAB7OrI3aLFDwTHOrnJNpfViSOK89aBhT5qs4SambG
DddcCa0Um0zpGTazneQKCiJlkErfAFB4tMjsk4KUQdeKSIf70/bW3hYjVDViSEcK
zgMJov7xRLjArXKIUsl5kLEw4FzjRTNgU/KQvyQNlQ5PVayYsY64WurQa1sqLSpj
9cF2hRlquEZXGMfad25113Tv4wELS/HaEQhcGiNZJONZIaXmQ99EYNq8zAR62Wxh
/sheRGzyoN1+v5RtOl60Ygee/bME1vfx3g/zEzq8DJ3AnzNQxnsgijpDlCVPaa2g
Nibfw7UKJcRffgUSp9B1PNM4+GorUnfiKWyTlkCharib0edBsnioNnJmo3nW8eAB
iyNXafHtNijq0iLVq/ubkWa4mdd7vyWQAvGkpNwk2wTrmuFXaNevZPIjeQ6QT/1B
JxJ4JJplfwM7Lej5EVuNlB6GI9ajI2Gj7Ds2Hws0pakTW5EvojQ0MtgAO20G5jn/
yRPFSHfQRSF7vH8UGlwsjmN1JZTYgV/mCT6+a+u0wvYqwLhJVNcnKNXf++OJZS0g
9jMXc/JLTCKQWvwWFGUDSoGyS0kda5qMb53QdPVMEfLr1RTh6Wmw5h6LvEwb1Nac
ltyKzqZtcne1Z2IqTMARwLwhOBmnLgyyHCy6dbn9FDXl55kOxrE6GxyS51fEPsU1
l/bCZiydl3Uo2YaF5CMalzFKwwKiFOEzo3Gpj/VAMEsJV/PEbUIIeVjvthRglTZG
Mhuo/IbWhEqPtu8kPEWtoLGJf4x/Usm9/kzeDuiESnHDRRCICfNrJ0JEhSCyDx30
vRYoA6d4V+bYG9PbpvCf4c7VGDZTzm0tiRKzWBW8eWLteWkXOnwqaLA2mn6T0cMh
kr2mE0vLfYNjNcRrmzFaWymzobuSHXEK5RVMYANBBkzqAaQNPLTQtnezHyto4JPO
Va6Sav0SmpPwljFqCqTLjreye3CeA13R1HF5P+FIv7OjZCLF1H2l50CUVzCkcTrL
dxqkCA96DMYekNUwNGnfy1l2yzWuH45yY18KDonrw4NKDDqBlPobCZNzjDDovzIQ
z8tzcLD7cw3F64IeDwzfEEvMgweiNjCEWHEonoTHrz74pbc+6Qs7nWXeZr28zvOX
DqETeDegfCzKq5VZIrzAU6XjjD3gc4LJfXdiJjSxqwTA8JTNbWNFOTkta6Xtdn5v
G6nEXdiiO9WuemQBM0nVCXykKono/IsRoClS/CbiGA/AUrQr/5nmRof51BsHAiSp
8bqMgX2dyPU2NQ8+xF+5CQX0IgQFbhv3j3MMztKYnWH1hN104D3/P7VQjF65F3LT
zip/a20Ux5D5GVhLXhybvYjhIwkaFiQuf6yypOMypdRv37j7z1dkTaWgOIBMpF5p
JKlrzuGTfEzD/CSo6tgbbvN2kuWPWHAPeWQYkDoTgb1FVoO4yJL155YfJUBLb49i
U451B5NQH5TW/jnXfhKRLx/SUFI2+7Ebd5d0yTNxDlomE9vFiYg9/ngYDSVTj+tM
gbF32RjHFrAo7/W1Ud5cxww6GKeecY7o2Axmln0NTdVfPAqw7Wisjl8ivWejyx96
iobYMyCxfFIzAzDtZ2kZe4r3vvDiF7oZKu4hEKij6/VMonrYhepsse03XRq5kLrp
UAfUdtfVBZB/8hpkITDjAJL9PD8Ey88n3jM+teEq3ED2O+6Ur+Y+bKAAe3nTyCsu
X9eDUZg79bjyY0V9bYi6neZEsNTFpf7pahl9YmS527NJA0+35lYcQCOyUCzjkSHs
EkUejxIXK8XnucTd6d7me3fMDAnU+ea6kEsFz8iwgibWxBZu4Fp/z+DDUb6R8F5c
4DV7MewupM+Re8tUJuDzJRtRpHDuTqGCAV22JbXDweNi76ULr5h29JI1DQSlDC/e
k2UyghjOxy1ofSd8ZwedoyZMilSQ3pVi1YKKCh8xbd1O39mjH22mOvRlQcVaaa2a
ooyJGs5L4FnVeXyL83H4scp4nwXiGhbH6bNgVYJkP2bYnynV453XFxVPJ3tZi6pb
00oxbHyBlZKyGn9LKUWWuLoTN7SEkAfEYlSQDO/XoQy/lr1Rw0V5anKF5qE8p5yt
HEDOk6DGGyUQXacBcbTLJgiwdLZkD+HSbyIT9+CE1EPf43FqujTZmAFCz5ycjhtj
DF5BzTd8Qori7+zUPg4c8qqACWSqKmQPlk82P3z2Soe2nRjDdz9QXI501naHA7QF
tWxbE0MbuibZJPT1PxuWDjkJsofXCUsMN88NcGRqpjM8ZhI3ex2y7sBUzXJWn64B
bosaRbDxrfcbnTL6brdFdaQ4c11Pl9cqJoaQIsNenf2ognoTZVt8LfOGfr1Q5a44
L8RZ1RAHvsHfwGN2umjqiTO2I7OwCrLCm1O6Xw51L99xfJ5wgRWkp7J619ijdl5u
u5yUq8hmYau22Xh26cCwfOxeFBRBZIJzbg5OgASMMGcxphUNuWNo0D/9mRxY2hky
gYTV6HDoPKdfI6FdIo8JpPRplaK6O5xV/qjGCT6PhWDUTzafERqHxCBIARtwqww2
pVD+mKSAHuNfnC1XJQ4S1Yjkc8ymS7J47h/77iUCeJsHw0E06QxO7akMWLahalDh
taOU0OmUo7RZGISTg95pL1DIk9TaVeT7iovrN4RS9DfDnvHqFXePtZEyeItTNN58
0TdyIqkOd6umts64hDUq1EDpqtHFT4GX+EcY1hcE/hRsRows4Iwj0ll4qEMKrZWd
6tUprFGuFV6zC+SEB+BKkpu7p8Fb5yPsjxMK98ZWZumJ7rD5SxgqD0RtWHPXiRIN
JUGgDl5jHyC0CpGmLW5kAxmN4UCwfp/f8bxlr8S+cs+K1RW/LDVUXb5CiC/VOyCP
8HkI5JtYLceGGlBczrjr2lDP4zfivSQfCE+xQblSWQpQKYqcaN2GCQB2maIHZ+p2
fUuIpNcZf9f+6Jz9uLI3a4kdW3RvTE8aMHKUNjZWGt1JtjS5JQRzuPb27cNn4URk
6FKE0/xru4EuV0BuSQ/5yKtK+6q3fCy3nrEmimpeuL08/U1rVmP+fw8SkR2Oi4YW
NJ3MQzXGwwRVnASdC/K8bP0p/tiF984KaHimf3IxH3oHpHtPQJih+QZFXSsh+Aib
e0GNmV+HMBqxWRL0tl7s6hUF4B0nWaNutsR5dtyxu4mZsAKhDLjVUFkDD3ufNHZg
GzI5XV/OLPIoMc5h0ahgBAmSU5edp+oWGquDehQ+jcxfonWewiwZyT+MUulLeX+r
paRaga6IbLErBmdkuSsTR+We0q8irsznYnFigjNGdJusLrJVQGL7J/Xkz13loHDz
L/CqEOVP6QzuTOwMbSYkUikPEPL2YYSJI464G4CumqhKM/q6n0OIVajCi8mj1ecA
4YVh3o0RP1hdx01P5158HsoglHfiP3r0H+4J5i4BSZrSXNQC74pUtpLvTrF0NQrZ
8eDDtPfRBqVcMV09Bf/nK+R+d0HA4E7w2vr1rTpDoueVbe7x4/yAP89MUCyVAdxq
KVluXzcUL4D1xwtHl6peT6saNhK8f00oS9J8xWiB8P601MHXEtnLnXOfnNk/f/7N
s+8mXT7CIo9F8suQyWmGb2y92aa4zBaa65mY/sYklrNkjbIJOiKrlqbmO/ugiHoH
H9XWqAKYjENY+YM9/E6VMBzVDKZbqY6cpWt1QRKV90p35umptqtCvPCU7cpE0EiY
UF2ZXJFR6nX5UkNw9P72BiEAtujD5N0g5PBazak+jnIOEPPqO19tsDjtBU7S2V1f
i7LRvlSbF3vAciOwRvgK4HW+n3aKXSr9OYIB5eXJ0FyE/Rb45g2bGQoevVbXwKgD
HH7GiAjDsMCr/1rcwNbynN7Hw/SkAFCd1uwjhW5YsiIVw1oascEw1Gnp+CWI5KHU
XeJVbx8enPKOsLxjqQopYtiEGlmWSDkcrk4XgDUflB3EcLw00VzTObCn1abkO7qG
1ISiuiHLTNZtN1gU2BIkwYFwjhWZfxq8ONpfqCKDdw8MOtmi/rNpIERV9MAPt06+
EKkDx9Qm76OD4TcUTLa+GGFx1ZwBuchbY7yRny9BfUB7a2Bu78vjsl1QfisyBmWp
2IOA3JtBXYt4hwD0+TNCPM4ugx/Za6+M+IZ3E/6mKburepwYo9ZqXemEUVKrhYxq
OXIaxRz3tkHqvArhJvbPkfoQ7Q/HA9HOUjILrEpqGGiM6Bu8/uwDTGcglE3qQIiH
c8nMxWeWAxI4IUpgtYxCYtyhvo/JVILfHh10d3u4of1Z3Q6KZ08YzcckPg52amy6
Tg32Z0CmdOXUrTMakYjF7OghDZwDQk9pnGxB90XSOtVyE7lN3xzsl/LQ1e7Q1dbD
4mRAQcMvtd1XeqUMSdcUriw54TrVcqkD2SgrDpkreJlC2L3VjStRnFVve5ind5Vb
zVmT4VjR7Nz+mSEQba/bIaZXOPlHlbNUCC0CATA0pGdcCsm/nWqE87PGZjj1cEqu
wAhyAfAyMhby+isUJ+eAWO8aTRQWnVazC82Xr1lC8+gISR+G8Q//UEnKjPPvsICY
t0iBTNf2liRQ3AXu9H2L0VcD0TUKinVAU3039RZx5LupFtsIDUxRjoTFT7h1Nqtk
eJMrOy9o65azvnqfXLRykIzBTNjyhGB/UfMJAo7Lyts+ePPygtOkLdGYe8Kf136Q
kMzsuQuo6r+4588UWyN82VTh+RJrpoZeVtp+q+vQcBW+574O8nwvaKAMNchqDlC9
Qp0CPnuwas+IEpUknEBf52xb+O2T/HaG4FRxJ/8/Mn2hWr08uxTV/6cWp+j+VgQU
Cnn9zHFFYoI3DbhEyoNvMEODgcTqE2f04qpXoTGxWYL6jHjgEvzAGRYT/SkVBnjT
C95xswMOLgi4Sh/i0H/H9u47pTQGlvOM/MP2ko+ZK31kJ16hkY/MTPpAPV0uM98+
x0ByyS3VEMlR+jOX4fxr5s1lrEhS0CrWtZoO850pki1j5q+lwEEvUepOiMmTzMy1
wMcLaKG3+qAnvsEtenapWWMm9ENO3Jx3RpVkz2zwdno=
//pragma protect end_data_block
//pragma protect digest_block
ABWikO0oxEMNwASyIFCsKGdQWP8=
//pragma protect end_digest_block
//pragma protect end_protected
