// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:00 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P2/D4PX6iCoXHLqXDq3eI68WFJ2hHEAYVVVHzcnKwlhKCVxUTr3Cnd98zo0SypN0
1EZN20ehlLazrWxAWL7PDXS50yV1TjSesS6kYkqG5M7eYVAikXCARzZkqve0mqZI
NAhC+7nJEROpi3vgZmPlzGGq1MbRH3hPZTaY03Thw3E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18496)
b8PB58gGE2FWqINNUgLvgD2nPwM0zkmBA84sdhE+gwzH+Z4WfbywHCFtK9/rV1fx
5Or+/vstDh+kJU48G1c+oLKpLw2QqAtQA8DeP08RAGuu3dRcx2IdyPR2iw68EkcC
VuT7MxK0Pz3PBFICmsi7gWJKe/41MO19KHbgOqDdVLLfPVzVwkn3HMvDanQz8OEK
iBqu5p5LY49o6NRGNra4ZTYRx7w6hBZS1UZttuI+lvLsAFBGglsadsCQVCXNHEvI
v4D6F1o9776179ODruQDBBxHAi2i7KhktYlqSket0kFfJh7Uvbv4OGSzLDKM/iIz
U3vJG9ImpduqR3peRXT4nnmGJIjihQwRJj2ui9lmjwaQRSS9hrkSIkWjruijGRWE
HeoDcuFGZzU2NTP+a/nPuoe/0YYexhc8qEtjS3hV66O5AvGXEi2iFTL1i+mHw9I/
kf3OeJpctj33PhCEJaqingHsCvModpXwY0bXQcC26Dhxp7DJSjyMJl9Uy67Xy0V/
rLxe8+wQIVpMLqKHY0UsR7rsn/66Hr3rmoApEhhUeutILpWlug5XtiWCWmvsYBiV
hKy8xn7AdHkEuiVKjyNTq2+YE4t19E7Z784rQJp/ALeXUxdIUO59nDD9yVKc0NsY
syusSBQOMg+DnctnsNz5Wf7NhuLeDGL2mpapW7p2z1SNRtaDQY40LtIsoaVPv44v
NpaJJiqIegl0MKHmKausJazme0lyCE7wF1TeSc71ho7KhYYCknzjQy9qElsfRoV/
kFtxHMW1rUZDlhUGYKknkAwdcG0mkWSzr6mcLjZ9YjrOfvc6pnN4KTcD+diSJA6w
fW90ul0YYGwEiLLHW94pbWDaukR3P3LJNun1BdwynCO/JVyhBwadovEykxHeNtIw
swyxcUY15Gt71NziYh9HRRCum8jDzjsMnc1Rb7oBpPpf25qWYg3UuBIWTzxpacMU
gKUmHBX9qlIDaQVNtXqG8U9UXpcgigOjvMDrk5Ms6ngsmuqpaVeyyIAmpWz7QokD
+sWHBEhbHCNERJxdO8jIhM7ASpTW9K3i91SYr6MuZVkO+xUs5vQD5cm1WhdYQ42H
W1WETpTbnG/tpnTJ8I0thr9vndmB/AgnjlC/TB7IFbvozio8nMhJISLhIC1CV6tn
OkLcWeCj9D1qjcWDPNc7zzLtyR5OHroYM7xBwH0ZU6U/dLyaL1IRPAjFk6kxldHx
9IGBSZVZ19c32milKApBCW1kAtHTCIBgJuq9utokD3oB1ib1wDJ10davNH/Dp8bn
xM3chBRGz0ZvdDZlWzANiFIF//JIDXwj4Zez1c8l7mSsh06d4ryOuErdF9CCYNWD
+DPQ3bInrTrMTWqfhUlTP6DeYwjWFzFaSUpfY/zhZ/LUR+3fOORhjYKXJ0XThNEt
hoBfegTjADgIrerrBTKGDUMRStd5JTo3lMOBzCvUOO1N8E2HdIzPN11KwMpEFDvx
NvnkPor95yNxv35JJYpkCHyV71cm+7YuKzxcVc2XJ09jfV2dzUGcuW5Macj914IB
NEBvHXrVx4QOBfQA401FVKJuo4OgrlzNlU3dOAxplEvragAnKhQJBL3Zkpr6fYAw
4mtDn46hHF0svNe+OLOhy+jCJNoM0yPXPN7o4y0kGK5myLA13tyHEUGCzTk4fLxt
p4Mh9b6fTPhYoBtWUmROWWvKgxUfUelfGe7sDTMhirHDuO1eDCQ4E3hmj8CXfeRP
yRH+JEK71rpNdqJb8fKsQQOX5VQ71yXrC8aJh5c4LWLeeL9FUyFvpD7uU2S1bNjZ
taqhcjNBTFae4+1uvcB1IkVcM6NvNjKFfvwK35U0g+pZZ5szGUsj+15H/ZtudZ0J
SRMqYgMWLZ2P2ZdHeBTc8AgV4VhGhAZjtAUDK2QCux2TAo6Ob19C9lWfAk3ilg6N
X8SQcHjdUOj+ZqnPATsxDREAJWtscZ14pZLX2YJFWDz15ddnfhe6Piycz1dZlh1F
C4z4EupqTX/YP2a5/Qnrn0ICJx2VDiF2uKYxhGw8dRH5OIldPzpgnrmJjc1DRcj7
kGGz31ifEY3rVLyca214N93/v6LDvc3tLnXq5FfnNUSURgWfecdHle+E2GKW8P/w
t1dl0QbNWYWnlYpPpOiC2kvNNiNAgNcq/KOnuEq9Mkyk32gqxGh091AzEIKjcbFY
OOzZtLahNe0vGv02i4w+FJghinSBUNZrxduNVnvXnKxGQ0EVzjN6GQBLW3W7YJ80
OzSFXk8AduhywYjnGy9DlzjQB2MQzrJmcd7S9ASWOKBnO5CKWFHD38skzleMhsVa
7ED1g3o2ZNkzy+VZvmuM3URaqwBa+A+41SpGkTBrGmSMs/r6Ef/HbmSNq3CY2Mv7
ZMsescRDaR4d023wwCQlP4FFjTdsPkAzzvqu/hDiucDLrKpCmAtZQLWuRH1A5rLQ
3WQbBwHoFW1QWig8Lmq1FE2MOwyP9tbTnucR1l76Q92IMDDYahTvcr9xQoQeYEvf
I28Y2dY4g/KVQgwADwuVHTaKBEJbDro0uVYeMd7DaacGUqWCaK7siKhIwYb3RVkB
0+j6h1d0rBXjbtDQotN4vG0hzafLS8OwxhWi7ds5/QEStyu8bsEBPq4FLoIRaKt4
odox2Eii082SNnvbBh7iWTPueMy17trTYh07tYYImdODrfuHoWZI5HNBmhAD+LHQ
GQn2IFRH1mxa0uuG3oZZ2YX6qytMEnK0f2S4tm4rN6gOwFAJGLWo+6AvNasctGdw
/Ar1QsycESizVZmjBxJM0Io/TZor8IXR1QewmPaLr5uWWenexwVWxgqSwkCNCiou
I0/+PzBiBii4/bqOGkC4EMrrgAc0IaXtzXHFb8LJUvubDOqSKkIx7fiaejyisqkN
z20d1aNlqWioEJ70aFoJ2N8txtQWLVBu9p2n6w+QTkMXrhY+eNr9QTcvqGT4pjKk
E03gyL6WKPzyKu8cBvcd9mw5AaTqycpyWplaxmQPpW1qiTsJ6G9etWv+lD/0yzAp
YNbCD+a4xgrhmx6GjqyhIyplTCQANsXcZDjgRmSSEvlA6RKH3y3VFj3Qhbx3rpTq
YWObjg/qKQ1RDftH68lvMBZbDEjFr2MeoaOv4/et8Lf3z7CNv1yQmb2mzwXBUVUG
uJLqdjkXEZCbxonAj9JsAGp9WY+ZseP1/hqDiFTKD1KNu5d+20QoB5SfRiAynX/W
CPNvK6ykG2voiY6Nf9AcBIFHHxhAI+A9VRVs2RA5pcqE7WRepsOVv3ByU4mLqSua
qkuRrwVdusuKlMeiRl6/rPzuCMeE/BbJhGI1hBF4ianxhAwE44EaQxAfQKYv+Wf1
iDgM9z1lm2Jg5+qAMNrqyNOmnYOezGhcnLZwha58vP8tJBHUXFCtgQhqDcx0x2i4
Yd8gSg3zJTLxUPIDKO2wDSTRskIYdysbeqtp0M3sKuNLFzawAX9V563FKRoLdyr0
QhLtNgiaZN2UDEs0i3iiJAGkE1kQesUNg4A3eWdlJTGRw+NklFCX+x85j6PhKio9
0N5RF2T2DJYc/8fghyochDcmqdGb1W08NN9k2ZstkNpgVzYcFHXIgzs0bW8BpVH+
oTJV4p9rthpftDm1zq9Wzv1LCLPqqGJ6d2z///gK5kTd0gCHP5V9DASeOVfv2mcd
OW1rllCqJXGFnkEO17pSNbYR93SMNY0rErJKs5JkKXwEIYC1i9n6FIo6HvzUvQdA
8J5QINmc+vKB8KMsybme6fHw5VgEA2uhuV4Cv9KUE/1vK+CwA5v/Jznb2Ra2V/gg
UkQo5M4JW06k5eZ7ov3qwU9vFq+Sdz7P2LGit3OLk0646FvUKaS7QyhWpEtePdar
97DnDpt8BsatPmiHUuk2VaeXqVp85C8gwmPisd3OIDb2DkovW2c8kBJCHbRMY/cy
B7NG+3jqRaGoY/xH4BdFy+ESTIJR7pQ3DwtTYzGdNtCGkrm5fKrQ4X9N2uP3aG9r
vN8d8r134q/fj3lGq6xPxlQSLTztrOLOYx1Iuq2suynm7S4A1uvuoYLgjGG7UQGi
Ytpasg7G+GNAUPJVisS8RA8OVlOEZUyvGVwEU3N12pQJ62BqRe28rlc+HK83ePtX
tcS690msHsdqIkAMUfsHnsvVOuslMGY/AEsiI9arMOdwLJbxwQMb9ILzTINKxN1Q
W7B4C8cMI8EufvqiqOfhp3Z9kR6pKWwyLZyeAPdNpvZ/T/Ll6hkGVHGr4SGENEnZ
V2ghYc5s6+ueEaqke/CuRhmTl7XPaohz6gAdIUj78sKZ8m0eL801520n9DluMneU
54E+GCCYl085G16vPvlqxbQmxXMHgKUpCWqWs1S+a1KYGIh956Zd3xoqboyRinfZ
kqvOxnYGCZxbiMCvos8D5PgRYV5I/NJJ3qTjb+nDf55t7AHpHpv162TpT53xyNJU
gssZPquxnQ9xVUHRNSqB3e15qcyTooneEmFt8MCefOBPTispLcX56gZvgc/FjXjI
S0mIDpbcTJonBVWls1oJJdXuKPyJjpHhQXsqc1px5U78qNNvJhwuMqvqjHrQkqTk
qWdZCKbKhbbqr768AUtng2FviO0pZXIcTIKfa+BkRaOxs53SKQWQwecvq/5HhgGM
46Xp/pVMDwW4Zn/o8Zxcpa5a1d3uLsB+wqnL0hsGsi5HCKQ4u6nm1ml/DBdYTjtj
aFjHK9+Pa24t5Q396H5e3kjSUE1vi1UrL8gmBu+cW2+ifDWAz6qEHJc27imosGmb
eryHDojdeEocNro+Mv6rSPpJdtHUYA/wIiQeKkj7K1IO+GloUmKF+gRKkTjmikoo
XUXtx9Bkr8RdJ1Bcsx6OfoUXLco3GHC98Pue6e4DUFm8GiRTjIIqfbYpqj9/cJEL
smGLflB1cZS1i/LSUU37Jiu26Gxu3hZ/Uhm/UxAQERIVdXi29Nfg+qXxS5gOpHQ8
S3XollljRwtAEYnS27XGDlLlegbKohuCBs71QBmY1PuejdiHus/waVTMSgqDSN1C
0EufWDl07U499BuTIK2n5LjM00ELgDtiJgyoRodPegjTQNHAWNixDW7pR4ffRfYn
2xbIVB/y1gb1p8W39eESBV7Z+scDRVav3t2ArqCU7u6lNjikl0/N5ciyMS+XVi18
Gsn01+F58ql+tNhcgRdYhnsAnK0AE5G/ENqF0Dbngw46ezihlTGcXMVXYnTkFDEE
FFQ7d7WsJXfV08I6GjqooXOFZd4K1+Xg1Yf/pULZI2qNyIkJmcshQcocZHaIPew3
qQjOkWxDSTcpBW9p0d7X2Q8Em40d7ZhWL3lIq9KL0REVxohX63vcYxuK+Je9Yotq
U0LFtvn/kqm/YcV5t6XPfzQZNWEBBLzTC4/oQUqsVVApM2t2Ybth3WVHvfHMcvWE
wJIxWQqzWMOC78qhA2+Gv9k2rN3bdNt6C9I+IjqOS+n0bsScoXjudgeh0Gk44siP
c/B4g4cKotDCHhkMm2SwCbt980WxNrYQDSh9LKidMRc7A2jeHqvxv8e9R3BngTZE
Jg/4sSikyxFJyEZolOpoNqY2kDoGdexjTBpkcJInp4b+wq1YkrFmIgrRnW4R6fDB
HcUK2X7Itnyt7BgOQXvZiYpcbN1/GP8f9Y9yTh0I7IcJaxgLb9B6bR/GKAj92i9R
a4hbrTG60wBNiw23HAu29Noi7e/3kuuTh5FDobBh8MFnuV9UNyULQ74gHENJcaQY
BO1FDHeX8k1RN94QqHJRBAWn9aOTdpZzO7RPWeFNEKSGC8pTiodaUamWsOME09co
HeqOtm2ya91YRZfYjWVmEguhH+lie+1pjETuUlZhr9evmiiB68tC7DhXlNiEILYz
Jw6d8NQxPgAvR3qpWhGokRalqBCbKzDXpOqE2Kc++GRmK7SVgY3LlzhxXXSzd3Sy
V79b+nwR8OaEpjTdZlzvWa07FhKjNZIc4bfGCfWYvoWBwODFcaAAqkx4x82/vGFR
Cx+qMKaXrjASlAj7DcePbl7NcmeksCvc0pWJey7ttzjjo0h8KeYmBXoOhsq31GNX
IbzDvVOW7uC2rho98OQNObjlk94HRwdrTWsdobtP+mVPLdqRp4eFJMJOpCmYdh6K
uT8VSPMsvvJ5zE7TZf0Wsz+1H2IxK8zFAulT7A49Cn8C6F8Q8ySRk4/Z3+xgLN3P
oqJupdSWyv0VqKKZ1jeXLjvrMDwNDY6V80pBSLqNMQfi9jw3KAx8WaaGwk2pZ32O
Qxn5Djg63U0GYJ8OC35K171d9USgEq9CxUMFky81QRiFy4VaWKkTx7j3quD4vhN3
LgXetthSAOQEMoYIxds0bQF93VlMNO3n/a7otF7LJQYHy4lJvFcQUX3fc3NGJT9L
at1xGiEKHRU0GOYGv+KvuGFxbPV5SSJMxb3SXhvC7n02BZ4NmE8fCuddVKIiN5Ad
mRnmozzvTME1yqLW/2/vnxIbSTMZ1zMdAzg8CIwhSllog3KrPi1zVYFrZFSsfk8J
LFNW3B+v8ZmDM/PtBHLo950Dh/kRaE14lrxvYMTL+vHvvY9pbc4m+IjLeztmN/gH
7txqxraEhYgBmpwqkmCs4gT+7+ibWKeyjucsB8J4v7N1BDnfo3Q234ihga9npJyw
2miW9lUzTOlt9lKXxtZ/pV/iny8ix/uJ8rPST/p6+7Y/vIzn29APa5b2kWiTOcT0
Fyff1zL4BGp839+COa5r6xk7G2H8ByNAxn05zMa4C880Isyw52bmHx/5cfVIhM/o
8p8TR3+fcJJNfteCmzb2yuG5OTI7eJKe2krcaP/VCOOITsMFfzJwnXBTSW2qPmHe
ZaKeu8MmHWw3WfFNDuOo0YMvA5XYwK2INj1of5Kwnzw0L3q/Tt7j4c7DYxR2acdL
+WI4QsujlXUqptkExqZQmrsIYe/4FA7BnUvlPpsfIhT3gqYvjsrmvgp0xxRvRSSO
8J044gfh3u07bIRniiwKaGgX7P5oHwGCqBSVKxp0BlKhvhnjkbOeRNyN6OwL9T4l
4qZKCjgo/miagBSFcP3s2siiv5CaN9BhBWcqJNSugnZymY76Bq0i1lFx0fDZeysW
M+gB/VkEhMjkF6nn4DpcP4hEdnHTQnhLhyya6Wh1KYfTXGZbdxj9kIcE8tFtdCx7
aLgJmELdROz6hwdtPsTeI9xAEVXH35saQ+LsawDEqeJvqh8GjysXNLOZ8eYvQTG5
oQ+BEMvXF9Duv7qR0jmJml273aFptraiIQ8Aw28d/7I3JZ+bQqnoKvF0jWqWpoJG
wsV6GGZgMoHbfnZPjLgOb0iR6MnsDzwSoWGimKYg7x6vYmW0Jma4YM2Ujq7QH//N
ppctOJljlFgSKe0uqKhpFtoY6NxDGUYiEQ3HtanTpwYEqHRY2Fxx6ZYqXObOtW0r
7F1BDqX+DjTDG3rqOP0OJtlkSqHYGClc/ylsaFVebRGouwGREIm4M7gAcZjOUwH/
pQOvqwhI/KI3QazkCx/LchnkswzkBsdlJd0i30evSp643qsFsjUo9+7ub6IH6Wvh
2m8dPkOgSaPDs95JQTZTBSWjD/JuXe6/M/mRLh9y1oQyIsgHrc4oBO4fNFj/OnGp
/uLTTcYUptfnSdCCZJ9wfk8oWD9pCcup/+mksX0zlW9beK5WGNcromXf5LMcpZ1P
P/7u6qtJ6sUxlAAmt9r/G4dJe2SWLi//Jz+rSQdaXa+/GrF1q3KeMLQCVFQ/0vow
4yfykavffyz1xFXOLFZ/IsC5M9Ri99AcNMNA7jTMU29QOx8rzTVi+nU3O+0gGW34
08gCSngF/fXJ66gjseFZ7PmitYTti2w5ssR2V2vAUl/zPmsVcaVgt5bGviNo9bpM
5MJivWo9qjc9yh8m8RQxBh7ycMIc5txcjPHpMY+W9FpusEBT6aARtWRg18Cdgu8P
8jBBkZ6SO3v4CczyGdcMJtv5Lkyle7NUYTcp/jM4Juu32aT3WMXqEkHlkpvLre3E
4aMTEB2WKkpPWUXK7TeugI0SjpGJh8xPt8sjNPPuRNqZHT4BA5mhwQFLbOPdwtCk
RskNCPePiHgJTxzUT5GYkZVQy58Oe0ITHd9ScwbWO5sHXd+UnLrzKLe6KzhtJ3ds
DqFBAO/PmaG9KguiHkpN7UAtRtLwJUo+/xHN5NBlTcu1iEDd9Sc7Ini+Tz03EbzI
HRgN97WX2gzTWXZyYE2NLFlx7QH5llzSR/989AQUUJw3WloYFXkYr2s5Aj15ZOcr
Eo1Sj16sv9nYqvJokL9/RNOKWrAqMibgme3p7q2a3bu/3uqm4E7Xa4mMbr2ZjkG3
A5HF2YbZOtEjx0R0T+U3ezMSF3nVpOIQQghwcrZF0s6p8debKHwu4Mh/oxlLQY7q
n/wcvWbJqWF1EL5aV1Yw6ZrMpuNJw9Qui4QZbmxvDzQkdrGyDUuHois8W7X1wKUV
kFe4tVtgkcwcXXdNwNql/OWsuqV5VxI8tqs+ONN3Ae4llGJ5r1byGdzKgfkPX0Bj
jaq5LZBlaOqkM3LVC/mMRTIB3snypafdRudtAUmzd9YdxihGiKDxHp2dVueGDAqF
04sbPO3vyPLfDIAJ1lFgiuauQ0uR2+L+yILWr0Uuh2gd8H9wmLxK8KnYxMOTzdg+
Kd8hFYp0Gf0KOSYre951Yf+Jx0hAwCAu3/DNyQ8hx7HeCIU5Dhcki1IsSxI0zwYK
eakCJD/KJ4ThyUHCi+bIPbTcr88VoR87XsOdmliR7NdhhSBcHgKlqFqqZSic8Ulu
fkA1J3Bi9UVa7j5sQ9lL/deF+SAoMKWRBaaMiMb2ktDPKQoKk6FIlLuPx0Q2dwjW
EhbDkI4jzaATRcHk56P91KiRd0dsdq6ieW8wxcuD8wGawdUpzY5w5jn9hXwG09km
bTFDZdwtt+802nHnSneYumm/T8vrg7kHrPVa6SU7UxEQU8ViK9q1FCRj8fT0339d
As2NNrMf1e0sQdLGSgg7DFcGGszRXF9p8cCTNhhxfOXu8FEl3dpwzmPFcB4Cvlnk
lU3SX6sCrMR5AwIjnE/CHfXVQyuhnlbuchAzTcGCl95Ew80N4qE4eSXVV+IkFupK
11E11AgoztRZXqh5x8VuG8guHt8rsRAki3tJXr3n5lp1T2aiFSDQkWYi90SPayEy
MhvvB3stkXjUjnt/Op60lbGrYKT3H1rUtFkkuweDc1WuAdrYztYUcMW69NOoURZ4
k1Xo/09PCmDGu1FbxYF8mDFH28kEPje7YxCRhB1DihtFNbNsSkTmO6hteDuKRcL5
OWlC8hVbgEsn73V79oxkJC3UMWdlcyfSxWYFBwYGlHmMKfqHjATJW7LWaE5G2n0z
DeBtVHz1SHlAqELUGLfVnrZQjq05xrg9GSDbiSEdWHmiyOWJ0pp6aAyd6tjjTvnu
dhrY/V0CJlsbk3CvcoRxbhHxWGjbl2n4z8iDdK3SisTcdFRT0uQ4laBgqSz8bq/Z
rPK5//zkuXOVIzWZIiZs6WP2tq5vqpgQrttju0D9vNF+UF9ZSXx8a2XAbTIUDoh7
KsJJOYplydvkdptHEuTSCjQUdxU+gNJ+1JB6z5uh4+axWLaDqAWytVLpU3qR4CHf
7yeJkaNepjlod6quZ7xWQA3mcPcQBg7+hjDMAcRC6ciV8T6520qTDBzXRN9Z35oM
YOXCUWa/+Fy2kpty9EpuIH31ZbqOEEbr1bfpNGaNCnDGQXljfuTCOavWGjFd83dI
8Rwg/bQcu7RPVEDQ/NWWzhGWrFhyzCEDyNlaz46IEXg7oUsQhARseitJmtZSGktp
ov5ZNHGNnK1H/hPT6kTyfJ8vppMMI6pLtwU7Gj/IcydTNhIx6Nu/t+LlLxzjojlC
XJvPkHuZcHl86h4P7xKNmDPMEffYCSMI5NaFuXKkTyLtMnJFGUpzPInV7Ru4pR4U
a41I71BziMzUdp06kswqID3afNj4jp9Fe8nmOKQY3WxcRihAyZZccGeRlTcEmV4s
YZQ0FnZiqxy/Ne+VB5iqjfkqZGVPTrk8tf8b/P5pPZncLVc72PtCGDP5oQjhsaR+
zoOD1Y0DtKRX/dV4Pcm3uWZHTT7ufs2l6lraNkc7ow6C0bxi/AzNEnRvNvdGjObX
Q9A2XzPjP0A6VUnZQjcqTr4Sbm1khrf3CteNDAzyoqhQRwZh2vY48o50uPSCCyca
NFzwuz+zVgPCtSqAan/wyPYXI3YE3WWYqVpGLzm2Ih2URNAbzrFOCGdThSkYGoA1
8c8yK0fMkEbmCAxxTzEvah8pIQV9Oz2Uz7YDQ7dWUkXlXlsEyESRA82S+v8sZcb6
2o4IQ0r82VA4f3gneBx0x/pL1BA/YVmv2RkTe1blqK8NgtrcO0uPLdMuZr1XT/Gz
ajPNFSZj/CmJV/AfmioYIQi7YhYKMqq1jlV+3dJEKZ2LSIJLWPS6x4aYF5areUOh
hkcjpV3FVVUyjsR5tT79b8z0Kpb1ak62GIq8OQLPKfpz8yaAnGRS8SHa4cDhAPNB
/qSc+Wi29mkGKbJCjoGsdB1iX5E+mUTh95ioZFHNrbXkwoCVhoG4qPOTJEyAVSg5
pwpw21CrYI3zMe9POsv/zZVTwsnsxdpMCctQa+y1QgsGO4o5ICEKpcuLdpQQFETH
cIXl6TViOdneYAF2VX5nrsKwQfkgpm1N3U/NVCdharVcoc05ZU9pyAoVRVs1/SQD
uqkzsLKuFJ8/oXkMcPhqnlVsZHeIqQ9wzZg2c9q6K8+z/lpb1m3MdykD0hWINmLX
7u2vxv9hzJ0sco+QOACCOijbuei1d3XfAiYezQWOdVTWIjVzfFNeKL2zBJYEqPni
+rHupZmQuRRkIkQkVG5e2QADJhvFqPZXNoTTxgkNwmbtQT9jXJviTSoQ6NStWVwD
3TmGi7rC12ztKVvovUBkVDID7FEKs3hQi9crRnBnojUxm/iZcOsXSbX8JrsKXcEI
dE1+PPKZ9FCjcrUnynYn6ATKE4gvSfVPXpgR9BxQX/hG3p/9H9wKa3jLNKmD5aZP
3pmjc1KlVTAraUBjGoZBajpE6gSFaU6Gj5/u/9klL8g887YbMNA07Odya8qE2eR+
AlGwm55xwhPG4it0Kh3bbhwy1grwFp7zTFcFZE5qxbPF+BAjatwsfdZ43rsuRz41
D33TmYFoPHI5FGLhfkJEy45NhFjEWzJrBnoTswVCDSB4Ft0mKsA/4LcyFj8BdKl8
nBFMbPS0Szk03s9+RYjZiNQwTKvZfVd8VMOYyiue7jxp3IHdJqAVR9+GPijxczdN
4mo1yOKY7ZwkE62A/Ai1uBbpdQ/5lYuiDEOQA47e+MtlLUQgIcHdYjgro+bZ9n1O
LQdH9WE604DTM/1+uVJA2QF8rjllDzsZJJ3NJGsgP+mO/giIH8upX8Bu93kiyjy2
71bGZDR1DYbPTzpsv/oH4Fy9z8x+eayOIjRsHRaJS4uru4bQWY1BDIDAleSCg/wN
ulGXNJMybKtBB6UunroWekjNl7yG7mZmZ9vUtODPEzMK+hIOf99CHTYI7kjPNhfb
q7dWpI0s+jpkz5c26OAvhyoD+qG3BDqPMSNU207z36/19EwasWsymYSoR3gse/Ol
Hilt0s6V7lYupNz7UGshPXKcHTt9Gorj3BDHFPVlTEfAZSM2G/mfyUEY2Jzd/ueg
P4loNHQ2k4LozAF7poasIrAgIVICRf92H5P9QhpjaeNsZLKZUa7Kvm4ywtKRK657
4o8zc68S9zCMidE0tb2AHOdSrEC1+AN76tph5NX6016PR7hyK19/yUuHQ1mL633T
Snntb/B0oq5yFpeRd/bQzQNJlHIH32C5LJyNqAQRa4fjza+bYEYnGHcXi/9MkIdO
Y8+nEbpm6GXMTArm0G1an+OPNqXQ6c63GSswZp/vOnshMHYYWhdjPREe7hMEvj1t
wqEsomCbTj7WVHHQVdqlYL4/irFf4HT/TNjQNREKE+mkKv2SheUvhaKmmCgr1xBu
IrF/BhWhYmrTLBf5WJA73RWc3dS/E/Xy/CsjcfFGfV0Ogiw9nTRwKRqDGdyg/YPW
p6EKKBPWVCnyBJAw1ebLRuNSzdpK+UH4EmXdGJY6kB6T/GDslI9PgJgiGrcr1E7s
pHTiJ8GDyHsmJAnufd4mewk0K3n3WV6h4DiCNToSllkLdYDRFyBwBxcEIgeH8Mk9
N4WkDF3DWdMczuuUhWq6g4Z6EoWCs9FrtnrHHCMGLXtj5Cx8PnBEYQN1j5tN1FIU
5LnbqvjyqwDmFwj1Kg13SSWLaVkCnC6Zeyc0tJJ8LQ6uJRUmgVzVDThmNZG8uY09
D9c5yoeRKLvo5bUv60ud20SoIZNo7HNqUfgF1uXOtGS3LNntN3GzlIS6NIf1OZ5o
xpaxu7M3vERtI0pPYBwaKWcMzlrq7s2k1F/tQfR+DgeYJMdtDEqNle2RiFzkpY+H
Ici9KKRB03HhBTZZvuNBHvvU5b5nUBMHjA+41GZZjTCbBbt1oM11dxtMqgvtBBHh
AfLo3zYaLusZm9dSIl3FizJHDhe2eoiFDoQ7iNmo8d5nVJ58ANJnezJbqDKINVYi
8cmrZKopfqfz+VCObZBRyKCNHB3du+FtJDtIMaAchiPGJDHGdVq2USqi7D5FzIaA
GKOwmrGB3p3PCV6DXQP2ycjwxfReABzOoi3cEVevsLgm9eYLeVNAL3qE3BrRknjZ
ApaGRkuI3B++peBWIM12sgprefuMjbcx4Zequ5jA7R45f/OyKyAt16/6nhRWI4sY
WH3witiIs5lEmiTGNRi+Tyi1cQD+dNaUmGf6AC4ARMRW9JYofxgNhYFby7q3OheT
ztMBkeIgbLJzlzSircmC2492cwJi80OWJcVuXUck/1PuJ4rPtAZi5vCcQBmhFld6
2rMGG0D1JAFymvd/BXmLm30W9I7f4ppa7RIpib1k39+0tQJGUzvzTD8X1jCO3CG5
5Vi9lXP9azqG2zIUxnkXBmNvtY7tixr6DHCpt0fE5NVOaVRekvue75H4GgMzG8Iu
rI26aFoOCHHalzvLPAMBwizuDHIgIRQ1gX+gySA+2ahKuvN9S9t5mCnOVCF8bLW1
VtLCGfgCuOTXaY1PYqOPODkNUhf6AT4mE4Q2HeeEnfD/y8x6QsKiMP5Yy1FgP5lL
WvzNgqmkBPbOgOxhCTeyPxEB45fKPsQo9p+mn5A50JbqnvpG1i20cLSI48ub3DPA
1Xi2zY0Ef1XNh/DsGcioR97qM7QGbo2xDNmPKUxjvr2nH4XnJOwSx+CnXq5i+rA3
paBitHqHUzzhMF/MTih53Vgn6zVi7Iyupe7WHgPGPwhcaLTMTWef4g/z7bomvfBB
TTM4aRmHQwLvWUvAdqOs/ulagRSDrM9qGEHNmyUJ+MgHoakOel1FM2b33ICuumj8
X2oY3s+J6vgcLz1f+yD5yJ0FXpt+i3FtusGYM6h3PcBo4O1gpd33/j48IkD830DU
4In/XieFFpGBsdxbfjJxdLg6bIKNFq5VGf/6AWg4cmQe91wd3UZd0MzK/QDvfYnh
Mu1Rixxhx5syqYDs0EjA5Cks/eChfpBzX9EabF5BTdCjKvVyN9vILcOYvHTpAJ1n
oJUjjU7/wtT8fcLeps5kCtsuNV54SfTSYBmW/SyX0VjoOHfF0Y7Bt9ifXikTkV0O
+RnxD8UnWn3gUcIDX3O00IRbJI/K8stddbjiqip/iYlW4zZNlZ601fAGe2C3S+Ul
bTGnDwT24tAmdSsM6QyJX6Y8bQH1T1XyYlQiFFqoaLTe02UHWqgy2nWAjSumMLVz
LEF9QVoKJa3502YMYFc/5YZnzEu3B4S1nH1IiZOdVqFl4Ntt0uXRyEku2xbdLUsK
KDZypsNCkM2BMNiV/tlNRKjmt3g+SZCcT31+XYHtRMKpKxnmA6tG2ZMvmNE5dZYG
yg6xs0oYH0cpiFTaYFvKUVfBdWzJKHZlRzJafdn117ARGp84QfcHjbAJ2kUVy8sM
BlF/oDyY9vdJcrx77q+sM4mr0jVkQIDta5ApYOfGRxOox5xPf58vwFY/0pdY0djd
hPlfIeZ6/Yf3xY3vDWV3HTGPTIWnfc7QG3sKFq1NrXTkJhCO6SU4ymru/XjyuHYJ
AQVxKpCNkItqoEq8ZosPWrFMW3HBuAeXylrDAAYleMDjGIIRLVnZmVj67SIOCELa
hhQc9wD0eQxxgE0Yn8eUXYqnPCS/IFuWBBUaaZM/V6vDEdGOdM7Gs5hXL/e5n4jB
YdC4gHEpjcasvp+MAnmnmN7Cu6X3qKhMl0o1l2BqutkPHKLxt10bkJh3LBvV8MHJ
4/EOpAgIIf6Lu7sVC1wUnOegfkkWSLoQKJNZKeFLU+GC38XOgwWYLA8zwdADInNO
r7AdIHXE8nSc09cpGLMlIpzwHZOhWD6IeBJK6Z8bz/19QzJjkkfTQOhNWIEJf8SP
krGUOkPsV3QAn2L4FnprOuLzp4nEyKVwQoSIph/A0CEJXYEDOufL+9VazL8foqPQ
Dm7j4BtZOuzl3dnZgMRycNmsWHnTFg/bRXprbX5NYDSvhG90ZBlu5gknQz57WHKW
Ow5RyrR5tTE/PE/HnZgVQ0CJRb+psiqY5PRQGtV2K/0JUHCxCeCSGMRf4aTuUOVl
zWIZTGXL14EhO8CapmiryNgciudcQjC1HUqJdZCmPPXtq1aWtRS33GmGdf7c8dvK
KYHPaAIy7kKiLfTOb5PT9qFDUdxyuVYXL49uZLgH14030Fxo/EwgdnEOmhwm4AqP
su5EaGpInzIxzJ2tSx95YGFNW9tEr8BqetPurNWInd3+LFg1g5XpPggrDAPjbExA
9Rn/W88/WXn/kBKkTYDG2BzZ4SfhymwJ6WGiS9V0EmIsem0JvquoX4e9dpc0h+zq
BcBfUnQV6LUF0wLQDHd7CxIrD6G4VGRlxGZfhttEWgghHxBnvaSTu1kc1c+cm67z
OQTIGwb7wfTlQGZHjueSH/JHrMY9SLHajcvWHQ/ZFg3BRxnpAHO01pSpqj1lZjMO
JT82wUCHubJtcp9fCYTtopF+KhD+wqo3gfWTeUJSBVFuwd2Qa6skJT0G+Xn4HOiC
FO9e8BlVpneoyiG+/PVqlr0WcsWVIS3jGDP5UqxpB9kZSTxoAR7KUsTfyFuachGD
ME0/yGK8n2VTmuLbhyOA2+LjFoETvl27Iw5j4MQB8rHxUrEoySa1xE5xvRpF0ctz
nmGj1RJv1yRLH6VU0b6t0szwhcCoTPb6KTet9u/SV1mqP+J8e+zUznIicake5P75
ewcFVXcQv0EkvjWMw3I6fBa8E+jqDRHWAUnntm2CFiEvmNRzzZGFsU8l7R7gkPDU
+ITk+ubHd32WeSQL5ysjVkOyuLyI8SiCB/IiMePzj1uaaBIvsMH0cWTHd0Uv3q15
rrv/8FunhVJ/J9wG6TBcWrpK1i7M159CbryuAgimrGQ6UqzXx+r8INupQS31PNss
Dcrbx/Cld72NQKUwQxO1Joz7yZpsYxUZW46DKLF6F+QJH6NfOmZZDJ45k39naQdT
jZZ7W+tex5G6NFiF7123F2pVIz82l+XPsE9QdRHCwfefxm3XFFvn4L15HFCBNkCq
7U/2+g0OpAqVvShsxbP+DMDjVI1BOtyc6PX3WXEfJZH62o0HYerRrjiw+dJS58fS
dWt7xW7pdPf8Sh6OwII7uMWfxj7pr8o9WxtJ07Ld61BPW9dNppW0TbFgrRvtiwyA
lFoJFhw4seD/mQYyyK7dMjHBmgLbxfYV8R9dfHULLoRlEsoJAGs6WnUBPrgmDUnj
m9wlHqxEftm2WuZFS+69zjKuKrCMkww2GOz8iPDuO2/OdClJDp6uzG/t9kJNqsHt
Bsv3EMEqabr0u3J2ENBLNT0qo7TZHpmthN4n42GLEt/wbpttgCG0DRTDaqcHNRWV
MxTYRm4Gj3Tr1lWRX5rk3/EpSzDYes1lins76Y+JJjxvX8FKVMlf0p5CvZVMneCq
+A2VCv6oLyT32ffHrcLCT4sPwCtNRhyp93T+kt4Z0ZAqqQP7itnRWwZDj7m0TSq0
X0FfZHg19ttfodiS1KRIYPNBv1tFN69rVazClhpN1Y7fD7ojrim+nFiyK6iwtE+M
uShPDqfaP/vcZpDt0bPClyDTCgLPzhSb4mU0025MDaj4hi3p5xGtlQzE2rI8gYUD
BdruWp/dipx/3X+fojQetQSJad4XSbf3j30Y6EEHuJTljo1PABIOE9BmenD4Fbod
JQt2yCIW1xW+UwGTxicuohPs0fqFuwqQlRhl7T2BMqKoJs2PER0dNWK9TX7yrHn+
DgjtRU3WjJK4nBrOUawaZy0QnE73vFXs/xMFfaPeBKuGIhFpUTJBUK7Pd1VZRHUl
ZmAK99DkSrnxw1asAseUlyDhwp5JrFLLTFNECzM6YLBommOA1uPwEKfJunxhAvc8
sWc54OXXt8BGL06vOxhJ2NNXlunrJys1lvtLtWWrAyrv4XxGIYSI1lSdgPC00l8K
R2GqOkrDIHi210QPNHV5THPyp2prQeCu9Vfq8aQu2/fd8+fYtiU1CrAIGnju9OQv
2J459PAPLFE6VkILwjvoDEfh3XnCt9NbpnKQf6E8ikVgZg9eyfFRTicV4PofrqzJ
Xrh6ov19qdAvgrNybAXn/7dsw+FMgzU2gM4eBAV12bIdUvKF8ALI2oUYWNFoNwEx
PJ3TUfzxHDSD1gjQJoNsltQeScDcMlXh8K3tTQhv+kXYfQkQ1X7hy9MQDGs19VIl
rTnUpwb5xDeyirkRwgICj6p5jX2XZqeF75ugotQHxqD333Ja16V3063NqYJ8Yasg
pNZPIbilEibobco52+TBVIJeD6+7nDOCctZYHj7rbfF7n8bKEbgeEUrwUTWMtDFU
34KRpFA+plNpTQB4y0ngCbuL+AQ7IQdxwksZnVhncFqwQ4iTxNZpCgzBMS6Y/BYU
oLMJaoiqozFedTzKBfKozvrlu206w4Fmjt7qe55cMKEKfBzcbGDGNdL0DRBi/2KO
xT6kIMBMYvyXSPqdZYGCITsWdIYb/1pRWVR0dEHrRi6baGUUu62UKh+uvtsqFyd/
KsgEHKmGniXPXfNeYFVDBSWOjciW+3DAvg1qGQ6++uz/DgY6X5iJrDGEdBaw1H9g
d4GRp1MpJHDmx+defFINrRT3RTpZwrEwqxPZZjfNZIz0PJ1Ggow7qRXztoHjFOXV
YrkNqAKxhnqVNlYZbQ9b3YWJ1Ko3JXumkGFbQnxpWNUMuShl6Q9wpD0LroXAvloQ
A4K9i4aGMssH3jEW1Rl1hsTHIaIAK+7IA3mXEiZU0kie6WHX6WFD/MnDGHIkVz5X
AlFa6xM1YtXNKX9Hr50WCFa7kYdwtobuc6job71F8NN5tK6LQJTWdXeGfnfeA/g0
WY5Q+YsZK9bn3dPm6phzjWfVZ5ovQ0Tw10OxY4O7hXJkm3jlftTxH8VGANowpBCi
jvnExxFQcSrk6MA+XlOHPWsxrDICIIeWIe60zRBV8e+fZ1XklkauCszi8E2gonBZ
9DH01KevmvEtgiszGjdDlCvmeLxHBDu7yY/faXY2pvPnBOq7Dq46QtfVy6ZHdZN6
7LwFF6en03JWRI9eDI/hQ9b4kuAdxlVpFhr2XX3b/VieuodXEr/1zjleLC91smIQ
PWMpZPl3shFkH56RrsC+XnoXKcAKyFqLaPp7MYJMoqwly0s+QW2jopc/6rkuNPdQ
WjRCigCpcDGB6eJkfP5gdWlZk3z/UdlYltgoTjm/7X+xacrRKIotCKyhaEZF8cgd
zHb1GHi668kM4CANVIfxV1sI5KLtFmIb1Xf22fW77gRm/R5cMiBQL+0AFrjlswns
UUOlRZ6eMCOhfuQdkDoH4tusQRNVFMyW7iVsBc0+/vzeI023GqwkKMmahTI1IERN
XS4E44FpQzfRvwgf5XWWkaHD4ki39Kbosjhoyr16U50o6RbbhjFh2X1jB7xCe5As
k/WtciTHje0PjXL7TKIKNWeMUq+fbUtzSwV82SEoPzWSN9e07cPMzeAkdp2OA1+i
qMeG8OFPxc30kUdC8GhXM37ufCg35lv1bmHbL0xZ3gxspM8/AQCHzSTPMlav0wqh
Wb8Pa2Ed5CGNkTku59mCssQgSaBuRtmn159eq6P0HLHeLNKbcmmoU4Ljn8FE3EtH
FPPX85tQv1kp+uZkqxmPx5aIBilubF26XEaem8gqFZki72b5qph2/1ZEO4iMBP4H
1W9GEQXApbWN08l7XA5OzP/IvHZatCIkfoJEiuTQVMXSxAqvpebsud7b5Y9iC0fl
vXZnoi1KIyAtkKQGfI5EZwNl/lc/2okY0mOMQVpLFLgjOT2tBj4+MC6K60ErQNtv
ohdCRNTYXOEUkPFoEd2RdBmZyYc0bTP5kvQ/yhHwm1RE5O+31CWiUmskjpdRh//D
xHjyLF9e55wcYetlKbYKlxsAC7/Gz/gtJpkv1eWtj+yJuUOF0hIxcMNBlt0FLO5d
Ouc8ixSWVpr2VQ74dlh/pqhMXt+66dp+i04K1jjkWESqU9y122QgVgTAZDSmIxqk
oaFDkv5o6jIpUFuaeMFx0r+fuR8YBa4Jf1rNQ07TNNnKO4ibQW0Hp15tZLJzGII9
8qXf47fQI4embEZmi5B10Uq4MXYgBP5THPfqzx8W6tM+m5Gig5jhW8JmexomFL56
V8pb+mB+Db6+tiXBD3syx89A+euECMWr4zi2nIDX+5nOfAmxfZr9Yw+P1sXTRZ3u
JT6TbH2V2sJlGGVceJj5MMt6fjN+LqtLLhpeaAPhlJyZV1u/LVn7M2oEePHxpiUD
NZM3wtyIxOQhf9txJVEvxdWlAO6YyW6p1zJU7YO1oAVmHh2bI+9VuEQwiDHX8wvD
i3DExzAt1Ek3drVi3F9sHSlDR5+8SDv02lxfhJKqpfy34DE43WOVObpJOje6jDxx
qQvVvkBQOmMhdaXE2+yyPXOyU3Ppu7mo161xQuAygUtBLVoW+/ZI1nLAG2xDAlmh
MCyfC+qaeT3Jhhg+m8gyMu+sVdOek2BmoxvspR4ZzBrafV8BS4MtnUD4nMgNOXMK
cPbBT/Swb/FVXnBLlC/kuIrxGw9ieMcMRioyYqjgWQHZkZFGO3xBN3YFM1M7BxpD
8WMBs819oBI/UXSmekEVLACOqdvBwB2pX0X1AdYJHKQd0QDXYiqWb8lUMYL0U1hk
JwFu3HjZz7VX/VN23D0kzMnS+jj+W9OyQijFcqm7e7mkQ6oeVg7aItj1b68hbrWU
GI0ifElptTvjPTCm2FCi4lxViVqYI1P0A8RU1mzfMOUATxn5aPDRgHZiRTa1Gbh5
3o+jvo52Y1tVzE4hsbPb7QNaqvck++CqSR7CJtYTKPZawyrXJJN3Ikwy5KIv3CMz
kEWnvv/8JBg3QnRE8g0+dOBUr63gJYn2bhS3sD9bbcTZZJdS+RKbqJEWWr3oMcN9
BsSxED4eIdSnz1uL4gUso2+6vYrHjvxkHtLhLAUnu1Q3nQU+9eqVzwDFAGVvtnrR
uPqFdd9VMpHPRE6EugP5WIvk/IgKtnYM3iF0x/xu7e9d4V8cOA3qMfoADE/swWNK
UcYLc9lKPSZlPlJUU+vfUTzZLXzd1pkMpgqARuvN7UNJYyl+Hf7gydpVuMoGSFnO
pHYsrNez8IoOgHeYz21CSvHbd7Rb2O0poYIqLccNi9FOsrEGe0jBVdA66QZAMJJL
He8YEJxibPQkwDlouZhQM7hl+AOGD0uewTI3mWPMkuhzuoHvEC3jKa/sO3QBcHBM
dq43y0RqjMSV0Wzf/bym8LIhxqWNVqgrccJ9P2kA64WVTE4MTvP1v9u7Dc+4QqHr
yUUYGSe9Pq+YZaVdYUXdXkzafDid1HSS8aVgBVL4Tayvu+dsVGa6p1XpZkHFbNxI
OjSjSYCTBDyV/c40hEibfKmSICJq8zFC6yXmMnw+slz/WGxtoySsndC40l5idbsx
6hasGacz8/1YdBl0zzICvJ7xkM8fr7WS2Ee4Zqg8Pm03hy0z2M4wepTDkoCv0Dao
amTF41U6AOXKhztivrwXJqs8AkFnG3h5vkX0ULSL8VC+KwaYVi4C4Z6aCvgDFfPn
iddV6xYyOWIPkaQHV6yLWhnuQFGvCFzgr0/MRtl0J9e19Tby6F0eYm8c8Y5gj8p8
aL/sJwrpfL0ePBVizu9ZbPVJmD0b+PKNIS/42QKIU1DIc838tNeFRM3r2X8sqMap
MNd+rYSiz1aV37luTZdBOghFX1K6IUUHu9h4mvccCf8c/pNsQUTqc7RUGPOAGaiM
WiUuEf9JRc2rZP1R0nmgHCM8uvkHmNBRXZl4waSL/4tQ+x/TzvDKqc3vpgIzasPV
cA9uvMUuONgCaLGiilAx01lJnDqLSoQXqJR+ap+fB99f0tATpX4/88WGyfAKwEFx
iXHcQXsJvCFfgjYMxMZIYsc8TXx5T/8J4Je+Uvy3/ThBMiZKYRTpZ8l8vjCfoFLu
F9ISyzCCZ9B1FP4VRjTMyTwX0Ezy0xhxtYWS+KbzQqfpz9Vv6Eayibe0YZcbwjBe
jpp5/t3a+2spUp0b24fLLPqcUMUYkdSTbdtQ2jnCB09cpHJDTrK/ioO1dk/PnD3D
c4i87rye49WssbGc6N+t7TDWgaHmXtgrcoNf/Ud54Jxqn8rr84SNhi+ASG3jX2Xq
RKsRfeLZDyDrbGuLJkyTSB67HHyveHGsQ32CI8ZI8s2QjL5vAhbw2OBGZ0z8AcEl
hT1/DVBJTV3OkN6Tf1l33bfT7dDP+fEmtlz8s67YRu9igaebOhd8au+1DZY9TIlx
n2nR0IzhadDKxrg1uAb1cRrWJjwlzn02v4oZtB7OG4APNHBpqO034S13bp0RNAQ5
oNcrqiHbniznNkhEnzGWalkZnqVCF6pE1NcnphkBRm7RCjw3dFG71RIeXZ3J//Un
XCoGspu1oPRzDQgBARzyJ2xm0CFSVGvYkvxM3OhhaVw5e4R7r1UzLDZKi9ZaKHGt
ZDL99/Of758SwNjEIbSPdr/EtHuzy8bmpv/Pvu+dWHWE38J7FFN8fx7KyBec/t/s
I2R/ZmykYN7+/eIv/tHulH4tP+rGv9n1Y0/n9ujVJbCqnLmDTMIupc5c0akH6qvD
m3Ioly7IBUUyvH8j7EBgrWtUNPyhMJ7alp5BAH7SEsDeFqfjHpiBpB/hr86S3N36
3IhYD2t/OrB2+rNEVY4dULHlis9IdEaDON6dT02Go6irD9Z0S5iwpHaG7fyvbznB
5QZw9ZDxeVpxg3X22Uz1r20jj1VTUx/5xDMTft6YHPZ49xfuVh0K+AyaM87HYZvM
+SsDhshOODbqNUggvRutjvH2UuxdVjjwop88jgz23asC8uvSITpny98DL0s/+AIS
RQFhQsvinTHQkegFQoOBDPFC94O3VCavFQqRbfi//vCcvsDNXmY+cBZrSjrXhmlM
wVT6qzkCbRy7pTJFmJDsrhBoZV2LHxjI+dKKbnyHBDjsYPUZbwQGiIorWJyx8b2l
WFqwQikhc5e6of8PJp8LRltFClMbR5WoiacZ/RGfUeSK/rtwXmfwKxVMVhXWphYc
dLuCU1BqAdzyCYLZa9eZtUhkvFN0mE5U5qOtbc0LJrLaUmbxoporKfB8UdblsTfA
gvqwZRqFmrW28t151Ht1D5FaRVaFUDoqhqggQXfcHOMqa+2LduUGstwiCks7eYIu
wpf//kLpHgha/DphRSeTSGEvHlmLrJBTIXyatbU79x0oKXUasYhVdigbGUFkqUuc
w4Ga9L1oeXxiTzNZVb/8r/bzLNed2ux8okFkv+oLFCF3PpCTBeGUh0RaXxRDkw3B
2uO5krd0mSBFwJlKFY1Kh2iwjhMQ96DYE98j65Ne0M3xWruSSNqjPZuLlc79ToQV
jNv7y4FVlScwQe2rpIyj0sbmjuorn0mYw4TST7b9E4C94ANJ3eVAzytUOUyO7zMp
CTWVnQe7lfPJpAxf1PYgKp4hNsgtDR48I+pwZGVsmKaHVitRE5JTkMemAaS75otD
XNvhuKlmWfUnsCgfYYqo/Vv3YhkogmjUkDYcljPazbGjImNK6GIz4lqbRU4ZfE1l
QRDrz2DQIGDobqsawhBr69KvFam4HoBt4J87nmJa538jLR7bcv/HnoQ+pcNj0lDB
ojH/60uIW0boQBD8A7xVfR0oah8YFElbAWdg8qjv9/TVui0My57oBXS0fHu/xTcr
Crnpklkpqdob/ScpuXtmLLmuG/JYxFuK51q6nBljKdruYXHnrr7e5epb6s2awb1Y
DfJPgcs/o+NbVpxDfjkVph/XU9Ms/lqZwUpoz6byb/2fW5U08Q3FjNFn2EPa8wDm
rO+NjrVmEpsNib6tqb88h76aO21qF4Ywlv1Vza7GahdR8x/Mzkunm3KFHleI3BY5
5OqAbwwCjhJaFCwcMJJcnyqez9fE7F2g27vwo4QIFN8c8hRvugTZLMyMs2m1vZK8
S3IFAkZsurSfEBGeYntQbst03+EF+jhQDoSnKxoai5QR4NuDxgA655bjJoaQD5AY
debwrii41T0khG6j9P6UeDgfmDUU0HSNeeLak/q7LZ2hrVxPcejFAS0qbB383BZ/
fhGm9tTbIc7+YBOC+xAiWmdGLypMcj3QZpisbtvxNPxnKmEACxG0D/L44WoakJYb
8uMooJIncpcoJT7TIgFVZ8mFqvxM6LcvsGqNXHK65++0DlebhUr8F4KncNuRUhqo
Wx46U6Ou2dsosfciyyFmFCuJdytWg8FppwTwVUIteCaOCTjZsJCPaUgurVI3fyUi
K0OIv7DeXFAMTSQykqOJfNtODnWr1D4ILybarPOHZgk0pN+iDQDOBwImMDJrE4z/
3B9VUvCgJ6G/qOcE3wNmS4jQWTdwQZMWhrBt4AqXT2vpMVOipZiH5S/JZEGkrHzF
xvdR8Ef2cD4R80qOKGVGJ0FpKicRTqw+3TePbbOA6pzaQ6TH/gdRUUHMl7ZGXpkf
jF09c+Uutr/WEXMf/XVZgnEqLhiWEVkwubgkYhFqzFJO9zlcM+Yybus1mINc0PqC
sYVHnyFmkejDUQnddVxUzZJ3u2TGdwSHUDfs+yUji9gNzuCE0Z5jBSAnaE3TFcTa
FYNzlPnod6AQ9sePV2EUyXoHDlcXzhb+1IHmTp3ZeodoxuchAh30f5pL8C6YUAx3
ohn2lxGcvwLiPIwbJcU5OdYAYuIHqh7BLL0qkp8XE1TiUDHPSvNiSkYfERu43BRg
ao/4S51I580j4g9wRhtaUthWRC7L658umJYOm/0JI3vt44HO7J7RMo03uQN7Jk3V
q5LLtYzkg3vcsSGo27u3WiNhaOrBnnxvHtIxCvWNTm/MB+Kl2GQFkBEfslLbtqw/
G2prfsf0eniNOkcev970OMsetT+Ng6hghnNvKA+Tg2QnhB9RKpd5m0JuXHBmzD6A
PZ0TIl4Mxy5jSyoohC42XgmfLtVkbdVUKnBIh6R0prnxtdoIiABVCUXQbYr7qvCq
NzrSERs/0KWp8FyzLIqREipBW+tVGac5J0BFuejkAFYxFhhzuPnOLy3qp/7hJ9+U
rO/ZElRIIsAMOa5HNhUqZopgJXAoxjujrOe8Rtl7pWPgMpUH/Lhgu16nO90TUKv3
ozMG0qr18m2KKoXvz9u8MVqN193FpIqtKwHub71ScFlaCxYXjAe2zGFmTUtqSpNt
r+oCqMWqZyuT7L5k4mKPu3fIs5lPgfl43D+wYkMs8LcCnzRIla+7XWmq6UywbySw
DCgbNu2wWGyWXALJsZvpKDrP3skQkiMy21X0ZCeUpz+2zmvGu6cAAPE+NmESlTxw
XaZyeZ8du6fBBtAnh812236oRBUhvGw98ydNBitUoiijj5GM5NE5/5JEg9KrwaKN
yR4Fe2QdkNod5qxcxmFdIikQ+uBqKuzDoUlqMFb35a6e0BJ6sXDozHNCpdgBsYdu
wn1nPbWP3S+F6DURSajOoBUFeD/nLfCr/s9AsuRVHdeZCAf9P3KEIvl+aLMM8ayK
a0JhSfjwEzbEKZvNR+qRKxC7x95ZdRL0efIjDM8LTiuw9VFF7AkoIZUrRTxzNGAd
dLh39lvCCFScEE6OK/96n1MsjIN6GOR+32b981vn2bEwMi5gb6W/5CxRXAp5xL2B
FX1goSaoA2LKM3J3E3C7Z6vR55cPlC7LFQ2zRCJBGDyaJ0dhluXek29qDqUP8eB8
3UbBsItd3s6Kz+GY48KM7dnQGGb1jdurVTgs4Cyx6iinAR+/FwzI5MqW86NjLcmg
2i4LikaEhw/6e4MrNTaci+z2eyuCOxZXpiJAfUmsCjyddFhX6bdpDNcmJK+d1x68
sd0+olN9A0A4kAjR5xQaFf9lRAskkZnEy3aHtDwCXYqu5EKGIf04JEsqjbRMD6qV
ZSIzYoNjWDNk//BFp59Qw5a1XqORSXn2d98uxBT/qYaqOak1rovxfKRmZjVj5CTS
NoxoTFbixq+jJ/9gm0Bc0RItRL/4rYfiREfpEJW4X7Uo3lmi+rumXA5yM2ye4Yjj
XcSm+kzljOjxe3ZGEVMmcC/xnzSQa0YlPXL6fTrGCQBRXsHCS3zGE4kGDK+3W6mt
dS+56UIDWoBUBHtIkEGyNKnLQ9q+d2dAb9DgDunS+XyCQZ9HJQjSuKdEn61P/Mif
fbTlL0pD7titWW3fU8V/Yhimahy6qV7T3/y1GYDNX8BDrqdS4Kh+p86+z7VaLr3z
WbvfekOVzy3cS3DxUupKNs/Esrqd2drQA0o/t3zr/HIhEDp7uKzQM8pGn/iVBFAq
1SH5lHhSEA9JaMe88hmr8g==
`pragma protect end_protected
