// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DwsLNKQNzujqb7PrcvbAfiLg5iGSgcIs3HRCQ8WAvwO2waOmDyMTgEKeSSnpjblJ
kP4dcnSG3MKxl0d3QPIJd0pz1AVRZ3atxWz+Ijup9164pWuZOgvxo8raHDi308wG
9uqT8fPOzT18EeiWNAXngPGL3thgKzoRjTcEMoUya48=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5824)
YicX2LLTX6Bz8cgC7CBndpMRsIe02FuGlu8bDQgMFgcLIvV3arCZQOR9uXrmcIDX
bTOq7apO/o7Hrj7l9L8QsDgeYZkrhMjsBhgh+909VArLAsWGwLqYcBCCc14ZAr3i
kUKo9zq+IQF7rh1FMiN1bQ7yy//JG2g+lQiO089j+d0Y6TCcaMg7XQ0w8NEk0Jy6
NNz8KzjeDRH0U4hV3+BdEd+4w516031PEh43+UlTjcLBhWW47Lw7ehVxAISc2G8t
aYEGtnIlfn4LmV+oNPauI8v4TQxopDlGx5yjX8FFXdYZXoM2Ty5wJjCPGV/KnCh+
n7tpFPMhT121asKm0jORcwfi+IO5NWMH3HfiAhdPOH3wP1jVIxswHRO5UtE2EuAN
sLAHY2TpFFWB6h9eRob1Qgvrjx6LBE8OzuOvjcwGPB0lEMeapzUTM/RSRacHRyBr
AtBnYJt3P8kcEI0AiTMmE7/mBsWnpEZx5DmLIR0POyCuoP4KBjAqzFDjgHqhUhj6
jMAC4zq7Rw32c33IayAuooUux3+u0kseuQhzXviUdTJEAyIUKEgmdlnVfR5QXZIR
vTO2A8dGFTEV0SU2K8fbbzw6Qjy3+gISe+08J1rPzLGLkiX5FxDr5iH+WBUSZB3e
b0TMcZD7FA3dgmiKEczUeT6M/KG0hytZShXCGy439loAxM6ywdhjM7d3IjjgEE31
CX/5fG5b9DvGRfqMnyuF2ea6F6qNpJ39GcktGPHBk8f1+lVrU1w4+OJq91e9J25G
kp/wEk28R5e7UThjsfLw09CqW6Uc13GY52n51HxYc+QjQBGeXaVpTUF/pnk0X/FI
wEc8WbzPetNL3NO8ReEwY6J3r02gOQfPH1+68BwjW23ta48bkmwzOy9nlhQDKgqY
AcDsngPonu48/8qvc2T5eWv7bkCLqyvot8L3GFkAOEMnACriT5kYs2Hqtdul5WVy
aKcRp1D9beQKCkyvrSW7nnnrAfsrOc85srecy/4ifoGzjPcHk/hFDnxOb1LRGS9J
Vw3ovhbTSKKkCHytcerzyPrElOXDJoAEe0JLLBmO0CyDXyREwwH9IBepjNB38Ygb
uQZrsRlDipRChLnYADtcHZ+Fmfi7T+nzSjXKn6KmrjdayTtXD7cF71Uvr2Ar6Tr/
vvtXrQ6WnW8kEX0nFu6Sq/QeAqXqRUIgaXyfY71ymuapjam1EQXPe9z1ibhXOQJD
9ro32Dm5lRn3aHWnMNlLkjm72NdBotdnfEteGWAisMEYhQPkEUJ8QIBs4/xBfcwV
iNgIPd/MX/JLEekUE7QPUuOv/VD3MaO/HwHdG+PMDc3UtTnr7sgspZURd/yo+W+9
17mTDgEjqVbQ0jnE4HDSPshGvuRYptvESU1CfU4vJW2yHKADJklBn5eZyCcBulWy
kPnXt5IbdoQ0ehEwNVQsJD+OmTMDKSVyi9EJiY6b4GvE7RCQbjSPUsJZ83oBBLXl
RiFSk+cxiaQwMXXG7/alpjg1xP/D+9DkfWO/xsKqr5XYnoXwGg8q0rSuHzRs8Wx1
te6JksaPiNf7JjrctpACg6XhkHGlbueuBqwX1hVOLFyfFOOLrNTgrfRmSVAltbvK
uvRfRA2FJO6XSuVVoMz87Y1JqcHeysEHvkQ1smJykkrGDxKUFfVP98gY+vLx9MAY
QlPRGEZiTqPA6dKWTSJSU/h/CEUbRsS7q9ktKZbG7e9Bqb6z0mVgwiwoGbWf56vS
1jQ2WL5cJuBjb2NCyV2C52s4HpBeO/54WhXe4LyoteZJGz32UI7QfmINeVFt+Ua3
EjfL1rd5hnzsapIqnntOqi4gEYvMHX+BBdYS/xZff8ZPkIOdIWFQ8+j+3llk1q1b
zJ9a4+J0kS0mZYPx5wxmiiHc+phzoE1lktMW8NN8JM0YUOXz83VSSxY8EBIdFmBf
Ge0EobqmbsEiXRG7m2ZR/D/JIlg7eAbpXsTosTLxQKg7EVOwgAq5qkFmaYoDmIjT
q50q4G+3E9WooMo4iO5F9VOb8RjvtwVuaMe1hKggzSxpwdJInWRzU5R71IKQuB6f
pR9m5QtZl5T/DH29DD774EJpVbp/kYcLlANsiU7YwCl+tvAt2pe/U0BPjBuCYXU7
heQkD+4H4F/XOnMliQrLpf61YjGHjiGFDmFo94mFzcyD+NiLlnxXmavAsF7EvnVm
g4azxsBVOqZrLvrSV0v8GmwIhbq//F1KtiNpWsIqmypRraLGviSbhWEBhvvh8XPI
0IGetXWgEjL4xXd++Ob38L4Lp//a2h4WZ1vDhu4sWZpBNZSF6Jno6dwEmXhedYsE
87pJt9P7J+MwaE8P61FO76F7ss0pI7aF4uuy5NmPSHRJ0pzQ12lI9sZTNoNUybvp
z4kSHhrFZsDOfhGteay/qLPHsh8nNIlmRwsO0Hx7nepDuQHRBJn9xGEVh/Pca/ml
Hhe6N7Eu05ZdI2VA9yfmg02sRF4bBc81/bqhNDpKcQh0gNZCg5rLKgfG/YiPV+wa
ZLvJ2OPrwFLTi8kga/lpl0MLjbs7ww79Q/cNlsVKxETK9u3WPxHdZ8pXcnyiWTyQ
GprZXJd/os55+A76aaTqgSbTNVIuPcHHXQ9vW0KnS6yZ+NPs5jFdnDXBffgirUj4
NAAseHn+9wRnLohiLoyYFtKaUW4QJg8uhw5TRboerQfMY1k0rJvUnsu3I3PBFG42
XGbf2vbLAWYz5fCftHTV6N8wTJ0UhEEiptHuCGmSgThtAOIcEkLyiPEzOaoY1QfB
KLLiyq/aKyaAhYSMHsW5Zmv7iqatMu/3HWpEmpmE0KokHu8eUU13xmGPYX3Gv9s/
ymeN1Qt6ZckHGPM990XtoMZFuUz8opxWzryH4mNW5H1SLFSgJw3mAx1r3Zxvsdo/
umCOHy4CoyJG6g5P883mOBiVjNNsHxePURa/yajM6waFETXckEPbqOTHWV710UId
XtBd+r1oSWYus0ipTCMaE5cKcn+Y+JkID2aAJUy5whQsm0GfF6NiT8XNg5xqc6Rr
U9Zky0Jdm4eotU9XXIJidaCPll2QjU2ukyaoYyQktunUSoIkNjSFrmaEaZQlDESU
1exfQ5oRikjdWsavIWR6pZNqK5g8wuAtBAZNC/xA2eOsUHsCP2AcbndwIADbMdH4
Q/EsGXLL+Uo54PsUBXMDnLsQ3GshXpNQ0MMQmMezB38ZjYdY3GTCAZi8UAOa4MOr
1O6gAjERJWvvtDddqH8GAi0qNx8me8DvJHMe0Bw+47wzqqSxr2gtuN1GhgbrtITo
2jmBsj3N4lgHNcQvuKyZDMCI8IiyP1gTQPAgUVx4Wh9UfGsSryXhUrlqB+JS7VYU
Y6L3emNxGf25Dv0VZv8+3Q0pKEB3jm6liESNGU9W/8MxtUzvxKpIKa4S0Jmm/5Ic
0WrldWug02x/TPuHr6NZrGxKTaNpfmOj5eHACAvKCNkcm0AYojVqb5+bs8+asQy/
XjS9mPnGRPtFAoM4UzCtiUCMcUadlVg4/8HqpCZnFDaGY2Jm7g43RIo6axH32mcS
O8TxzXyGORrEFy2XNSotD/IlvSD5aUtvs4MhfNjdFC+vic8xZgU0eI1zQSO30SB1
a0a1QvpCnE8YSHrs3oDXhNOnTiXYkR77sR1cxRQjM7UWBCWeqKaZpBJvDCYqlJ7G
h5m6KBVWx2az0umOWkgBUrtkWUWuTuf7sZKUJKRNMQJM0zPTTwn75NBZyErg7I7O
Dtr2R2lWI6XZuSH9xcWZFV5sPH8OaKQs85mSYO825PwjND7iDVTFY/OibBCTr8RP
l6BJH14230jYz/sDr9Vt2J7HMTMRCTbbYM293tr5BWMwrqlNA0NVKG+HwFeAiGYZ
ztQ9WBMPcivvSPbBmIohZzfM6VW6uWvm8tnQrg46xpoHO1iATR7BiU65Z3BLYJiz
RXDEac1Fpa2N0eLD/7dUwO8jxSnh86DKYwLrAzpBMTwV1JpruvPyle3EXZTo2CYI
WNzyclCGEbq4zdJLPJs9uaVXfZ4FZPNgS7YxQ9hbJbTWvaujgPeQgu1tokGEOkq7
Gr73bd1aBUoRvM1gEifeA117yel10Ob1sZ0wNT/VBEh7j+YZUlc5O3r0i/G9yhTm
KpwuuBhA6EA6I3YvLSYGQr9Z8j0V+iVTfy6BxN1k/kgpGwulu9suNAYGkXR5S7BO
m6auExhotoFrxVdm/t/ev3Gf797o5mfJPGHMfDIsxhsUnXPz1NUCUE6byJfJqRT/
l/YfmEu+P+exH/Yw264vHKiXTDeipDWF78M7D3jE1XGcUO/TzvklDmQ+5GChxPKG
qYWPVNjSRr5d5MiRYpF3EY/dXwJQmvzsSu6ufQTKeFOp3qszHixa97n/51CsddSx
tKmWd9jqVL1uW32V5/8UagQnozWAgAuR4/CWFCFjsAOvnnWvZqHD/tKd5Tw5lUrN
hY50cnEnMpZwZ0PT1uGlbYd4I3zsYpzcBnI97OFukNAW38u35Y1er0gH9/8dj8wu
lmaEySggDdJeMJo5jsW67W923tLtaYUs+JljAFyO8+VdOP2IAc4SNSdfOnH2gKnz
6agtIJK539CmNegB9bAcOq+Q93r6nLFXv+P6qtLFZdO9HWzXa7NKyLO6aYEMsLqS
M44/SvdOA05bKj/5jCJmkFbABwMCevoO0PMFBMTqvNb7INrPiAo+lCwqqmc4KO5j
MxOOxPLejbT/5xfvE3pNNOUTcCesMB3IybAk+/n+jSpefn1wN9/xTpwS6qGaEmf4
thHw4ii2NiU7hgStq2WsF+Z7Em4AGVShdI9X8iJlcSv6Xt4TGKzdJA1RrzUd51MH
TY7r1KPzCieg8AMvYH/AOMH8wK1v3hyDKbfAyd/JKQpD3muULPOrW6AgbTHXKFrT
FTD21bYrBsp1zFinmCsgliW+JDjhy9DPHh2x1C7ftHisBM19gCO5fAl/d6gyuJLK
4DyRvv7kZtW2W7jztPy+vSOPBvV+FUF/mKcxklu09zUqwsWf17Gqe/gKRnNd2PU9
QaWYid7LCcVmjA5FE5j1hIQcvXx86QeC1nRPLxQns9Bk36kJZU0jeoNu9wuVAFLm
g/WJfivgREllFpxi21o+PUgJTPTD0QUZBye0DPSAA31tleei93PUAr0oteepnAfE
tvlv6gs/Qswb5j7XQcwa14kv4s/L50w8ODrowGB8FwRiuc52aYCuuBzWb+/UG9vm
2i2u5qBjdGfMnRxevvvhGKPGhfvYCn4nEPK20U4yOM3sFjoIHCOSudrfYfH5pYD9
sRIdhTpo8/E95hDYvz6kKHQZv4cmEwM9kshlteMd53RLN4vUzR9n9KOYCu3GvhjZ
awkQ2dKwk13RcuFsvjdQ0LLLdel2VAFugY4Xy2tsUtz/O2KCn7O8xh4FG9Vkoc0w
t/cNj/99ILjYaX5QqJa9hb/pRVKoNbic2r9mGyReIJ7H8nejYmx8FFq5Z6JcOumX
O6o/jeyzK255qmZJ/k4SIBNsxBVhkucGp94ixpOwhD3lSkOsg01lO7dzMSdw1m1L
KvVi7xmSfadcQeqgsUmvp5SRaF3rV8hUvhrzGVVi6cp83MRUN0+J/UGR7eFgNywx
WndBSRoxY2jKASSCa9fXhuDqtXHANnQAwITTK6FY6xJLRzbuSStuFPdfQ/5hL9F6
Toab6wyubR3qwk2MZkQEPMxLgUUxSIQB8GgbUqXita6+9c8KpFN7UrWr0L9SCgRF
Ui8GVmaiVFqZbswYYJIiGzZTjUhQ5Lpt76LqcFtzevJ7lkUNpt1Vh79r8ToaA98Z
07Eo7N9sUVGcPYB3vyMnLKIec5OPuaLshz3V8dE+taSrd+cJ/E+ZdA1Q38yb0a+4
ruBpPu+4A1JOtroimwYk8gTP+TuvYIdndZOSSChKZVc95dJpIhxIBcX5lrV/22t3
6ps7ZEwU7DpfaFaKqeQJEBc5g8wGdDA35EC84LGfGBVQuuiBK7h5vXH7SkIbG8sW
HWeTUZ51AutPPCuB0SOiq4HSsp4yrGfRHARZfV5Uzy4dvTm2xWeknvZ29FasRB+j
6lVJJj3bJs9BnO7b95Hc3xHe67mxtF/VLxwS6h0X/EeTb/1Hb1WZkBsL323igTGW
LoeYRkppxqUvwcPi8CzGiRlKIvT4k0dBaNcF7cuOmtRUMbx9q+PBFeJL9ycLG9IO
tPa36KTGdGKAz/jncUWJYmsWd2s1HJAQOHj3kXf/NW6vqg7jx5Gj2HKFyqkCreIt
aBhG6Yr1hDvS2AvCXXRpQyh9WocKb7Ko+zbWV+Y80YsHzbncfHv5akxp9XzI2Hqa
WXvIu4mZAlKcN325MLE9spwKlFi+GDa0DWCCdfT3oBan9kb4hXVat374sVbS8ZGD
TxiOi3tdwUVzHNM4J7UewdQYI3gxtWSWh6SMEMs/Em1qzuic8t9CyHVEty7Fs3nG
aJX7b1kW8HuOcIiyXwFi+kFdGje/RPewTt1aBqVWeHUxBkrky1CMcPZdMvbdehbJ
lhjOSg500TsjDeI0xjS8W0s6hagVrRT0uFBSN4BpqblwlShnBCUijNPUPpQ5KrDC
BCvBl24x2cGg+QCvKIrvoGYIbD+WCmLZz5U4/v1Tgi3mUkFkaMWeS3kibcyZ7my6
zuDfAvoJZE3IdzJDtFqyfnqoV3luwfsK9GQcIMiyOoMDV3QJYOwz02zSADVu2fRN
6IKIHszU+lpI2YBEGQS5FxvLIM0wGENE7M7vouWFKjBSn0AZKDyOSYvfGxBWh16L
pqUVKEhRfAI/xqLY8sZ3gNUXuhYVVX7ENncAHmmoTIxCfHGcSSlM1jW7HaXYATd7
DAKZXFGg5Y0aeRUjSV9JGusNTWQ4zt3XastI+pDASIoy4N38agtdh+F3iNLLUML6
XaVC7vNrTQ5nlZfqshTAkRNZYRjS1RQALdlLq3RDJXmkK6bXFtCe8rcJMjdCK3y5
SNPh6exL8S9KlZMY3UKN72CgVKrb5HZfZgGnOq8O0P0lX83Y4AQUwK0xzcgNOwhJ
2l68ma07/dX6GfZHRmz8NsXZM6o9ULyFr2pcsY6ipv4ys8rewWgSUzM/zdKlaOnp
aLkcv20Q7DR4RsZ09/OiccHy8M6dVZ3wYUvUNpaV5IBFp0azmT2h323Qv2GwSU65
PVQprg+kWnrMAHrVGnNLSc4/vxz/+r8Td/ovyeTD84cwYdeLFfq1RTsK2d9Mh/k7
4srIExFrLnd6X1XnpSx+ldD9LDFUYjldpBALKdFTozLllKwsUmDTcR47GdDmZU3k
IsnIBcKOXoju9vLZV5NFeUoz703+ajIl+jQeUM1WUIj9H4WwVqrDlmrKKkl9V3VS
LI/WKPw7UJWCoN/903W8VbL5vk1M17rk7WV/2lPFJqfXR1LfNHDYrxhXrF99yq1K
K8v1xR3GhdJ0xe02MN/+yFgK7pNpkXAFmko0TXK74ZlQMHo44jRlh/XrwC64IWR8
EmL7vT5hKVavhNFvwPq2APqArYEj9mxpx6mB1ZGgjr2nZf5RzZFZtzUrNht9l8eO
ySRsQL+mVlCuqmJ505PGljhkyTwJZkxO8x/ZxtlwAMldQF6bREI4QLsSkCFX1rYR
ch3USgNKv0uvZ+XVhfACVm0+rpSYboIASywOj6l1ge5laRU2CS5yMUGBMPnEwuGD
weY7tWtqJ7a/owidWxCL2LgvuB2iz6ugvVWSCBABuAlj3YnXY6VtjvUH4xEYOHUp
Olk0YOOCz7HaqZ0JfJAzv9BhCoik5nWTjnOFZZMM4JJLSf1nhHJJhNcYRVM5Ded3
LdjZzqsxQ2yZ/8Muxz3gbA==
`pragma protect end_protected
