// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:46 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GGzWbmhZHMsHo9c0AAaGdcuEJssvXpzCrOCORy0oyntbd2rDac1823Aau1L7lMqS
A3kmRrGceXIURD7s2Ru0PAAmUl14UvDnBfiw2el4WGecZs5Wof6mbnaBpH+hti2d
ODZJsm2OuZC7zJY4+GTTovtBFq6xrdc+qAMPp8akego=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31456)
p0qA97mRBrkcyH4/YV82HcJcivC9/eULYpkMU03XXVdTsHg/QKQZnOr6Ndob/fx0
SgeTnY298vYPhVR7kz5dVBEJdkOYteSshzwUi4Sy7Cw8EytyTPyQxXl/PUbWt7/6
TEI3IQDemfppXSyHyDrsciFg/QORrZ5JGnWuCWazt7bGqGYo6ei7B926pAuuwK3S
bNJC5fYcRYov3auin/nK/wv0RtYGe7/Fu8qStb2gx5lq6E73iVh0H4mHQl3iZxd/
z6RYWIyumjmG5XDCuA/AQKqGv4MR1Fe3lB2ifXNe0Z8jYXn9bwhDjQWcZzVcOlZp
NFdKA1bfortRAO8ukZFf7f0h1WiT3Y3L2Qp7s8FVdeaNSdH130UsHZ3kdpj2qlDI
T8JedU8aMP+Zd+bEbM0/XhWiMvVK4mxCXy3n2bKkZgYOIL2DoSElsLaUu51mj6do
7GjLwjYhSFNBAtF4zBFQ4DyROT7YCWB1YXfBSNTtRLuYi+zUkK2tQGQf2qoBCvte
299Ex0YOiSR6KZgGpKBKRyn5aBY5jOv9iPdqNnqE/CZOJMLS8QgHEZaAb42Ig1X2
Dtjwqjb6BRIyLuH0FGKkQ5+tISIiqZ7WQCYyUOKlkHyDWXga0sz5O7Lj7Fi8S7dl
VmHSmCx1wGGEcIHGX0IVXzX5I5f/GTCHdnaKUd4XEWDIxINuEH5OE/wNJdjgKmTT
BNG8e/zK2i/ZocktppNsjZHvbMW2+nuqH4naC7qNwgk34Hy87CBsj9PiZS/aWDcU
t8Rg8Om08VU9Re74fZqvC7jyr3i7EI0ix3sfrku2BLQG/DfrOL005YDuNUVmp8Xq
//t+3WVhqeqoTmF4bMsvPX04+EBe//KEW8vC5/NSDUJZBPCjRmhWMRetRULjpzsR
7qzi0BPMlc4EBxlNpyv3MEoGX73sZi0W72JUrbOP1zjFbS5UGwb+Jifvantzbw1b
iVGYzxVeaqiMgOv3eA/qj/U0v4qXQmudiKTJ71gcOKZR8oxCl/eM2aoApp6ZiLba
6ODCAabduFHhEUWAO6trUFqxJplpAlnEKRihFehnyGBnjxVyjCeuZMme+mYD3yZt
gpfYK9u16Lb+40t0bLwrjcI6nVpu4jh0PPEgdTMDHsFE9mSp+6EoE7LVCBxAi/rj
yzyqrtUOMFv3ZmicDPTTz7vGsmRJvxXg77jguI7JBNUvPW7mb2rLICIj9AXXvhSw
QbpT2rcudIXuLW3F4UEps1QkUznwENbM5DvF5FPGjOJlBugOzEX9KpKRupTS6S+j
IuKdwC1rs35+aXNmPl3P3dkL8pkHgJs7FI1O08X4edV4v5oEYLt7OhGk6KIORQsd
64jZXMnp6RoZ+H78NuPH+S5ZP3DyrYqYftiIybohrEFkLogj51t8TzvtUH3rH7yg
mnpdpPuKltARmsztqmNH2FcbljIa++sJtCQQ5pszhSVu8yZEBKOGqg1jr9BAJywS
Rn6lrMQSREQZfMTQsmHiZT2Z89UHpFlrc5qnpwQHnHUy4G2drmv116GpgraHV6kl
tnb4ay9l0SvTvmTCJxoSWwLkQC8tqu5O2OcNkErqx52Ky4slen+RqSKBfA59FSX4
Zi0HcTiiEu9QOMOl91e+wc4hmUX2qpKmr84HhaKroOzyUqXFxJdAWCXH6hOIp4st
oWu7VThji2lceg7I2aJN/L1hUzGpC8JEr4GKRgWPkDbFuTjb1NhIYJh/1CMAkRF+
18B8xaBfUDOXohnLwhXRIDk5vxdhwc0iK0qNGBct2rLW+6OKCpJU047VqXJAizOl
cds8tBg70mEAUFiD65YVkHhCWccNiuGJBr5BF6SQhV183Gc7EDgZBeX7Ix2rf+W0
bsAfFiZITt0Auf9vNDeDWclx03TiWMDsb/tI072r2D+xTTzG+E4eJK36l9ZgMVTg
oXHXJjEB7jPJuQt7hEO4ijKgV24oldRU7mQeAIxR8/nIAvrndrAnyvmWiSdIaHuZ
3WrU1L9Czjz9Hpe76mhKQpUjZjU9+GOL5IIKn9wY+b9hzRCpmU9nnZpgNKtQkrme
FTFXshCCrUFSEOUrcb4yFicpkN1YIR5a6kIiRPOHDxoUDA6N01mMY+FZp+bzwZsE
DmYAaEfoea3fNxTJ0U9IGAbbqgZxGrKccxPf87OpS2aQU7MqFP1TFX5trxBmA9A/
GiyefzIdUWilLFsrJR6dgDJcKpWSkG2V5DYw5jSa5GvoHyZJDqK4/p3ooLXgDDO8
AZPFbxQYVCcIr2mQ9rF8wlQlbvqL5uVFN98aqhujVZCIiBiuqLXYST3+MRDYRSgQ
/0Z2KKsQ42Ck37M6X+4qIEiUdXuPd2o3VjyxHWr7FDmZXRhVZRQ5k/KCbJ6PEYqg
z8r5zuc0sfWWAWCsUohKzfBs6hsR4OriQJhuJzyrWe/6SVR7t+RoeXIftgsjHPOv
P1B+6XC4MXkX4NxIe9I3IWuxc2qr1iT6xRbFNuCEabCxVoP+uM6fgdz7bVJqDsYo
ymvXWach0Do+/ECVpWqQBPhje73+JZ9ssAc0EmqizDIkTchGKYm/EdfswyFrNyWa
Hfn1pF3ZYI4Ih0TiPXE8Crv+W7g3ma/9j3F4sXVL1Vye3f6io0NSnZ9ryAhLlZ3p
eA5SxNsRJU+LrRdJqJCaALby9528mWpd4NByGsjKwSXbdUx/V3AM7vaUz1/QMv8J
zT6JczMPzAEv6KJ7rBar53ilus1hh3E4t1JZXuLODW7irkM84W9ogvibjxJZQTJU
RMHZaY1p7HmBr1U9fx57xyTWw/7lII/d176v+zqcEJueX0Ycrc2npSsItBqHGgJI
dWUwb5u90/YzRfv09RrzGcv2nqmvJJI05Xm07ivTOiRQmSz5lnnjEh7J7x5DJOcv
oFrVCnCc7xdM+iEVJmHdOKGWUm5p9lnnRzSk/eU/AwI0eBrYe5KYu9KJ8MKC1jDO
JGVvx5iRH+XGWqgq04+4KNZiUuWtzukA/IT0bMYVQGJZMsII/oay8G/Vd/LVUCPE
pLYh/X/U12vDrlrUPFJ7u48V/UvgAt+iEb2WzLv4/kcIfSQ3VIthamlx6DTHNX8I
iiEl85jo/34AJM/PZjnTaUUokTICEKsmmjAgYaaSzUAdjeOY2WzhFIO7Jato+yiz
9ATen4Qja0DhTQDQr5A+KvEe1fNwUc2NBV3J5Ope5xxGhU82blzE30pTZuw20mEr
Ktvs4+tC91YvcYpP2dmdiEoq/Wkw8UJHdsMXYw0QS/LfbtSpJSyexQJ3W2fm4Xmg
M8AmXZPV6KKXmqD2PZ9XoUkiaFtLHSZI9Ycc9Dc6aXbor8OUHQND85KyeK2JJZX6
8FQI1AJjP3s4uyNdQs3wU8FZ/hecA3KVMhY5maYfxGfGSXojHMyok8huIJ+Xq8YV
RVp70NMYR8RyKoQDs3PgCCsy9CYOJVz6p2KQLO9Fwiiof+XcyFVx1NzObiJA1Fvu
npq2x7OHRLReJIb+NPrk6duXpIHyblVma0SFxgb73goZ1qhvPV23r5NezxGZYVkl
wJadmFWBkpY0v/Z4oUM6GD4Uth3E2eyztSHPVHb5ZQhZ4rjr43764QcZ5voSTkIl
u3D3iN9cD5pEv0dSEDGEExZe2NMpnzyBoNcqxH37vZ/QcCoqOTj/ONbEUE7T0yEE
zp5fFbmkgqEpojCo6Ar/mzqa6nvUJNj8+QYu973VGyRS8zbZDKwcOn3BLnOTJWsn
4UwvzIXSHMYP6LNDcRHgCfHU7WOi7zW4v8MYCQbUTAUySbyZfqI1cWmgqVX1cFub
LR+nCJzLSdfI9GQc4P7cBYq7yOGexZCIckgKZ+GDvWMulOv52yD/6y1HdsL/U5Kv
xT0UTwkMFWKDWGx14W+fe0ftl4055I10UpiApBrpxU23vleIsoAD8pPwhinAUJQq
8yGX1M4Cspl/RAaJMvQTHuwEajNFk4mKa1kXNhUw+IYCFBUCAVzcSc0ABLFYa5Gs
AA2WVmaIkw37ndncdGk6+foARyViTWyduSPC3sYec6oz6V+i8l+i+kL3RfNFVOWp
JtV7Q2TayARxyFEhEiSdaWZtXcCvbBj0S6I23lD1wqO1CaKl8nVAMjXZ4KAIfuLq
PTCGA6F39JMz3NgtJl7CzGEPAaLI4L1VAPPTPOlFDO3sh3c8xKZCRklf8KSoSRCj
X4IOaw5Ux2Uol0naIjQEQxbsM4ih9oO2T177OAW2iAnVZTnBGYQDsi0LSlwY0D2N
E/U7RJr69rVZdLWx+mfrmGTgdqBIRnpdJlQTgW0z97NmWyIX2D37uQqAUaTJK2VN
0X99D2L7cS+jFO7QvkW0zXtDg2tTTIQtniCdSiMMyGxbrGC2mkjfqorj62hObWBy
zDdB/ij/QPazdXq0GTLHW9eQU/2I1RXzZLCPGs8A+RNx04nraFbYOIE8GmMPrNYg
rGhhuyaVhqbUUG2aQikyRxYC4SP1GSjScIf39oEmZgt89k4jQDn3529tOaVBnG6f
huo/Nt2Y5ZIwdrBnafXD3VrB5qx3rFbIWTFP5gfKNj56PJmiv8ODohfwBATmAVX8
btpC5A1sdknR0KR1JjAGxZ4HxehoSgsc+OUq/WmjzvgBgPYxmxRVvKl1qxFuDOzb
Xqoop9ebPWUzYwZdgw7mW47MJAfH4hLQ3msWnySDsC7K3DaDgDeT66MYIbYZBew2
Exg3J1FtqCsx6kEs/Ed4NROQeMrQgNfwZhjdTgtdYZT+FYKlX3KRtuoIU2IT002v
EgyZpHdJZGpNrSjQwMVWWUEpYwfnFVJ34IxITHBXnCDyLK3qt0gUtWnLRBSwnJ1u
97IY/1FbBaUzUtG3MKXl5NF96d+4CNiAG/BlKun+/WLqK2QkYzrjyv5AZ3sWMnbo
owxA8cTVCjoDx6uAXwDx2xZL62ULbPLc8x4tjnNd2lV1SyYgipsBW+UK+VVN+0/N
A4iFu9JTLRXSaWV8GNs3lE2TDe7t8/lkShb5gU1y8Ak/g+AFiQh2/8Bn3TXOrg9I
tq5AyRAXTU2CASxAeEqE3B1xliBzqWhK8oO7ODos1eMYOa2M4hEZDg5LUXPwD0ge
y2fWhrPkgWWUCfVQDltrH6kh1GVHcjGvZ9Vcx1HAitKxdS3HwkUdtGbeT+VpZx1Z
oChf8omvdoF+wbpg54D7z4JNhxX8v9g8nR8AW5vFxftNfM4KdZ6y68ZmH/fbC6nf
PHpdphE5U9nhy7UAq/pGVoRQogK9huP64UTtoGb9bj5CElEIT/oSVX/8Z/vR9Ziz
rbJMmQMJr4RbD+NGLDKEUYGZOFASAph3SO06p0T4wnpq3zhFKtPBIwitYkUddgbw
j8OpRdk5rOCgNBhZOKP89za4OP0iUQWSqbFqRva4qro6dP4wJK6c3Hpus54WM7PO
7LOEbSAeVUzvQUHl8Q4wGBo6rGPNNzxrxmx1QfPFzoX+CyhkU14ODp6qh2PBF/aF
Z/dowkYUT0ZUC5kI8nt+ZXLZbqSa9AXk8QglEHOHD0yPRiRR/712lB6qRy4tkyXX
fx30XUb19iBpCP7Fwb6cRyy9+ZpoQCtKzfN3voOrSu5DzuWGoTfa9s3zefsGuPHh
f/mFrEtSaOpNcSk7DpfueeQmJTZ8M+dTfsNmDZnKesqqlep4uCa1a8YHwGJ0iUaJ
TeN/KT80+I4tbf0OoYlnabZE2bqbx/8bEvuBGRNHb/dMIFjbbv0hmzNHqnAcFyMl
dtL+tF1sbovFivJv7543tsUAMr6K89F9ZZgba5wpyxBRiLW1NW9jIUbsjsVnZM85
xnQ5I5PPDJA9qjfwCHnKZ4sPFzgyMlH1FWmcI3AtDf2gKJZIVD0OkhHz7c5m5WT9
hJz3Wgrd8nR3p0548q7Z4U0OQgP6YfO1IAhdZpVBPkASuGcjKd3rtxx0g2id2U+o
vhXmH711yrCucXc7lpr76H/BqqoPhOn7jtmzvXMRoivhda9zo1uPgnt82VwR7RlT
FvqCxX+WdQK7TI/CzxIs+Y/bYgRX28CogGceVMOO5RT2v6dj+fBvyxfAKi+7xmDX
u6JQqL3qjDbIySjXp3Uqy/SxiAjU6c+IoTgdGs6R6rFTwFMPb3lAiGyoESPQZ0bc
jM66HQDGWtUfC8nPZt0PCqseFzuqjJYLaQ8StDQB1IuE0SgFtMLOZfitzXtST9jO
Bem1MWjJWaQba+upQ77x4S3PgZrVnVCvxK/AukuE364Rf5HebHbglDlOeJWTApcB
ijz7yENaa+D8ts8FzD1/dDcaqmmkoMY9XCSzQ/QrFZKnqMtKXu+YIuEY74Z7ypar
/3ZY1VRbweRWzKlfe/UmwMvDUcPQJcQqx0dcEYQzt678dykEyagUUTXPlbNaw60O
CMyr+fxs3O0SRp+Pp49I0BmYMm03msBpwqxlnnILB355a1dnQdfzmjFRaav7hu1C
xDEg6guI+U1dv+gKn5kSQQyh7jBYZFTeen1oR4GNmyopF0NozPgWCPulySzsUKFt
aFlshBg41XSE1gm94eZoRDOqhHt61HuWB71XTYC7vtcO3v6ZULf3whhzB2t/sgJl
FAyLI3kXcRHlwOpS+QUBpXqKRUE6da5MXTDikcssVGwvSCYLvb6EVehCqnNFbrgv
PW1OdudlHFaMGRoVb1GZ9JQdAna436X46hOWMdZhh3hoDQTC0hFIA1jXoHdtKPSY
WaOsKsjuJGVPJf+q6oUmfylDHscGaql8RoYoHGwiGYjznC44Yvsg5j1r7U5S9/xF
7bUOWzZGFGXfI5lGR+qACMz8oLPACwTVXJ/HKfKcnpOgcNwnR6QYfQGkL38VTJqt
ciz4mI0iul8lwBKx6WlIXLokFxxRunZ6+AMf9D9O1D9l15PIjic76u+vAWAw16qM
gDt8ZzPSE/IFk6UcmhgV2Vhy77WpFSrA3q5xukEyrSlA+sc6GcpVjpkSsHxdiLgK
I+fcVZimB6zRJli/a5QK3ldJ25Gg9/T+KmD5nfz1jntoq7o5ANOYogfkGKd7uWaW
aVX4eChyVyrJY81FdcRgkiHbx7UlisXivyhfiE7pW4Axeiu0ymWu1r6KfB8+si0U
QMggpa7+gd8VQcdO67IYj4z60O934EBV1qHeZ2R5sWSX9Liw1IPxHar0Iag+NbFj
LKiar2ZYhg2GzC4fmsn3sdjZFzRZ1kUquFNpY/eXmLIZbenmeyqY/akQTJXB/EsQ
JlP2OWvD+tpkQO9SNfQqWovXHwoLOZ+TVM8UCoYlhXJ40gJGiNKEY+JVcHYe3fEq
R4nZP3cZ5fyiGK94LykAIrZRowK0XScrN9Rv2w3DP9OKPqHqQaucROXprgipxu0r
I12Vl8KMWA8ztP0ZO6LhnUa/iQAWYIEd9Wqlxx3op0mdrRj5SixLJBHcZLOK09+D
7I7Fj6bqtMRVD916WoV2KwYOKE9ePNrA30KTKH+GolCJznEXgtg5PnBD6g8K4SnN
7XUxzfDXKRTDxtS0mocIslPdd7cvq1X/NNu3In2pw94jcQsVBTJgLjGYqx5ldch2
7MWBz36F0oBbkIwncw8E9L3jJukbgu/T9dtFFQiXgguoWTkRNmELiViVT54i8sWd
G/D0aT1+TFhtUvdS0jutOz4YyzJVCcOnCiXJJBYQKrPqR1NJzYIaTmrwxBQiEWWA
ZVWWHu3P8SeCmbC6fN9flKJ5JO9Go+dMKHPV44OEbuW2yNVJmJgrwSvBwYGQUSBK
i01Z0Zmdg+sVa+A3MkG8B5Yfi16avEPVGamqTkyBGqqFQVthjVy2rUyJqPr1hMnO
eZrlMRoZ4lPhfAs+/zsIyjNKz25mZNrPtpHJvg/bWWxee1uKoyiaJl0mY1/3PGzb
+krdQRkN7M70g38pSNLRj1u3am9LAYs+NDGOYHfaiYQjb8IQoFK0RS/vBqI3pn50
+o9AkBOqd57WvS+ZDP3Gh0EQ0B5iseorZNuk6hVXpBlPAy9vKgQ8BvTkU0DuAt8t
eshKHL2X3cXSrs3msS4N7bsoqJLCbCD6YebyRh9stOD2Myaw4vSLXqclbFZPEo8f
yOZLmrjiuyiv+MWQ2uE4AnhWb/DrKUhSnwmTaISEJHSLr8N7ZA5Zuqr7sBsVh17P
WuVg3wOY9nlSNhPl99rShopSO+B8945DIoAXQGmu7FsPVzWM9z3DTB2V8P0Rf8N2
fGM+WEG5BCyWnaDItlyWQJnvNOZaJlU6KnpEDRWfmlOmJIBNSh/bGLYhI07Ys00v
iVMRadvsxr1a9tGoctKiRXry6RNmF5ni57eLi+8GLo8t8U7ZJ84TKcl3nQe9EGD0
EEUtfX7oUSKA8WO3QaxHehDklXB+yVZrX4Cbo80bsL1zXAMVjIY74lHM8YSAQVfO
qDy1zqE2rYhXFs/3WQeT98DmSEBLg+ld3wTmmMmLkVCMLnpvbTmqXHE8OkCDcXos
C0KENvExTltnE7uJ5AX0tqZIZrDEFnqzfvDDBjOvGWMd1F3YztVJ/JgQi98M4RTr
2Aqh92hnkAnkSE1/b3x6oC8FEIPDGX7Ce3l5Hb9hmGQaXurUrqGLN3LbK66ul+9v
IzsGqJIgQIkDi4hu61i73jdGUPYZaFtU4mqgQohBZJPGkGulFWDXm47hnJ/TiGv0
fHT/baQlae7cpjGhAlmOBsd2Juy5JuB+MTowtPLkFhUcVyvF40AjWNQRicV14W8a
hLTRDCbDFy34TyWrd83Whc9xixpPDVqxQP2/yP9jKG98It0JfaVReUcWjEw5ShdO
X0k0if5DkWTPcSTJMTQfjKUD4LOtv0DT8i2TopEmUTwKMV7oz0twH9NUBsCanJzJ
r/9XBS4XkRw7nfyJtOkVviDN3IBswp6MaP06I3jFqLOnkf6gUkdo/grFqayNgTdx
tTQNg74RDkUFuH3aAE7vCxKBWv0q645JeBXey2crUIpBqUj18cArhmI9lNBWBMNS
mKsmxBfRciyLIEci8tUf7PyNiVpF8XO6SV5G8ii/kKmVqVQ8J8aPdTOHEfxS8CJu
JXr2KSafhg4QKYwA1uTvLJClKHVzn+stq/pnvbOtuNB0+FaDxZnUPhv342aCXtv+
HWYqHWxgBVCnVnTrWHLko/dsxeh1NX/BrojB/QJMuqecLQedlnTbG114efB/G0Ie
qks96v+Peicg14+9ilP9/Fl4H68BW/I/NSLQh9Y31otHkfnil0jTK7RYc1j5jEyP
UONn5W38pbcOSmcQutg6H+ggZP+SdYjMLdk8rITcADwe81LTj3y4TC7NMnt4YW3R
bTEEZX75q97VdXhPy6NuxBfeJGSLBgpE1XOChX63hdHiYgAgJzje8gwUyj8boUeE
3jETMPwxnpqppwIqQ9kNJTWZg3JrPrA5LvjFpLreg9a+naNhZSRH5gxPJTQlw7mb
D+60rYHosUEO+nNukJ3+N1XrZgnz4o2TgzJPH6JLTCQhm0uLVDICJlGXHduJZoIG
sq4odxSnCdBJOgo2pJFUrCbO1PsIwy1nTeYJ4eTHgi4xOsU1yee+agzkXz3zqzl0
Sk9kapLrsFakjTFTmP1vuI0OzJyiduB/N7TDvO3p5oXPCjehqP6hcNWZGJSp1xHe
rSNDmVHNk7sOSEl6XozyTpfJDrDasmoZCLQn5g8mzyPsgjC+Ip9loCHnJsf3DSWJ
EgGz4oTNoBJvTww2d7bIQYqMeCazLX0VatUpG2Bcy44p2X4yfrJTCePo9CWMHvwg
MfC6eodZRuBQ2954GmNrH0MNgtlpbXNR9e7jIy2pvZZZ2DZAjK+xMWNjdJlA6gPv
dSo+DvVYAmcDcz2eMwklM8ALM4wl4Iu87Li2K9nGcKVyoN7FZF+H7Pwfzds6Hoq7
Yq0viT0ygEoTGVwCWxcIcxwQDGCRW7G9NcWA5WaWa7zHhLBt0WE7JtIbI9m6eMfA
TtQW6fo/O09UvfUPLv1RrM1cA3WrEHG0A5qg3LmW7F0OCsx9PbgK7KRSaBz3nFdY
ujGbkAGVjntEgQyGji34q93wmnWe+j37/TWKGTVaCdyTJTGG6WUteAv8kV9dRIlb
F+gG4F6FniSgS597pxO6/vVbhKOO08XNvMzHLfrxzILHPteHdYscUvwvZk9ciGjv
ENqnvuY2x6j2HMuBagRs4afr/2TYcelHNhKJKcPOpOkaBRLf5A0WupnHsTvAQkPP
tRg+Zua/hN0iMx707rtdWttAinYUmZ18XBg7RBa8RIS7CTvVl8dz1yNlVnCKMvqH
OjxROXADEgiOThFjUge/E4Pfgmi3eRr6uK9qvgkg1Mu1nGLImBZfwOf3cYJ8+Ok2
kutix25bD/56poRHGP0ksJw4DvqiwLDyBO40XOdu6H3P0atKbGXopJp/PlIxEujC
MY+tAQ71rvIEfpsIcL4Va5jTa2HsJYmz7p2lK0YawMhPplz6ANtAYMIjL0th2py9
1tv+Y5CQgqZle485TK8/NUoeVdP+jcUE/Grgn6kt9A6bjRecYLjrnRMcVsRqmG2l
y7IamRkT1hD8DoctP2tDjeZ6bzGrrTdPnkKaHiLXMcU6K3dGTGxl22GQ5GmkGqgA
Gq4crjt91+5sfQejsyguCY9nx1C1tFE3wYFcrutA+Nx7y5gA680S3JkJmsUWJegN
0BGi8ofj/F2CT0n6056pesb130HcoORqR1NeqLgtHyjqdkMHTY2/7xKmq3T13dZQ
V2jL2SMaFdRx5nJ3oQ1xPej5+FpXvDq6D5C0fVb9HFoUhRgzlTpL/vabgGhc9tWM
U/YH1omWA510KCObfRehxcZsRAfjjDy78XBTtqKJYqX6LlaICtreMJ3IOc9mYjI6
Ms4xKdVKeCRe1J/Wq17YCM4FDTs2GXKnLUZvEu8NZHGa5mvMKAeRFCqfGIclA732
6WZ3rcTYZAqXZxLmMJDeVEO4PXXYiyuJ3cJvq7GpAIxJh3iWCCQqD0YM5C26N/TM
LMlrkf0HmsDQLzyeX4ympKfhkrCgb/g62RjFO9FECxHyrElHcYf04ZGVBxknQHiW
od5aWcB/Bz1Z2M+ET01t45lRpKdmqY5qqmetkU9iWHJIZivkCI3FVpYA9r8RyzCW
bHTAydMfCjoeJSU7KaF/++VDD6FW8c5TEa6GAmxDM62PMNfd/CgJollWbMQ8CFDV
WXVtomfGCtJ4IDaaeICAHlJiHJHV0ljmfmgWwjl7kYV4ApMndquWD4TJfaTRp9Nt
ZIFDr5LCxXDWS/bwoxd0dhlY50oVaVw42h1m/yBSkZBY7xtAsWS8eI2Bt53vT5MK
yun8iF/YOMfEwuMJIv2zmmKjZYTT6C7kisWoE6WszK3wPx9xIAN+Gc29Uix1QJ0w
CLz9k8Mhva7LiVEAMkN3D99V4J4gSr/1wX1zdR8YMhmmT+b6CHfgZ4jYKqRvQpqO
/eqgYNeNyhCBo7dqHOzipNHiS3SMkNbUVcmDCEV81W0yNhcvIWgNuntb8qpBnnmK
KOjOlx33LjDSuftTryHxL8U2rrkPOnzNX5UK/xg/rliM5PuEa0JF/9w7GiQQJfxX
MNAcf3SpFuQvqBHdXPX4oL+wKg9LkobpKiCIhTjS1jdk5495xHEy9hFoLV0IxgZd
+74ekB5RFwFXojzTB0lcZhd3cfoN79SoQI6gfPB9WWGYyZt7SFmR55xcdT6eVnUh
wVTWqJd519wTGeb/5yd16alGMeqqAFzQKS0HfAiWrmKXKIQZ5iHtbdxsrPmygdG+
NFNE2c4ODstYnI4KJF6eS7SFAu62GNcaNEngPxIiqSNd6pPPaYuus6avobry2ZF3
PuYzmZ/Wpb7BEnQUqBRLlOVRDBneJRKTCeGbGpuDsdaM5OqPkaKEJEiW/GwEw/TU
MRecA7R68P8fSgtN9iJ5Y8RAsINQYisOa2zDxwdcwJlBtVSy0htiWLtNozR0t74P
hBLf6iWtkuBVO3pVR7YuvMzgA1dRIf6AmdDWYEd0D/hIWE9Q+3gKQuA7O25FxCCO
CQodhcVC5JjLepFxhVn585OVfPFeZijADQk7NpYqsgFvlM6mIH763+0ndWvxy1Fm
OVYOd76DuaqyfDDWpUPnL6gGhGeNdP6EW0eZ1c/FJsbooiiqxXj9BrEDr/rBFG2v
K8o0cnBxvkwv7ZNRy34Phz+sbUc1Ljxf97JlWdOQM9Mo6Vk/oBo84fsWmBJvwyNm
rKSL/UHrKJ7sRGhzb0EgO/nw+6oz55Afo8qwr4oRIvQUVyD+L48IiwqlJdoWrtOp
NcSGcBbop17+NNOHM0RlApHvUJReGSlQKfRIPrviMSeECwQ+YAxpLlySt0kzIMuW
JHNeIo2g8Xb0viOTinu4e2JURjymJu6+sv2PYKyCjC1fMTuvzHNIh3GBdaSZckN1
isBB2Q2hXwhAKhhqqhifz8BR+CowH0KoOyBDx2SC3616qeQZGH40wYTZJXaazjN9
xItYl8N9I0cF3rszC+oivkRtAWxy0ZUw0+cL8aF0iqAiZKynIrHM7sFAZJNp4iLF
5JcfIC2dP8U5C8e3dTH0E3PgOvAbKFfUJPJe2TeqRbnVvTjGlBjJKiArve1qLR3W
7eHCWdDsmV1F19buFLBkL7OtteFtYVMpTJZAqEf3lVFgpOJOHJGL1w4oeEZ4uoZk
cJTg8lEewYTBXPHxRdmaDWciFVkXWGFbksz/g3VR55s//zyDLh84Sy5Nd4rmKLek
uFltzMuhnC8687yKJBz0bMscilFrpKd5MAfybe5CMXfG5a8eLiGPQus+yWBlsZ1k
PCc/rR+A0u6CCWWa7QmapaApQE15e5sPiB5k7Dvl8U8VsJ9GidKyGPlHPCV9ZgtV
kCHOBIj5/hQWhU5oHrA8jng2TuIYoO4A1AX+PHAqv36wp+gx4EO2Pob+0ULgFqi1
LIaDbod9oHh0GfMdJQTtYyEPdlnAmjkPtKqOVZZL8XCB2DDL95eayxUIf8/CVJbV
4kFNccDtuF4kX+LcNU3o+aI8CD49u4eX5fVSHWst2x8/LDXoBHU1ZzKSEtGEMFM8
42KFV2feObr5jBuCtb1Bvk5LQiDqaldSI48LatQ34cYE2l5P51ZQLC4x7yRzlxE9
16UkhdNEhMB7bQGyDWC2BLNIQogFi9yjicxMTCRtCPJGpiJ21xZ6Kfw7KHvnV3f4
vOo9eEvEWrdhW01R4tkwjYXvupmk2Am+ykiLhYwdFL4qD0kZ2GubHWwANx2NioQr
HO9fCJULX5RC7xnWnXs28bHfOB2y8gXOB1ZOWNZtrnL9omp48vq94ejvY40Sm4dj
URQH1ROU8uyFtxD2k/jNfOQlgcmy9rK2gVlNIBazIIXAjl0f52k+pDAwSqO6aJAy
NlASd+YIRS0MpF9xg/zvzxms9rORaPus+3/QiU3hVAzoO8DviaCgg3JN4vDOsGh5
2vMehlF/Z0WWW5xcI8KOFmaB2vARRQ4IOYiLLZLykPgnoI5Oej8QrkJOxGmBz8kx
5D1K3RiFu+a4cwmT0Lmoewn+AMVL6twiXreWEDrAaLnTLmXOePWPARGPjwbk3Hd2
yCClOpRBpRkgj7I7b0MzdqC+fm7zWSSx0sto1o0uBt1mSYVqiYwuNMVaIaohpyRt
Skumbf4sBsImjBS13xJMRuUiVxsjje2k+/Dda8piwhbn8O9zQre8t96hOX75IAPZ
t5qZ5dQqN9dlk7uhtQZhyt8EYqXqLyCidyJMyWLwBTb1BfCXDjNorpLC8x9VAVeV
zPFKxjo6jIdx5OhAlkRLWwLOlCYt2TyRoJ/bRrBKxDGMn27OSJkpcyrgtUtYKQ7+
tjIGePIaZS8dOVYhABZtzZrpOJi439oPNreP/TXcoLJsElLhoa9yBNX0rZQ8Td1j
vu+kixPKrtrQZuk2RYYXuL/qoua0MJOSEPfNRWqTz5340URUytMoF4xg1Z7D6Ysj
p+kfKNiErCsTSUvvnFw20Q22ld/C99dLUCwHoYig4o6PlxGqLBJoJHp8z9H++EQr
vs1iDl/aY5C5kLB4rAj7twFp9/CoYxtNqyt/km6p4tQmjdMH9f0HETmOBml6iEMP
LGxGvGhO2HmFA3gTLI0yVDEOXZIbpJrWhZPeNCeMVi2yCyXn0gBVCUoVBw6TspAb
FNIe3qyi196/rL9EtbBVkQMa16bvN3F9tWfZyvkBOWGVlmCGEgt1JtbeeXCgeWak
5DTVyFK++PrO019wI7cYG8ks2akNG0L9IWWaQkafoSd7QT+RL6Et3dt3JEksyx+f
INGt3QOW3xL2fx8D8yf0HDEfwd0RznufwDJZTKAmZR2TNlt4aUS/dlNaQkkojQKq
EId1gfuXH36r+eji9SnGh/mSHD/ZF5BJPuwGDieIhrPHjMjaWWznQs7l8N+WdJl6
sRNcCnxhcj2BQ/Q9Y3h13BsAbP6YjvNbLFeobJ7yn9AIsaAqHDRUdQ1oIWc6aBkZ
opgywbdzsTS6FgnACeOlFY07dnJEkxYv3xC0Dm21dUh+XXzKmvebMtdgnEndLWd7
ZzJQpRGTgs3WzbX92JXk3tVP4pTEvdV+jogsAOcmv9LAQh4txTG69LFlnmWzVoYn
E0GR+sVFLaM+gdpSWZyWZ2gQN6FJP8DzePRbZpAdyWk4O2kYZJxm4kuuaeW8sVY6
y5vXpxEqbxenn0lOuMg1mx10q3rF2A+vo5BNwLYMfSnQkqRdN7CQj8CfYYWpB50A
R+CnFWuOIAhXHWqHJ3mH8kvo0aKrgm2hNituCBVKIBlaJ7hS87E0dvJ7vzDPUDnO
KbdF9gf3gjs+RCzD5CMxISUvSRV9ukCue3CcxEqgiS0dOjJ/0b2+mJohH3Luk+v+
f+uidV0CDNpL3m0mT8GWQhSt1+En4fUHeoVRrs1f7BJm2ZOs0g/oeVVtxP1rQDqG
z82y2FcKMuy6utGxwBIomGXRaNJ/HJ1SXA0f4KFZ/xExdu56fOcz7r/BobyDQJCF
OQBU14EpxH16UNqO/qfvyiUhSgj676eUSCALjTFgxnKzm6WXov/TL+IFABVSQjgQ
KWTOYIMGlC47yfaAKycMro7acHYUKncv3gBCkTtGFtOXRL1f7Bg7uoQ0T51Pu5Hy
eigHQkDYcO97l5GCgCtKZ4kd3jsKPYX9oyLfOKG+6gVsuqBIEIY/3shoD/1VYSQt
ih+Clr/JfllQRiTEzCn+86B3ueM63q5c3neTJcSzytJD1Gu9L6DXKIpjnAd5udvr
fvuAnUHhDu7xrrajdlNobTkKQznXobUReIluJEcyTHpdDJvxoLNrwQG0BoMd3avi
E9BwY4Fc+zIfFVJdxQI9U/HZ+xHnmknfycXk8VTDIUNAftqjZIL0OfWWDQ+pmT0J
Kuo04Y4c72QQAVym45iJp23nUONdgPGslX61KhiQtoI4qmaKbol8zc7Axsd/btEe
WC+aep2jgtPzM1C8dCwrw3G4K99MAzirSnxwo/cRM3dvid2N4ryU+Vo7nFLKR36Z
XBqgyo6wJUVNB741FZSwR/0Oh24JnqWx2XY3oL/K7QfOPoiqayjPSRzTX4F4nppV
3lqbzESioF67x0ZTisFrBM5dmW5huHOpMO+gHTuc0TDLCTY+ByGxhNQWCnc1JqT/
An7JUDnFfXWaC/thOtRv1aX8OloAG9WAzISCjg7V4rndYu8yQlwM3BPb2tXNVFj+
rrqMToAC22SbLHUakQaH0e28FD5OcPr7Deh5uYTS7cCsapJUzItoJYsEydmUx5G5
SMymVA6XVbyDaKjOqQ2UUXhzYhWx78I7IvpzuFm7QqgkHaw5LcYi0dhWDO8Mfx00
jQ48N7046TjfAmP5t+rQASZAXeIpypYViZAYSIRqu28I5t/2wHn+O6Swvcj3HvZu
d7xvnqUwEyr/v6l1JBgr7ZHIsnyijvYK6+pIJ0y+XSyqB3K4Kn8ruS3WkG9OgAAr
p5BuxPvtxq+O5XzPUr6PxOpg3dY7rbtrsGeQGr79nNruhgKrws1yXOjY3M3uhv5H
Ap2IxsUYoGAAXKAtBRCmZIPodOMf96w27W8JkBtv8wdY5wlxfv4bRM2vUVqxjmF1
goWuxqZtz2qjDzpHSupBeTDeG/kX3RZz9A0jwsosKEAYyiQMelW3Dnq6JaeuVsgH
0rp5DXecQRMMY3xVkj/e321pq9p5QEOAaExKcbz6BaCE8ENHCAQ+ufEDXB/HCnVW
XenQ2sRT0XDnnQC0DLOK7bDtFTzv4T2smEwkql5gfxn0dmIUdP5nxMm9hyA/SVv+
XvdBt2rvsfGcuhdQzvaUZ7NTYMsMDfek3pZFg3xlqST5FJkrAc/fiS0dvqSQvCsg
I452Bc3ZU82nWQi51BM9pK9WnDaZ33Em5M54/7YuDpswBa7cQ5up03GEhbc0isNJ
V6wh2/NWOjFcK5HluHP6uk9BE1R2q6YzDBmkijojdkWdS2556Fj1GxL7snJ3Ppu5
93RBevuWs28rKdn35h06mvggF1vIsfF3w46lXRTqItSh7Z3VfAeKRkP63y5aqQWi
rdJJDkMIXxPH3U7UtduhIGEWQLUMtLGAyzwPfOOfMwKRH3S9qb3t2cIqeqYirHFA
+YulgJNjVjhCkieDZ6hC4Hx1wOm7HRlg/Gmgyjpni4yia7Ftzx8zbttcD1s3urIr
Qcywp249PSidN2EBIAaGwtnE3q93xVePfFK41nCX9oa7rnxiswizySES+DodTtV5
k59qtIAMhuxlZfggnlGYcMspjA5JyHFu+WO0p8y1cKuwuKyoaxonJSe5hSPiQbHI
qKUQ1ghcfAYpZiCP3JJj9lIm39aWojpZ8sAb0gLm+9yZYBG/Q/bao4QFMXzNSvMf
cDSRaK0tQh9+E+X7sslOMJgTwDqObzN0RP/TNvGRbgFhMYsvBQPcqy+TYzJ4i+va
cZosqD0FZ5HztawaTvYXJFnxpb2fZkrZA+ZcTcmxGKSRX7UxPM6iUdav4E9sDxmo
C65+p0+dOVt3tZ9o5GzoRhyovI7chhsMaoAMMy3AZFYPV1Aej8hIt114xLSqPViw
NugY5fbaoyofG0hMqdRM2upCDDe2fTc4L56OVC5ek+yJYiQAcbpf3xsWL2BTzLfi
ycQEvCszfPJNY158l3W69Gi39uh2dmWJJvE4cwCnDhLAZdylDvehbTBIScRWlCI2
4cNcyoPqQRjoHuvXRWTq3ZMK7vQtnq4h33gxSYZ5Izy28uohJBCIPLLtUtKAN+vQ
Ynsq5O736mfKDBdUyk7uEuvv6NtD1HU5bqcGdN0vjD/r0Y5vcjGxMNAEE5vs7eCc
r5KZ9v1n7uEbJ76YagXOFM271p9meMAb+6CgJ4Yhk8+ljyJfMegjf4pYhI5tmks/
RCGCjkiM0jYGwz5yz2Fi1u3Opf/pxhR96ogmsPveYeCpAMwAPA6LjgKKbDJYFJFJ
TvxUOKfup8yTkziWiAdoGfcbZyAOCYx+AUvQ+YLW5k5d0ewZHoNYM7mk3CWdfcOD
IfzcJ+S1KM9ZFEY7Ls+hxyMSeiNjGLwwfyIopxnSzNr9xZBmeG3022dWl+cDuGq0
OcKesJQIcJDttl+gJHzxjVJ07xsMtWAbRpwQezyXNjrAhQUGzwtwop4kV03caYaU
DNM5PRbiDMdEftwSnpGPXavYNTfwFXLIJwcbRvXLpe8M2K8BASePJg4u400gAkNd
5o1j0waXu3QtI2iJWUxg9RUlCdkDRNKMaEUzldE/3ZXth6uWrXmG8bYt5+b2BlqK
Q7II0zqelzwY2odlIkq47yZ8r3rQLt1dAJthCPaOsNMTzpn2rdOH+lGAyr8D6F56
Q4qVTM5Bfqy4y6ENATI95VWe2gYU9/5Pc7MKH4fHjF5PzfOEIylSQ+ZFHVO1ymjW
Flj1wJ1pYw+jCGTmE8zSeInK/Y1owplgQk9Ok3geQM486fZtpoK2qE2xcDwuwJ3c
37RfJDFXRkK5Vw22etpCxFyAFBlszYmVCijtPhaPlaX40R3HrZQnNv8h/5AeQ/S7
TSx/zZHoWcTY1Yn6mX1YCYdAwzhcB2ajvVB6MJXEaWD04JL3/IGGGBSIZ4ZHns/+
juoZ+nvGwBc1UuMhIi07s1T1e17nkQhWsdtnLUJC+4/ULsdOTdSCB79UNK8WUcb6
UjoWRM+cZ/Av6N3Y9tydV6qjijIOnSHIF0wY80hDlTR0eFY2QW5M8PqTaLfcMopR
fAjrBPQ2Ua3+8GhV9DcGDaF5w0ZvZ+K5zvHi/lDL9IRh9NPgVSOo2f48NQ0L00yr
GSz6opPiTlK2tcTwc0IW0zfzCrHCsnhLqcL0zA0HvDNdEEYv7ojtNiF1gDDMIsLL
bi5KoOmOjNJTZzRtXM+5mTuFGK143dFLCg2iC4JSg9htQedSZfWzGvIhps4ifuz/
Cl2j1bADe0gfs3VMfd4QOTXXxUH+/H9JiJPJNtv++ci43oSdgKC+ehSTW9ZQtA//
s6qNq1vNaHWSKcGk7V5nQwnznrVaB0LBwcBWS9xEY6+VD7IvN3DstYxOigcdz2Il
81tRqp9sb9R1ShNmyFM8qJdxBNIw11cUE1ilF2UuOLkvnTR9TrXG9ze6KMAtKQM6
KsIyC6g9T2ob4DoEJ71H4yrfvSAak/cP3WnOS4kZ/gs2XkpJe2Jx98+4HEqFe2FL
IJt38mGtJcEWNRGNENtNJFR2R+r7gyZRSOCAM882NU0FyZhZRAu6PguXxVuJ7lh4
AI4FY3flinT774w5sEeEFFxOWsl383h20TUR4Sx3zRjZJ+2VgdOP/ZIVtBFGYBO2
/LiLWkMPOAixUm9yj4ZuupqUe3OidOjQplu1cOIxAi23ULO1WfWahcupPaD9Gvzu
Nj/nEzR8z/tJPn2o4yjGiAnbn+ECSaQJuE4GMotEUVfhw74ajtI19xxXz6jKCE9V
O0B91tNNnAejtt35yp6c+dmR3pU9Jp9edxxC3Yrfw8dS1mL6D1WF/r0V0JiYjaUP
DHg/j3cNmirm2TmNm5Oh0lvtkqIgwlvblZxFvZg16dv0KcvVem6CkpxwBSSKHzSi
wUPSoLzObi8F9vPT6/oZio03/HW5Hj9rrAPYOZt+4Ep+qYpfYIZ5r2v09xbeJJzV
iI4I0tlaBuE33NPIYkOp3fs2KJfzBuxRoEaFqcP+gK1RdXX9PoZy+jhGevjXTZXE
SYz/HrD/K6gy95H0F7RaBTv7f6HizT3aZBVh89DE71wifdFO6vWqsvDxxVFpEzTk
MmtEqo9vrFLv34rBlSmm6E/txshANo4Oi7IW3O6Ik9RPEo11H8RsW06xcd2Riili
WPRHH+MCXkygyv3SOuvGXyoMYBSw40hDOBuCUsIayjrDrjz9byHY9xLlRscJ9opz
Z8T+c4SFCBxBrCsrThAe7qQZKXdskEm7SLTvStxcDfMFZ+Ut+n/9oM082cCYtIdb
wWqjJOPvP/MCkWL61nC9oGAoj5NYfRtU5ly0Oqy0jzfXbo+nJW1XkV7Eb2y3s2vb
2iOc49AzwKpg/EKpWt+hbqR4DyxArURIreD3+Sbs9vKYQrXljieEMMqvrUZA2ALi
GWs5mvyFGT8aLyaZ1/ziMB33JJLQcr6RIklXygWt/0SPlK7EbcIdPFmWfGq2VnC7
iLXJBG1AfAdOgTsofsVz9qPrGjXP7RzWQLPt9MJo/RAWMRYedISbRwQxSKM3VZWg
iZ7I55bvMRLhEEY0epPmMr008Z+Q7KdYoWfMSgqp01xmN1wzA/xX9lzKq7l3wed7
brX0pjhZbkovWsc8MOokK54+61d6w4nJPw7+GVWIHEySfKPLIfNi7zi6azs3pmeP
hBJWda/qrrHi2VnWl3pRF6PpPvGHbZuqW2POOc+iP2gZde1OW0oiAGrpisZPRGAe
othBg2PG5sC1Q75/zK2v11OjNaF40H6Q5r3clc2DLE+fH3xTG7pDNVIBhQ6/4swg
wb0deBe7fQSfrvodmtjHbE7yqoPERGqRsuyIhKHbyoy1kCRJZegYeDgva2gWlARl
3yibSECfVqg1hdD6j4kyibStgOq/lh6yoCwIOz5c1raLIQaCO1mN+E1+Dhuc9S+s
CyfJNS7TUOmtKvRPYo8nOxd23PPok5jSSKLvbLk64V9HZwwi5zNYFiv/m1PAEcBb
Mzd/0XRrGS1W+eHuXjUBsRcgPXCzfGkR3aGNRyi6k9/2ZQA2VoHMdPqJUCkuPApj
tuAjnmzEZwidO+JHFLEaUyexgHM2c7KDxu25NVKQZCdz+ylDR99XukGOjsYMLv55
dKyfYcV9uEi/gd8Zzpus7cwSie/20/yeHBJqJMTRzcrhQewVzKw9AYpTlQXXaUAr
/+3s/2OKCkv6ude8OGYfEluwqx4iQUN+1EqX7BcpNmVWZIiBzJOz53kqpr0BZEBT
Vyk1WFJItAiPnWFtoF/5XUVd+uXwUZamWqxX1FtLsO9uRm1LNwLLZgcIgs/8i2kj
NnRDNDf/T4+8N3hzmVU+3N38N9RLmtt2N+5wnzJUD8o5Ig/826/Fh9YQk3/y7zFz
SPYDNyZbGUkHK545U564TnCJwosk9jppIXj86EPYI7I9v4tJDkFRpdE6YY5ntY8C
7ITEoflNhCg0gu02396QFNVOfW47xcau3AHL73eHZxs7g+auxbjWbSKWJAECIguF
HtNPBXDNz1t+4bCqSA4GdyR6xpB9DrnHsljFtLMpPMWsgXZM632VK18oBhhxk/g4
iAgMfRDfhydYF1DYEPpyuVu/LwBELOBLCsaiiD7irb7gqAMDLj7PgsFDb4kfN/jQ
vh5PAwr/JH6jb0SQmQoyYC+3Sw2ZRPF9fvsX4Rn1JR7W2DoDNOU5/gNPYExjwpgA
2oWigTBRGm0NCNPYLrHzPdX9dBtIvwVrdHPr/9Y8dMlVha1CdjJ3vkkX7CHovifn
beULJ96Uro9RVJVc75HCXvypxDytfLiIPnxYAYEhrFJKg7uOSKZ6I61e1DdF0R0l
CSJZBGZGlXhhkWbW+tm8OdZdfNJm7lwkiXEm1IXKgoT+dPhlkLA7jJOYFI0gQqvi
0oyDikxUM/8lX8cWpZ5wsuc9Ah4bajPFT1+TBP1zWgY45TcW9pcOa9NJnf8/JfH5
U+j/i6Y/8UaJd+qcdvix6rNyk3CcOb9H7z1Q2C170TJ2eT1K6lYd57wDA9kVoM7F
Ysaz4kCOgvaXUef+3BQVtttv5tTxHNn08dl1mZt6/hF0YRzlQNOwNNhsz+BTmvL+
mvtsYAGFrAecMVl/3RP7F8xxh4J07gtWfkdPJg+HqOWhmMAO+9VnOYGX6gkoprRU
1j2l1G+ZRpZk9grDNps5aVugW/w45fnIOUzl3UFVMN/PSUVNocGlTFtErtadoiFY
qttMoo8yCxnDIAQwv4rgu2jS06YBn70zI5ivkVHu9h1eC2cTPoRo/xgeQ+HEmPRw
nfJqZbGJ+1hLvENtMgz+ov6XXg4WrKwZmdiXQnJX0gQhNMC7NTw6WCUjTYiODjim
pqg3I5UnCLUQ2/Kpow+ETbd9bOB+EsFGOfDTEbPSdkvqDbh4WpuuxmQlpedcX14Y
7bh6UJbPHMzBTiw7YMzhJwLjICcF+JDKppZhFJGu1aifdWNy3GfjA7GUSQdga98J
hi5bHPeNBcMKsfcJGOdiJpNLsjjLw2zK+1E7GkWR2uqEI6Uz4KNQ/yC7w/U2YHky
yk4kTh/y29WcLtVAwISsPETWxmUDDhLZYHiczE+16IfiZdoGS7yfkMdh+oj0eg94
+kJCP0hr8Efz+9NQnK5j8qPJVAQ60fljJjYrnH9kjSxCM7bPhw9vEuEWVTOMnzoU
A39drQSNtZdxsTKPShj43ITAsf/fGUO3aXdsaaHvAvXnPp8bOsN/KMiAewGAI7JO
4huwTCi7lRxF67a0pJLTD4QcmiYCDYki79tI+9r4/dr+owpH+SE0eBOJ9dd77PhR
YJfGwdOo9Skm5VDDoCET0GNA6kBAt+NjEP2XlmfFgv7e/xktcg/5Y0VyU6hu3szl
G65kAi03bIJrZQ/Q/ZSQ61y/7ff7IOM10xvDSL1lsA0fCD6WMh98elIe/+WMu1al
5QHVn1vBBeoL90lDJ4LFyPNGDtrtt7CEDKA5j/ZNXwEe+/CmwnESo45coN8dYFbx
1/GZecDWmqhDhyePYl4RUJmE5pboVSNjleyropNSLNyWA9lCvZt45lKi94PY6nF6
eXuA9TghNpKPdQAv8nYoReuN6S8q1tZ4ge5u/DH5y6pXQd/cncu0p0D9QKJwtT4d
rn7dDKGcg2MWgcGjC940Kfnt2t6LQYRoeYxeUI02h1cEwA5t+zkgD2hbkbqRO5PO
uxQIwhK6WEXSXmPaMmly3civ5jYRR3ZlKlwP6z3PzzMbn3CshT8CAaaA62YS2sGV
d2D6z8D9pQEZzK1XqXjkS+vrzSpQXZqn7d0qEAD5CFVxiHf+2lgOGeteE0cbXiMv
EN6cHlf0rCs6oFFQ8b6xSYfdbRu5RxiA6+HOxcXWvR15p7WZ43ZHLvlxje17urfS
qPgl7mZblV53dsXlvrTQw/hB6tTY1aV1QpMPb/8Fz8YVeyszccx9dbxqYKJmfH+s
oZTju1oiaLNkKGPRSUS5lTUhbRvCVw4rxucRCx5EzvmkEc9i6aG+3IpXwt8tnOR5
P4Hn5PYTpq+OoqtJA/EWF31zDDa38/aqQD/sHh7T+0J7lsYsPCwd8CwWxsJSzV5v
5EnC1Vsd6qSnsgcTR5FU2TpYTiUGgw2iey0DZX6YEk8ee2BN4O9/34+/D+w8fmIb
n06EPUIOen/RTYxu2WXyv9EqwDZVRgQztsE+8yhkv4Fnt6RZLjDt3gmiwcd3fVMh
88DqEpfitMB7P8Y0gwASPfpvyw6DPc6HNCVwCPjloitrBYQjPFNq1sZH2O29vggD
t/ghxapTkNVjXFYIA3cPZb9nAL3xCfZcqODZrEWuW54rWwxDrITeU5DFbcTbY75t
8Efy9v8Wkzex6O1e2FwTdFpaLXGoVPPxpk5j88Yw4UPr73j4uJTNpgg6hfeDORFj
vYdrlxBpIbOZ2kw0cIrclPo9ZVilsuaDNb53ZVFjxh9MGA9E9oJYN4b2fpJ7uaYk
Z12JGl3QbLV3kk4K9cYIXqoxn4qjk1dll0cXNCVl27JfnMSTPxt4fyQ8BIaXeB7d
g+5ALRXWj3p+NMlQYf4yRAY/SBS5zBSbt3P5aV8A3QVBirx+m8WQkZ+6isrRQYGz
kqt7AdbLF7LyNEPNcN8FZAJrGueimI5nbzl01vcz3bXSFZAKt+yv2kNiYuulVR9Y
4PIxbMsCGbk3bKZhCVU4bWbqRuYQeDAB76PcXv3NuqMeOnn8k/EmzS7gvZT8aP/f
VPHfGAKWk4sD910eXQj+Ad6aXsLliObXTt/0baPHCHUZvCge2jS2vJ+zOQbycgi6
zO4uhGkm1mVMIFyKsllPD3OMy3+GVPkf+RQSoPZnvnmc4fNzHrGxMBZViBRqumCi
i6FN4OGbP5teaXSd7BkZde0tjA+Y2d6VSolieFwuhPSuKa2yXOPszLZD968wU3re
yaBSc338Wa2RQl7u12oo/QZPpESWEDaJs2G+d7IGkl/TT7kFcOxOS15t4ly1F4uK
Sx2RE0Q/UQyLYtgnEUGHPLhXPF1/C8L91AYIZa95F9gC7CVnESfryuCcIFX6Pin0
9S2af47fuMeQdRIT/DWnlGDxBQ5dH29xL3uxQAqbnn+VwRSwv6e6MsWKVpN+rX/2
UhOqYIumhIpjyO0C/9Uhc3vJop1WvKnBIFq8HDaIdpQqYTeocKqjnfY7XFU2PF8v
8aK9IbTff/j3A/H/v8pXQjmuc/8qpW+KyQQKeBp11eY2f7V9Ouw32oOh6JmquCl5
PYJsKO10p1n0jx7boaacb3kwUn7S1Svy4I8b7F5TGoIOg/iyryImi2y9DBgfJCA+
csvwJwXuwBtGKp8j+HsO5+1Ce4SKUe28FYbJGwe/Ky6gl5GSvaejhPa/+DfnpiaV
bWbiSY8ftr6J8IeIh+KyICWkUviafx/9h9bsd3fJpfXanrIIqZZGIL5pzgoUUMe3
iKWWEK8qfYFGh3kcrC4VkXCJNiBE6EUzqOTUzBEIRBFZP2JwI0URSAH4DqmZvFAz
ixo+gxMgPWLPY/XwmJZy9NLhy6Zr7sD/KprisxQAfiURSaDsBZ1RuMF8Q7Nnjdyz
f8dIOiqJXqSfbFDzSMtzuyIl+Rx+1MdOePZ3NwVdysrP1QGbobl0K/MNabDI+5Nb
AcQvVZzC97m81YAV1DVB3DXB6Yl4K/MCUj+AZE79Kn0nLCpb6fDcMwN+ch5s0Qbg
Rrt8TRBznjZ7MeEHtHMqu4IUJpUPlmpB733QIYQpxGngoUzapSCzo3TmKbtjQrAs
8tQx3ah3q9RHpIiue0sJIECYqjFWvEYAKyWJWnhQVuEBRW+XZlAp6BGRGDL+okLq
fC0lERbK1/8aPo/+BMsTuvWbnkueT7KEcu5xjo4LXQ6pJxM1KBYbnfSKfq53zL6I
AQtQZShypiB65q+dKAiqffB71REi+OTOaqIlruCqwsf4Zep+fIW+bRcdPbOziJLI
35xwNTwRHrCBGfKAPtSX8qnWF1sNCOyUlzs7H+vuq2UwaU93M3Rl+cbAbkABSerw
Vi0Nus1KeF1QODvEbItoYczvY7zRDTNQR5dLk1Xvj8cMsRcpxctLw9Uor+aSTHYb
18ui7fhvSbeViXHlrI9rfAndmANEqDClCIFd9mTLTxGTPk/Q421p5sz6nQONUNgZ
KCxcemvtBvmISsLkDNhG52mNYQiVM4bLWBNoeuhJ3A2E2ATyIo+Y9aQ9S2i8t58I
Z4M8xrsRxKEAEYdIq9pJbJ1386kxp2dJQPAL5XyAgLev1F13WfFHrEhHFGPq6uRM
hbUfL5Wks/COxgmvP2FAKVokox/ukBsYADSXle3qtN7X9Ordws9dXe7Q6O819Ttf
XlpTeD8n7yG9Be5W333eBlVGvmJ8+G+o2OMdZ6WBxhYn/vUuWCWw9ooPf7iwp2MY
TeX+Uw7wbO6ijB5NjW1ANnm1PgP4YisA7kPFWJX/Ly4HJ7Kz4VKI65Lo6F+RvNhA
o/pp1pdzlRec69sJSIjtYcf3n7eNP/0sDT3cqaOtDyUXs5gOgnZGD/hzj9RLll9/
QADLwB1u/+NF+LDbtMyEwV3gInn+gOOL/UnwTkm9LBLai2Ft+QVdS+ZRNjslfiVC
BMjhcD11MICOWpqPOtkjcQXamFrJg894oTuPE8sKsriDVTw+FZIS6emWWhHMslCp
cjYSN53QZYEmwtE+YMlX+eISkIi/vDnKDkEmL/WC4g3NphMcDeJyAaRu+vPQGtLp
QFedHdMd+1zt2TTgJbu7hCNoGtupiuxHg+eC8NBW0SnjsQT7mtxvHQHVD43QQPAi
KFU3CjWQo3HMM+HuB59zBBuUKzx8a+6ZJBjipvKSK7o2uZdGkAPhx43WxYJ7aHL2
4C7EgNY6eamGLYPvHwukOuMI+WcjC0Oz9DRqh+cGaxg46j+kio9UkzFN/bjq1s+2
9zOaiTmHKtDIfsz0o4mjxiXaGx3ZGvmUUMGydMh27d/2+1l+ye8gjaX0P3Li5xfD
3FqcQOHzUTcBXXnypX05bO1vZhNEB4OzH3Osy7J+TYR+6uJuvyFaZaIwMoCF78sm
OWgInC0RKb9RuTqOPMfccKamXzfzWJQgcg26FsqxBPHSf5ZAedeoGYLW60Nn2ax7
rg3FD/Qbr04gmIwEPkGSxySQKYMRWCB1ZF54lCu8Kh08rtx5/iuLf91QzxBsE5l2
Z8RgzFUPs0CuZq/DELtPe2j9cmgOcrv42RuJfdBRi1PQ2KnOv0UWhMU4D/A4xnXV
LLRDZEdThA8gKsAsZM8BkRsHwIhZBaajT6kLPs2rdadHto/Mm9RQRIkUEMHB6ICa
5W5GyiVNCtWJCYUfl4NkGlhIqANtCcnRn+0KfUBi7KZgjjRKpai2yNwOEUITrc4D
dj12RYGNGzztVv/FUUZKtEh8zkJK8fcVohUSqxqrqCiGPE3TgqTyKx2AzpJQSlpv
N3EnrBiePmWeRT05hikrhw0WqAACFFWLMgu/uL6I5HBaHi2DaJ+UGdkBVf5z1BR2
WCza/lQkpNx2tiEIMWXdxtec557MvinhiM2ViBowr6xNQMVx9QDvuU7GIZAoEjvV
IsEKk0V8t+oCDR8sP6gVrXGtSZKG/v10RvzeV01PcwiLjXtBYF/CgZ+lDSiiyROe
RtgxRB+rt2t57vaRvaAQR0lc8J+Nywpv1RIriolbEuopFbS+g2QwaVPh15aarX1O
Aht4/zFBoJbsse2EgWM1DLZJ11n1pi5N6XyXzifDVLDgBGZdNIwgL6K+kq61u6gI
Ku+OtwcNaqefjFvnhwKPSjpIKYTFzT8x4fdnLS/9Wb5PdkN4aoiCoxZW3IA9flKC
CEGkbmww6863EnenSKySJUleF4XoXaH/vrY8vBIolyZR1Eiq37i5zJGny5ApNqmT
AQ1YeTWT/84e0OeVkRbLlszhPrhazp0slt9BXO1CoiuXtHU1w7as+z3xJ/1A5snV
J063Su45abvk3V9KGIk523bGzT1oK4bOVpUfP8oGCItjjGZXNSWRqA/uzvUUJRIC
hGOFMVmCxXlyM7gQmMqvffFrEAzXgAglw5i4Mvpgiy7DPUdygl50msRwJU05HR13
9UYGDcBePRfr9bjtE39pmaOQtMAwpJ+sya7E4a1fmMPrY6A9ZEqam3Z5WGknhYFr
pnB90ujhwNrequjLHdR6SoDALN9mZvtbag1Mwvk8IGSgXUtEblurotvMtOjLMY8j
nGa+4V3leTYs0vGeAaUYWJhzbXkEpb0ovrozWEBYdO+DLVjPEKfyxw4X1rtBMx2p
7etq1FIP/uEfDOdDZPJh6zi/CpeGbeueiPEURNqhnmRXYHQttXaft7olDg5poILR
MhunQu0khdfArQGqxDqfWDKexY4n+J/mYPGKOUMHjk8CZHJCwrSi2QuAGL75vK+L
wY02MdeMDnWPuXVUJy4PdkXeUkKSgHBFAM56y/9kJfAtlly5InNUCe1DjYvF6P/I
lmgPa2Csbovrtfko7voQchFPUBD/GlolEWDFOdHK97MI8zrPmiHcRQC3a7jYvij5
njU9yHuDZru7ln+ppr7uHIiErFsxKmeyjyo1KhiWiXMaO47P63pB65TFilycCj0c
beHxYZtWGmNUNGhT9jCyCLh/A70MMEhg1QOT2TaQg0x3NtLU1TJXTjB1wRjh7pQk
96/73agfxEDvCS/z+J27rruGrsr7ZcNblPugxeAYDnNMcFQlyB7F1vvkdBc72txM
+grqd4g2oFiEoyFiRCA0QUB2vfxANpgQ0SWODpkReEa2dHg6oKQBuYeIGP8W7q8X
7ZV8mogRRLyBbaP1ohmiAUcIu2ffqlDQIJ9su/kLQpjAIrfUPLdS9SdGoZe5yzHe
NHw8c3mb8+Xxrq1dO6Bw6PuMKBpNYIW/NsZsx/6jRnwo8qnCITv9BUZeK9alGCM7
O8HIsaLA2s/PgsZMbU4LniYDoWrBKjPWtMEgM8uAnrNXgOyI4nfNzLGZACZdnI3f
xjn7GvO/qsqYy8kVLgj1ZHWKQ1H1/f+u5CazM7NSqw0nWoS9F7pO8I70he9aC1Ea
C7sduNDHB6PBFarOaud6XtMCosjVoIamOZygCiVJIRjpk+X+ZcM81rxF317VB1VC
L15UU5zEDO9vSAp6hvFmfQKx/PLsNE1hX5PKELpqPds3iVPV+Z9sZfvH5lZbmbz7
RxTGU99YNFZ0Vgc1LY0JSgVZzN/TeP54wfJject89lhPL5j/8/Ra5Me0N/7nBU4y
o04Yowr1D/6qORZA5l8mxN2pr5js75tLWoRs483j0OzSgwxa09P3eyhnKhYjM/hI
eHxXmd4ESu7XiFiB6CnwBXiKmxGN5RL7gnq6O3ic9GIVufUOwVUm1V6tzB5eYHJB
nV6igPTYa9jY7TgcUUcgyZ10KznyGgRsy9kwD53kZgjq+U/8dP00uYRH7yTozvwX
aFbvLBN+UFaw9++qNHBeoPIlexw/QtkYEPDKE/gc13fvSL8vw8jU8UKgY5KF0qPO
kkeWefoFi9AytR5IsK348qzTpwy5pYdsIHyATfw+T64Vesc+eVckuROVfV9vIxMD
MRWKEox3qhe8bQDDoYsAlUwy7sy/mt9rmnuPjwUmUQyEiqyhATtwr4UnajcSgD9u
lxTO27peMKxlGrTJo1TtT7LSBbweVGJ7zuvEk2JuAE8vfeSBVMPOl6NVKdksq5fI
jOA73DjEPy8Cvp2auGFEZgiKbwJ6P7B1nU2Htv7C5+1wHMC68TaKj1WXPut0TLpi
geyn0NQpQ66DiDqTp9/KZdqBzt2eqlbCUr9rJcAuKreEIWs+j2iIDVAGdh1XeZWM
akXJ36yehvBm+CEFv7uRB3MMsk5hqauGVCZmocJRkbwgGwNc7yhxX1jewmVEYNsx
xO/zBOSxmeGHhmiyEf3uMx5yZtutxCCgl2IMc8BIGW2RL9Uj//axnedx25cEgF0K
1rUGVU+OOOS8JdBe8seXJpqD/vSpdbNHT+eZzgmGZgZUUFTAGsMZDxIS2g2qna5i
0Xw635r4RmjXX3ZwDnJaauxYEidCoMPPX+LnrGULNs9YrEOvRTSlhtmhFOSUEGKo
gmdx6g+38gaISfJTM/7D3akoa8Joa1Af3Zsz7Okms4ZjmD6Kkdy3fO9DEj/AJL6A
KoFjTyQw20G5aDQjD3AHzA7qN9fQ/8N+z1yYunFBXWEQSiQh/zYW7mbqdK+USIr/
q6K/IsfLwQWUajkVjPAh3/LdBffolQ0Xt1Vx/+n5Q8ykKeB5XpPxenlhg1gAwfqZ
SJZLBeRAxOdBeMpl1STCYcKazYiU5u/eMhREYFh95li/GgBgRW3wdvi7/qjy/arB
KoNXQe21aEKxbO2VUp0DGM9M8ZC9h7oV32Muar158XPJ7xQHGOFd4oNWyPLZHEnp
Z6erocM/nfymrmoIUF30fMj+2hehmF7iVDmwpHjk6/0WjykYNLwgS1Jq+Vf+4IeC
xvVVoEeq/SDkWqvjT8W76ozs1jdxbxwd9wHHLR4bFHspUTPFilCWQxR4A3tnGLUx
VdE88LqFBRhNu3ca6/vRoiOtTqvHrrxy0x0htf0z6oQ8wrE6jhkutD6rQcMobhsi
JYzzH0CYPEuZCYL/u7PiuaxeVjv3Q8z4ByRM6NT2vXO6QwuGnEl24XycW1TCskAO
UR6bLG0+qR+q1vY71FiiYGJ1DArifqdS+MkyKCSYPEvjHuJchRnORRvFGlomIAze
MZatx51xutHldn6v5dLtthbZJIrX3Lq5+5bWd3HkO5r0hbb9H7Mx+2i+W/tX32CD
pnOD9Vz6ycPbL+1goj/T/fOYd1zt5qVs/PKb63g9f0e7HIl2lJ4gdjS+d4pa6/Dh
kANAeOhyvovR+/E2xOsj8oqaLVtU0RWsp3HT5htiO1K+gDa1zOoUdtOSZJMgsVDg
O/cIP9rlgA6Wi9LbXeK/rx6rvFAJ0Tgdo3yIo/2lU3PoyfIq3Y6kiFmoKlin7YUr
K6WvOdwIkdNfab7rv/BO3kNeASEOCVo74jALEqWHzvu2inD8mKs8nRuS1hJsQD6X
K5IKgCOXot67scIPtI3pNaEmW9mlBwzLhR9XqpcsbW+sNf4JgfmoxQ1ZUj1c7bfZ
kzs2ZM0MRyxoOivq/+W6SG5nsYzNp1CMx1QOB7zn5Bv0ZrcxUy9nGaZR6n8sId8h
/SnckOA1RCipw7ErIyZMTN1FW9MSlguYdcohQRj6pd22wrsmD3A1Z6Aqy+HC9Gny
RdT90oAs0KuWzy4BGXZoQn1eBqfwgzdVakBE+Ag/dm2gcpJgJ8qLLv75f3o7sKop
KtJt5cBgQYwHbwnb9F+h4DLCvN4IWTaih4NudND4ylAZoNx/sNa6jIUrn0ZWDnbC
GD0h0zGz2n1mbsRaEtASMz2g94X9sqch+ixBuJObYgH0Z3dtU89fukUvBcid7yqA
bHrcPQYBlhc+gA3G3mJbS8vxG1PUrx6vFZOeoIIAXU/A+n0FfZ7ycL72lY+SYnn2
x/Kj1B2pivWUE8WJbV+loQ1ux1iVjF1CRmI1sm4UzKo5TR+pguhxTonCSQdfT1wB
P/eLgpt9rZ/gxCS3Hy4drtPOBtLSAXULSVBO37ezgmaXAPsEJF5qH6/UkTHFG5q3
hrI50p9RN3aYPbyiYvA0cx7j86E3lTIobDuRmA0vvgIpkYv7+jKdhPdXIC1Ep70c
VY66xp/ZZdLy7x1lHCOmkOVEm5pKwmYO0OZhKWP8s7eb46SJn5+phRzvD93Fjsfg
AaZjkibE7nECYNiE1Skp6UHYViF9fJolFYG8eqAhtQY+Z94QdiZ0CccMI7z28FOP
YBABGvbkuSGxpZxytuBBouV/1uQpmlXpGeiXGae5PgVFR7VmqaL+VgcMOR29HQyL
y8YIukNlXJHDbTpuN9RdWjigs7dPGIZinE5YMS8CqqZhwM5hgtJs4NcRwP165gq1
wYWZXL1bI9GLM4ZVR9865xZDN+EUHJsRGfD6sB/FWLKNsFWI9rBGOJm8TVrw3oBH
JyRcz6G8NeZhnKcLd3yA/yCFovc72aOEToMURKBT8l8AZQKjZpTZhB5QZhzZlOZJ
2Y1ht4uYliIEXfmdV5S6izxNn4wnm8o8OH/1MnzGDY+DPGPhwR9aoeErrVGVesIl
Kld48Bf2f9y5Uc4dVZLQ1qWf1LIS6JzhFBU7U7j5BtSx+RMZ8I+n1OZMULD0U/aC
1km2CXDlx0vIdM8po87OcYNc0w1aLtMl4/YPBODJoVW/v0YDnVvAMlJbTELuYuVB
3gvbqs++0WHon/9RAbmI7bhTAh0TkPkve44NGtbQHaRTnsub+RzQm19zbqgQSyn+
n5jW74C43uoUPaR08ZNoLwswidVbOhiFWULqt3kAXWFwiUbHnn2396JwJfaREg4h
UT7KgS8UeO8QOO9JWY6psvhVybq+k7qVJD6SvGPZlsv5Qfoc6FPrACa3l+O6MHOR
0o5j9WC87VSB8hY34ErUiezThz3b+Jt1auNnnOyoGGdLyr5FZmZSGf6xIiwp/cN4
VW4kC1NTSxaYVxsTEaMuHwwToUnBaJZyGSQNjdRcN+EW6qxYr21IZpmfPB6cQO5C
W8JuUZmdZz2TRNIiHjMdEJGBhH+YrVqDFi6s+ymDj7X7AAEvz3KT+0vEJ60EczOJ
LpiKe+xzm7RxaLB6927THne26LIFvbX0UjfVetQGU03Pw52Nr4wVrh5VgZIixVF1
D+4xvOc5d5cqxPZHDdshjES19SHcc2VZBJuIQziEjAp2so/DfHKRy7Wq5pOAbcE4
49lSnj/3CqFrpFM5A27daWzIJ6ZesamgW31O2Z/U7pywt+T0u0hRqqjYm/TunBjd
OM2Ia+xosbJvghq7pLx8hLLJ1L2ZMZF1f5cS4urnBfwFiAp0wNnndIFT3T5dBCxJ
igR+D9ggrlauUEmPhyMFIYCBJOeMs8JVNqxEBHrL7sllvKqms+i5PM8aC+BY+2bt
+lTgfYZP2OjEZWRpEvpwJ7iOYxWx5u9rux58sQfwk8H9DyPijx2AfxGhzpJFjIvP
PV5A9IIC0bNBlgNhkCwgqFDew6wrhmSL9uaZAU0y3fMWDrUr5DbubwiGIqmtdxti
/Ix6sSm5PIkzl53d6qLNPU0+z85ep0gcSbEC4XIdLUvDybNzY4sqp1InzpDDWAAE
0Wm7bL9dK01N2JeSZecE31GhUcZfNmjBPGInmuP/0V9nqXKEygfrCWSg+waV5MiF
Nbqqag1dmXCUzYOikpOXTz4bssqoJpmLEg8mMfuq8M2tdvbCT9bEejBhRP6Z3h1a
5edjK6FAqr72XNQll5dgoRCoAOJ5jwbEtoRbGG7zH14w6svgl2+Q882gwPmO0+iA
IM9MApz25tSLPETLzAXr97AD2V2DflhDmPm2oDIrDTW4gzngkfILCrEbY2/vB75A
IirQeNRN6tB0OIYMClWSM+6hCCYBmpL+mxpb7utoUXO/qxMFUy/Sl1vL+Y5P0knq
GT0MlMDupl+vQbXuKh8V8JqvkEIGU/lzoapjxPrWMI2pAv30wuanrN4R2R9Hv7Td
h2469MkqInuSn0WfwiHQk2HK8tZTER9XTKCxzPVyUYGQXGVjkWW1G7Nd+dP3VRt0
3sEC4zyW/j48pmDWZD//Xj1qKobu2rvTrAE1PrTrhHUWCIFrnhapYsKLFvdjDKqG
tWua4+vixkd7MRdYpc7zG+KQiI0qWlgeT3op9fONsVH8ZS7m4xcuVJFnRnM3QKos
lV62RYura+twuLcGsXhuf8IY+oZtQy713Ss3w0mdKYS+4Ff7u9g8p+gQQiNco4NC
1QSIi2cmx1Vr6UV8ryyTD/tjcG0zDZR6kmGqXN++U4Hv9XK20dJznc4RNXE3b4/q
1Pf/jqjDr7HTKJffFTfgxBcOvjpR+yFnDrn0six6iNr9S0ZP/sjKzUWyDiV4XZ5J
ZdjT85QHF5pyi3DXol/zWqN/zWIJRgXjSI7eZ16/yOAOqVZog3isWR4f2ddGiPBL
rmSb6oWIcWw+uVelMmY79iYW78MABTLlAxheQU8QMLe65kiD39pVwFbRDpE247VL
Z3ezDyUK07LrNiFfxdvFNMlJMwDV3fL9+9c7pYQAMskicvQ0ZXpaycASiYGxXz0G
5FXkuzMwG10W8RmRvzNqIBKyLh1IRhLoGUZDLlJikFa2LFmp5F/quUYjVy8IttjM
cMrY73UQLpePL/lN0kt001BefyvfOr1+f40jvNBdet0PSxlo4IrbSOkRP5+kCw0B
2PerhSM0xEP9pfWnqXwtrTC84G7fjJte48rBTyY6bloqohpCjXUK0aticLC1t91E
iVZ0373G3hNdg99Q5qJkWJdAov/nUWWfQ+/htEmiLW7oe5YyexKPpCvpUP8Cv/Ix
J4k84K649q1KA3/gAa/HA7uVFIGRNC00Gh6SEyRKVM7v8DB2skjcOJwBcRBkc4P2
WluZJtaC1oR7/cqReyBwvByP0L+n7aDo5xC7LvRklYCtj/4THgo5hXBsumwUoBdc
maVR7CAmoGQW5JtkKra1VvBqP57leLYwyPE1YVuYF/r25l0+01mFGYCqbsQchowM
KoQvxbJ/DaU2xzj3g0XsR5J+TKZP1u7AKuhVuFWvUpog0ww+s/aukt06xLe5EA5v
LNBwYTYUHfA8ky8MOq81xXizovfExOJEhwNh/TXTbJPRlOuqoOH0Rg/edokzeKfN
qeK+mIsiOlYnSrVLGahk8bgN/1QODpG+5MgcRXbnwvbU5uxtrNC00ntjFhPyEtcE
FFdUefsCBpArrLkBOBOJkm4Ya/xKZsG2xRNsBWoZFdAOAYhCYxZiU7WUcwZnN82v
yLG1q0fWs4fHG8JWygLKJq3F3RwQD9qo7Ec7Kc+oi92SuZf8f/2hTDqWsCPYKsfk
JfaZ2ObDEY9Om/NtMWMc4FTV7ymwsnuhDn/S8IKB18FHEivGACchbdwaiQbHegLD
pWi16x5V0NgflfxJMt3HjoKEUtkWJZQbi9wErmDPAfg11k8rA4hF/g50BTs9Eh2j
6cAr/qCQNyBALC5NuxRafDyHZtYWsWsDUqJ7ed+HpSxizoPVfAvBB/nT7DLlTAVZ
CzIqaA47/yXoVPs3LvMRu/vWK5Gp+ApMTnW1cNzbrR45fkc31JLj2HUwVFuJIdMf
UYrOHZHxo7Nf1yGjzllQ6NqZ/+6kOu0pBZBu8iddAK4PK43ep+bsu5/T1yl+qsvS
ZhMQhiSWHWCq7VnUQ0zRl7mWto0+dYacKeLYoNiI8WBH/au/EKxI7vdlCfDGSm+C
wEuM2X/vPQZDdevgSvlk+DLpex9V6OZ3hOhXIUmGBnrXQlNE1VkoS1yUwzJ02ksO
Sw6erfb7B00Sk3C774zFQSVFqRsFKVanCgGgj1ZeB4nAdF6bcIiT+Whi7t/KwgCI
Oyr+uTV5ke7Opn1T/cG8KRCjr/oqJZmtnPTjHUYs8rVQLB8eZNRnvKJ2G1JnLqnz
6KmCKqQGdlgQzYRNrGSWMJjdaRZXz6udAy6s2WGQCcMKBv9Wuv2IQJtt76YysC2S
wPF+VxFTEMCLY7h4p2yoIxsnXRG+niqcXV5bmEx41U09Jg90ycRkF/1v/XzOHLMa
4X7GWtiVY2sdTNIKelhQzv6EACSlsC7IDETAOF+JYNiWi/4iq3UoRnWFiUzlhLYF
5eM+1td+l7zegO8pa7IwNW+D/m+lCEHXvh/2EzrapFIzEFrJFz2d2NB7MkSbGsBB
QzD3mDPOhrADr4NcA7T4BREHzYjY9k4ha6Mi7YdF9JVyLCOAGUm1uypeH+riKGtL
XImWHy28e00JU7cXG2R0ikh0rBKBhTWY1nVPWApTTPLHwaW0OzY0RRNrWxHKr1Zj
LMyA965GQua0cNPql//5r/supElFWESDM5RFkV5XwpuMe/QIl9PAsa3Q1t9Pb4lF
nfpjwv8O145ep6LyDny4NI9h0HEuYyD7SLbAVf669f2AiqFzMf6PpjrGDT2bj7gi
oyoGBgaDUTIf5YPx9/EAiE0ryn648sUjkc8P+sb7Dd2tcgQuLBSFTnbXavQ554UN
fGLZWM2Wv1Isi+N9wTr3tXyCmalQ8lLQ8HktpgT0kQgBqCxgfy2vQLeEcW65JXyZ
lcUetiNG+Wu81LJU2gfDHxkVOKgaMaXYU4YlnsZax1xqa1eBoO6cgYDh45Pik0zl
d3r+n2HUQ7jY9dVM6MyU9nikkQ4TqnYNrJG2IEMBMTSpctEgOpRf06Gfsj5QEQA4
EJUqwILWGRgz0T8ABqLgqENmI4CzwbXfKtfFJfAjY11Im/+QzKl8OEFRYZQr0ieq
MilHiRqkikOA8uvkmEa96k4/n6TVrgMGhe4Pg675qTizCOKQj986IrUIRbFl/hiy
AV4gJTWTj2h0QSqPPYDoHeeQURJ+m2dKdURfuZTN1g8UXw1zEHxo9smLMtyVcd45
mRspjOtE8jUvAQjZYkl3SCy1xAjttDoNDvIha4JdygujVWvMfbHhwCEGB6aqtJCd
fGRxpXbCI3L/c8/ammWG80TE2qUzs9VMBi8j5zUGCEUsY+YRSvrbv1sPyq1036Ej
5qCCZauf77jDeV+y1tK7A8r3iWXgn//SHxi0JJpY5H//bA93vvks2rcVQfQeettF
4XSzenjjKTGw3He3IOOfdAywA9xtv1svVn6wHsD2Rkj3RZyNxGJk5Bp/7v8WXfBh
qplLMndkUBiOUXwKPPgro9A7I0mnkYi6yyXmXzQVDJ3ytAOYcZ4OI0XEQ7ff3Mba
XbCCRsxmDC4a/mjmhAowqiH3aENy9rPUsqVIF7T55Od5LZwbDcx6+j+zIAd8J7Pv
Pzzk5D7at26ulN770XHXuNuuVw3XhQj0+3B6LKFHxZ5fvI+wT9CCdL0p0eOtwn1I
QULifMfSCpupdwGZEnAIBiPvjpU3rkMa46SoGhK3C95Thp9Awc1bg8M9Vvc9vBD/
dW9q/TOgycb+DSW/oiaoavGXgld8y4sKJftSoiVcRKY7SMLqz4LqRcOdMGO4eRoP
aE+j+rxICXYvZ0+cJS3/rq7I56PL6rISdjLCl4lL6FPX08D3SdCc4lE8dkewlFTF
1uBMOG+7x+TQnft6bIKw0XzOMCPi77Mmqio/hqh3GLSUBxghHdSHK3MlmPrzpKnN
t9zBtoAlln6yXMWIdZDvnKX111O7uzzjmKxkkEkM6UP2KDQ+12lmY6TUtSdTxZr1
vy1J4MwHBhIovfuTxC8S59hRqaXMtgFI9NFZ1HnI7BeYM9vlxhb3gJHd6i8sA00K
NCvxDn6k6z++WSBdp7NSxkwpzPSf9jaGl4DAwPg4sFwma5ouPc441JyWWnUQoov8
5kXt8koMQHF5Qjh5++Di1UjpwDwf8v8DtkySGTT75/OA5KOAYC6x3HT3pa8B5gh/
/aclxCecHYVfvgtj4Rf/h1FgMXrCWI4i0+8+wP9Jqlbx04K7LhRvzEpFPEkf8Itm
iLnUilh1nnKVTmzfPpNUBLGpVj/tvVBXrl6yiJ4DbqfTCQaM/N6c4k+kVvG8EVzJ
aB9zr1coitOkhVrMUGhGg/ulm4ut9KDJZCS0s0llbe3wq/Rv8+YMJnrSzGSZEa5c
t8cPz9aIT+2FsaeM4GJjUsQZXekKTqIVtmjHyq2hylZXB709o+LkGhvEEggIBW0l
JFbGJYEa3vWE1nY3F7nM7/ELRBPZNARJ8PnJlI0E7UlPue2BezU+gbI/0ICbEVZ/
JyPpCFbTnPthfyLIZzGVOGn2UNfU8Q4MQ8KYVwPwtFBlMg1amRQIqcsCN3oZDIkq
jLP0Fnn4UP5lZAKJmXh8MObhWdx+3ndUDT5jU+MxR0iWsj/WL0USLiTjZPEElZev
Iu8OzgSlkwI0zlGMn73nbbFo7hwqnn3QFfARUD1piOpJWQTkSPdxJqw5FgMMpuVj
Ov1+OsNGQMTgoBqGLi45WeHxKJniwXqgIGE4YhsxJ8wyaoX36ICsP0cVfqMCxhRF
qeZvXWcPZfQxRGtm+jDYd+zqrRU2vjuHTRPhPlMrRGYq3ZjNQukRI8OukM1UJiuS
vuf8EMpVfR76Atv3qagvz0BDLxFbdFLrE/okmk+DS/0A+5bT+yEQE+VVxLu36QBy
UQBP6re1abWIm0jG0YQvhbacNcrxKHY9kHTsuE0zP5GrCZw76HaDrcc+qAjYWm+u
tL5F5zTKu2hHr6I+JSUDKOVvESnPZHlrywa0iDVAaNDgwr0KGOIL9dOM87X/dtQT
Tbwtw97JInQmdrPjIhC0L3p0Hxo6uObZofFG6Cmgks0JkTYTe3xmGJkxzg/q20ls
7WTmfU6TF1OmgNEFw2QzvpSawndeflkmOnJmpIt28CcvJChFsHXgGBV92hxwr2wJ
QwvmH3m26rGdjQAXxwrrsUL21jIUCi2PugwaT6fAH43m1BFWR/3wdPYcIxudyvU5
A7CkbFdpjLOcD2uLT3/qg8co/kjxf5XdvjqqUwG7pgRqQT8BIYTc1apmQu7UGe8F
j6LMi5c6srzecLQ/tA375bJYnJoVT6jDHgYK6DuoIomqHwW6oSKicC/TcnBcWxZC
L6Wcaq9rZPHaM9Rv/7bxdL35yBizbMiaN22824T3SF1FHmv0+Z3evt3/eVh1B28O
znCHNiS+p91qbjr8moglm9yhigjowyns+JUY2aeqli4CxCfyMpWekV9pP7Miafi3
uCZ4XeEZRtzS4px7xdfmKs7ZaVd6Yc1oFW2zc3WhMkHxBX+TNbnBwXO2pMwEUUzb
jUZ4M7dDV0/+w+jPC3tmA8GukzB1JBM3WmG2Px7RvflCpIVJlZ7igDV9eFrqBzYd
G/FeiFRcrCZD9BoPP6eCOa3DI7VQywgynPBzX4sYIfrOVGIZsUdULA/a22ptQP/F
fc6jEDaZGd3kfMQRZE7vmDwyxtwD/NvEqhVZJsr3seNN4YX0MazqIQ24dEkOCI7Y
kLousfG2wEwP54fJYYhR7uoJcN7YIHw4MKUyGb5rkFvrqpaMpn6xALbAZCmYRIDl
xKTdZ3lqhTFUEY5gXSvdougza4bXNNf/HWkH8ldcZw0UN3t+XWWvxHcqrWfRXbwV
HqLlQBVGcki+rGUl6eMzm57u1DWrZ5Fygdt1QmHeV95KEsQBjO+9umWGOxmvuXGH
+qk5RVosihhQ5NNTrfEfyTgnMKJr1zqzoTbUpcXNLvkHJNSygcSKRRuxhySwLm6s
B+4Aa2+wEF0PdI0mo+la3q3K0H0NGU6tkw6dXoRL5m983az19+MwCCLu2tJNlNSf
q65+iDfhvb69BFzLS7/tCt0RLPgoHxRtMGUTEDwVB3FNw3Z23CDCm9smzi8P0DBD
Y/UYbay6+mkPLFFZMbMoK58V9vG+ZMMpiDx9PuxZ/h2Lmz1j3OjypTdpJui9w3z1
lKt9IwwvjH9aSExlSpWbdC/HorCpxoKQ7fs4E0mQJKuxV+3rPpIGnTrBJyR11uCT
gLdnrvPpl/xX8YuvDoJ28q5putoZeEXQMdP8s9oDsPUpmjNegQWU7i17Fl2fEBqP
nxkb2Z/zCexMT/QBNrQxTAjzPk2gJglfHCRwHuCDPUBk2DLZfKb1Uwb1/Bck4BoL
DXhpap+cCiZOp1Y7lDlNSKNPcEAOC6ppgGRrqRCpYSgB6on6iV/1rQnGfU0bvHCR
4vsXhYd31Igu/r5rmXivD0QDFvPr2tCmvEiRHXhUBlkw0qaILilSMZ6p4jswtdqp
ukLxd+yXXqL/62S6rbEX49k/zNy/NDHJcp0yIO3Y/jAik/g3JCROEIkfUZN3L6LF
A8mReVKLX3KS1Qxc3r8xH/PlcRQKmzU1uG28o4mKTbuPq1Zzek+sm2EQfQEbWkql
44mIXHyxhPQ43UtUESdEtDRECCEkFn1Vas1isrt7f0983JYCmGnebz+iE+n/un13
e5ZtyECYRQA+Q+EgyyDebe8PlVwFH5cSbMycCkXSk/NSnPr/K7ITW5HagOXwKMaw
fiAXyK0RdYH9Sed17MZsrN8gjjfQOHjmUAJvC1A95AsBgLoY2fpenasdaB5k0uyL
78adjd9RcztGGIXfJFPcU+gic645FlanXyK3uPewtQsnyHqo+a0kxCtP6K0wM9Jt
r2eMLY90siFIm31N8U53BS6cnM6ato/KfXOj+7DGb4/zKD3hlYV7eOwTi1xau8yF
jwx088NU8LUKmgCS61HjBey43JAG5uwvK28uMso5WXZlFHNUdW8yEufh2x6+b3Gh
W4/35TXk6HebK4EyrWLzdPk06dbpzT/YQ5HOXTW6zEvYe+/97e4v9xZUYOrvn2Q4
mcfBzkcT+VMfs+np9DcBNf/7hsZ+Se5e16/FAsUvfY4E2rmCRhwZc73O4e1RiFMm
aKQ7Gc/H8+bpLCJekL4cxb2mT1foCM5U+Qk6AQuEf0nkfnh0UG8lIiN4Dwwmw2e9
0lAF0uAVOe0Ib/979Qypx51DvcvSvY8I/fplg2MFW35SrcdrvVkKbeUdHMIOqqwV
j6Y15WDz4//A6TrUIxlaNjxQ+bpKCyHO56jHz7oVe02xFR2fU4teptKxXbvcDGsL
oK9sxn/j4fsLocVRL5Y3Y9HNX7YTK1jzGlm2SfuQDeKBZtU8o1aJ+drdtqMhKwI6
R5haehT2I/4pHewXKEHwcu/+6lY5UXLzEQeaG9j/GmrNi30htL3GCrZa3HjuvquZ
WaqfDojgNKfIssHfK4sguk17Io12O1pHZNNy60QU271iky5YP7o4EpT1etPRQAMD
2dqeBo0TTClpv6YGGnbGZP6CBGB43tc67lh4Rs2BqSUhhxp8uCsOZ4SYJwqjnPMw
2GjE9iBmXdwqPaGuUScDtNFfnpvv4uRDpe2fSb8Owts7IUSrMpR554WZPrFbuFgk
kWfuY2wfprGJRFZUNwizL9B4NuMz39MNexdG76+j1wqZEael62o9iOASlbfb8SMN
YO1bWEXT3+b/JEczzQ7zsg0mAXW0qMo9SwyPebioccKxJ0LSY9ui631fZL0mshhB
p+/YWiCNvu9s6qqD0FwFrdgIgqoyJxW37ZuHY4p9G1BvUW3E4G/rHDBuzYFGOGzs
/7GUElEcaT6rUqiVqG4vLSEftEmbJcyPPQ2sFoqLsH+Q8DDa1ys3cPfXmbb+f9Yg
/LD5bzZ/U3G9KN38rCW5dan1S9ez0gP5BEVZWxLHZOEuGrOlcf49VtSH1OGjb9xs
cdFPpvQ832J4FNmyCrsZynrYN+fGSjha1jZRxmomEEGfAHtG8oLTsvIgjyQW7iDk
4Jac3OtC6zHR7g+ssAZjlE/FG56l91mRxSoep0Nt/FjZ4lDYFajlPg7Bd4iqGidm
3r9nBPsh0/8LZefpWzFUFB5YktUV1mARqzw/Lgr1YdGQ98zmeFeTlsPc3gSp0fr7
hCilfQ3LC9TfrTcxYLdaMuoYQMXz4rtmjrqVgRw8QEh+/UG13+8s5O9KGnj8wRZn
HLrJ8TlX8Facq6nLlKn/kx6UstIv+62tAVG0CDgjEvkby85q/hVQW5PDpltLsE+m
x6QMydYmddcI2DQ8fNoE/+Z6CYF9GP09dFKbA59qLjiAEsex9ji/rHvOQtHSuUcY
BMwaTfJeczlCypkPHocWareitY81zOTRYSjIdj0RoxTs2UgFkuLHoWOztP5RIJPN
4IlbgzD0cQOMNE51UbWa6M14ylcwZBebQxUV9D2bqLxZG5dyWoNYX+ZTAShUEh94
G0Aipd13sWG1eqj9B1kMTyPfK9CeFq65yDer+OmHwZaBxO5ZLdQ6Wx9QSdyGb1FZ
mdHzi3Wk/P/EuYxC1qEwklUOqC2BJ5ROCNKl2WV27m5ZWGbb+Ogb6TsF07yP+Ys3
CIZNW2mnS9R2VoVcYMKok6hP6dpXIVAmcbqP8uXS4abRRmpRUTi5o8bBnkSCewR8
O83sA7v3RUktQ3KycyLNDfn4qwxiwGeVRxXK6Nvqr6KWxNnt1Q3VxoiabeHR2PWr
cY1NGmSJuHW9z8Fo1xQeijXo5BBApOGmnN9Jo2RCkn6Jc+n1ZifWXkcbo+R2HFCr
RaAeWkx+cT7f6kB0JHfehvzLjmyAIvg8HubSuUuXtVS6ZqodxatR3b0ugWoSEcB5
E9IqBKrRCbGVLydtWoN45HUcWrzCqG9Zaj6yynC6WPC6ZZMBcyu+DahqoyVqorM/
zJjAnaUuW1ShxFhC42dnl7dskJXk2qehBSJfMSP8mhgf80isP+em268HO+T75Ti5
whgEvAEYIFUsvlyOZmGQPeQA5GsUoqJWguuZUg6JpOXaNI2JC94pADhTWe2C+CUq
VJzVXF45uIsqFeKy0JVY1o3I6+INL7MC0M6WXuDLcHGIvoc5lFIJdQFIbq1Hmsjy
plf7Ya9koOjxzblNk89MQD3wc7D3pEnyw5MliqrrqAzufSe+FAiHNfMLhIkQlOu8
omOda6ASqAitLZyxNkv7oMnKu0sfhkt9F5g9QZjYXVafMZSdgGFQFqyV76paNhSX
NpEv96UFddRg5Nup8f6mE8geC+WvMP7mFJ2N2vfNRlBjLelnam/aiyqnd10Mugut
qHrVQfFCjbzLc9MTy09gEUlcXg/i3jIPNrh85xzdRgkj8sMPY9+QZI58cEPs2rzd
HPww2OlBlUJtOrr9bTY0Ncau2WaMO7ZPiwSF8EL3a/SO4zk04Qnjix5HJ+/rvAzA
VjNgILcqHlhbFkTLOCHn7Q4SU7885GWj1R+cmasNKIg4vG/uVZkO60SowXshR/A1
XnpvawDSvmZ+nyATxfuvi9RIO2jY9mOI3Ao4y9gKWXkYlqcv1ho+rmXr9xgCsTTN
KemByjYBQKg/TmOuEXLjD45ou1/wfCu0/B0gK791W3pN495lPTA2YBdLuv0skVBv
PeckvpxPrdj7LrU3NC6I4P6IVzHlSdmvPhoXzhHVu7vWGSbzPIb0s53ZvKeIOciN
WGBt25LALKOm7vqQscWpFrQ1JtKPveVY7BgU6BLN6XBdcAYdYKU+CxIK4tCqcaGf
98raG9hsHJY1RaHDYESzNZsA8wyUsMU/L2+juBJuNjCTV85zLGYqm7ijaPj6L3h4
0uSAJXFrrvp9zYI9EqiWaBYOSXmME73fYxUySmSClua96sSn2gmqUFrOmTO3pF/+
/VqikdNd9olV82YCh6pbRBWhOiwSDNfyskhDDc0yyHBwbcWHsQwb/nFkK4T0a4An
0e7v7lPnIV4gNeNTAvSv3yJscHiZkl8G0KZyegjlbyKyjICiwmuDGp4z4O8Svqw2
Gx5hHbnVn6WZaS2d4q/+l3SQmjguRd9HvcqifAijgs7xg6hYzsA2EAk11rsFV//L
6yaEhHeAdCSOIopzGXxOrq15tBjg7Sj/UEzV7eqrM6hXvO3pyzFCF1fYzQeEsfIR
HevpYUokkK0zq4G6ZSUQSOMgFwI6TRaps3aLgXSKN4PQ3xADhPz4KKP42yRWPZOI
FpLiZDykdpy/g5AbOOb2uybDoDL+90WnVvW646jMnX7k/zZu0ze3ctuZBpY1PZyT
pSyxendprYpNA65v2Mw8H9h/YHxtfE0mA8Den7zO0ug8BqDeJkVO6ZKI2mRMdRdx
AbJdPU8YY0nZGrGGXH188A==
`pragma protect end_protected
