// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0d0tyd30mvzX2tuBFTS8VWQ03fwK106zeMgggtV8OTqhNO+FbNFt9mTHpu9AwdNp3OvE9aT0DwGf
qRNjeb66c/+uEcicSBL20vc6tltvYs2ArjEpQ1cRqFhy8cWs+ixJ7LSaeLH93O6gi7TXTr2LVwLl
HRRr1FsVZ4T5kxkcIP6xP7wQ9UHYU0eZLXfsEfgVjexk+x1Y4x3XG6Pa9yNl87Vq/FpjHVv1duAt
xSRWYACQTLSU4ov0r9wM0Hn1sR6253i2wOvOm66sn7W053ePzgw97r+1PXLu6V5oGrj4R7kiEoYV
VyeImLBR/9e57XgZHUf4sgH/VCuX5oil29jcuA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13744)
uGIeNVwYcysGs7+MKXSQX/PUQ2FAoCSj/Uwd64Y7lRZRloWMf7OGDkOmN8J0Jew7rnFFOB++WFXW
ChIS4aIo+9TlVS3h2EmqNq2KVArKrqu9VFOoiH/1Fig23r03y/r0c8xeBd6mp5k6cke0UNkIV65D
r7WvwMeoOI61NACd11wadyODcJbq0NJwiaFJZiGAIcrUcQKYITRd8/idfAPjNzf0Wz/MYeKRQmKT
TWbC5KDX6XOhBKYKjssLEseCFwAPzWr+005waYD6Ln4C7yuS6vIBtJxNFRVlMowyHR+P05P6fT5H
gVMcmqM8ViUwOd3eRCPBVyvfAzFJZ8TsVi15Io4V6y5zu5lKllOYUWkQRp712yy0yX9WelGwljGM
X2xiZxAAx/U6Xbh7kE/WC2JqsEUXhMBew5jptPH0nn5pXHJAt7ssQ9RDandAetkXPRRr1LaVAiu0
cnYDBvOP49p8i4IAF1Mtyt3ondpKl3R8bcasHCPnAbeYMWZWWQLpf+YNLINKEjlX6xQoqr3MjMWK
6wdec3zYdoDO86Tca8t/lz6lZAAaSjFnUr/dx88xKg/QBtd4tK9t8HN9xOS6AYBYm6uYJZXkw4HJ
u5CBEQyuOr+izNbST/wnvLj4H5L3ZgxJvMQFla+z/+WiHRUjq725gxx7HdlNMzvsBF7eMFtpT2eg
xbgVnlDzbXq4IbkBxGuwQBvuxfonvr+FX29KhfZFzb9bvKW9KrQsIZdkFRYfxxmnHzQkI6xQ/r3A
qL2Z+x76W9GWBmPxDwJZm+b0gkjHvWBnRlFjtUQqJf2IMR4mG0R27fgkana49B3uky0oLe2eXCUD
dDQjdmz+XsN82p9zTlMDxWu+N87XMD8rGWm6t0AclxYM8fbAssQ22yxy5CnIJ/MvJ6SJo5d1Kd/J
51rOiGtv0EVFOw1D9rehZntcbuac7TCPqdIruxlDLwjZF6t2P+V7PbTcFkfeB+pmeFyCQdqfrEF7
VWC4Sl2m1P6Q0zYpDoB/2aZq1dXWccddOdet/pe797gL0rtDeEFKOLSejNJ5PYkhvGOlvsp5a2Lq
7xr9CB14KT0e50VdNIcPfVazoNNa/aDyii54p0xCJ3R3JAr5sdQI8JLqBVH0pS/bqR7YYAYyVszH
4yeZ7YMDrQmBS2DIXR6GpTxLN1XXJkNm2yKstJC0LGO/NtrauremK7y/xF86Vivg3z2cMvQvfldc
6cmJvT7SD5RLfZq29SD9Zn6qktY3XZu/E4P5HBjkZgoIhe2YZeSrJSukc9zHSzWp9t1kora4pPFz
49onBwJZdQX1he4W7Qcrvc/OooWLgyE0iRRw49M7G8pw3/8baIIO5/BvLkRdj8PJ0pkwYh34iI49
/gjMoX/t/j4OQgTtsmc71NTbckcOU3fFUa58g9JZOYR9HqnojxHtf18ESkYczbHIwhFWp7lf6Kid
lddeb12KxQkDjHPor0+ExBZSReZOVHa3wcYklR1loDbKPyR4wTvdqhFkoRojQfb5BMSG35vQgfOO
qiW4rULqLtKtO2VWjLZ5mnhTjScYi7FS/4/iETnw4OGamSmuILmXY4Emxs+JqtsacWvbw6PBHvaj
e3r3nOLxZy94eJ/59DzA2yXttiH95xBtbMfUBEB5evR69H9OaE5SNBLHnzfumx+SZLh+CwStnQMs
jqr/nSSC4Vqp8aOgzfJZH8BiPeDof80hsD2YNVDCVQlpKYRMIHSCabjgGOFZsf+vlWcrbtaY8oya
oofkE7hCP46Lc6hAoAJKv59nQPe5MI+hJhDi2L2TRqQtBvrY7YooPVu1DMYKFdbMikvmDG8OxKWF
kYCbxnsbSg5Jzrbu/4DCgpPC2dWuPROJxfMTk3g16J8dFK7jVnXTWb+981vzHJ6J2AR/GHpcJ6/+
kB0gm2Dgb2usBWkZvTTDnKEszdgyGcOOkJ26Sj17P7PZyGDP7EuY48sSdXwT0dZK2a3z/RyECQYg
tC9PgRQR4Ak2N+60ye71YY5+lzp2TF4MxgUlrCYWx6JNK6WMNHmfQqbAZWmi0PjDKWmnkfl/lu7m
IeqySEsgQHjHZYYu9gpukryjkWnj3gGUYzaAdsBoeZw0EUAcsq0Q0TffC9b2yzcd2LoaCLnVuFqC
l0bmsO+gzPtrVGWvoyBHUSjiJuf/qqNFSXWhwIC266kEtesY6cLNf0YM15VyerhXodKsSWYk+eBU
T3nt6Z4X8gLj06vW3rufN0wQluHWCPKtdmkr2xSXuVt8+ovj3dyv0Q2T9ijcXj+OyWOT079MPx4y
UvFtdUThFgZuQJ1Z+RMZIaVhayxVHcJx2Z0pnX4WSZ47pLgurYQGUtu/oOj3505YWiQ5AfvVLIpV
j553mHuaTTLsh4mcnsgxNdmXAmgfU07Tg9vRW2UTXez4mUE8VWetN9WIhP1P4uOHk9KWwjoDNdDC
qQQWDSnj3LQKQ6vysikyRlzJOQ9vJG0tLrfEPeT5tyuohzYRq7Ny02DlM4d08wjmOUF6S6MK4Aqa
Hh3BECNOLsB8PATX+Dd/akPnSudiPPoGXFl0Ek2G6JAM5e/8GshbM9ML5tbBcIVtICdFAcdj2NVJ
NaCPSOQRrLOQEV1f41oggjpBwnE7W2YCtqRNxh0DHD2etGqhEYrYl8GBeIOSckyG5oRSmCCJOwB8
CySLziZLPMSZpuF811v3KnwBnuezC5hu7wTCWPiWAM1w6DRhG1oPree20Q/7yKnGbfE8gQzOw7c/
DxiNtxtpKbEEPaycQ1JSe9HHrJHHySYP7xIzJZSrlPp4GsXRLtlD/BjLKixC2DUf7l7VeYyX1ejY
OZql/wJLoD93kmkv0FgrVh6FseI/Q5q/WocxVMLLPkcbp9QmrvaSe8rxpC5LkgSXhztZP6Lujedf
33E38IEC7s56IOctBZ9djBs36UM3tDUaS9NrXsgTPw6EZLgTeDjc2cacPiMVOaM7q+ka3kz+V6gO
LezkeZ18biL43NiWl0lHHfaLylkEjoDjUOszYHjO4zzGZlnl9QnX1D/TQvuKHfl5JTtogxUyg1f/
nwi8aFbCPfXmJwLGzZryZKXS4HgOtEV7PVUcpIyAKexmkFHtjDj+0TDbpjfYYx/S0daYDiZI5pOx
9ViEchrvkSzvNVb4HbavH6l6v+mbvpAUbbl3QZazT6s0d8EOIDes3hdTuECaRJHRdyizeYkaVM1M
KkTrmQJkhVSzS7jYz8GI6+7adTkyU0lGd1dbVBoQRRpUpUJI4PQuNa5coFzEDLRaFhuDxXWkbjyi
7BB49hDF5rX6Y1LjwetCPCgd4T6v09gxyYLiLIz4rfYzBw69vf5+sjlR+DiT5CU87hMRITxTPDv9
mU6wK2Fsf08kaZ+6aQNr+QE2f4WEs8U/NsxObEV/dPVYg5v5r+FCSOdtO8SKfwTcfpKtxG0bPvbK
/2VvUx4Cw5C0D19bfigsHYY86RCU2YJLWwtcwDDUwt4CPI1lYHPmdsSUtRqrtgUOTQ5DhOWtpDYQ
1w/zP0bCarXxftvyb4Cr96B4qfSJS4w8t5XYzOiN4fra1ZazNKkEtyutzMnXiTWxNXcwQlTXBsY9
WbwjYEO2IR4li8P9NICyHME4DM/OxPSdiNQoCluPu7L9cfRl+52yH0x/LEKA14ouIW+/bSD+tlM2
ZR1bi/SF45GNMZ2grNVwflSRVV4X4ON7NI++4KJVMT1PPDQ/Y+GG68Enrbw/uJ8CmCm10xrH6cIm
K+clI62gtdy+n6/HwSZA+pJbMMFDzC6wlVzGD0eqNR9qp2h7UZc+bXqIVfdrwDwnNL7oC7U3keUD
4feCmqYW/js8kCcL/D6AqMckJiBjLi23DjWzSiIbIrwdBfEOgHtvwdatlcmvVHhVEKU+4IXpdUBI
S+MHScuV4CFWkoIWaQtGWc84mI56EhnBpFbCJO0A7djCp65G5dgD8pzFBDdJsIvDsn4INp412mad
6+90lUlEYO9ub2jISsSyqiHdF8oAmG+QDXbP0QS73SHI5jBo0JFqIjvhn+mkI4bcBVlN7z/f9XFA
19aoFib6DRqsanxt9YEPZPjMv6B5V6IOWrTR+NYHHf3liNwcpTCHJqnbxqlPhGpEao7tf23bqeFa
Gkab6gX1Ihj9o3xeIAEy8zd0v4RTOyi0SAwpZV0JmagkLFAN4h/duzcQViEmzyFvAhrfk1e6dOs8
uo4lir/8UgTcdVsuJezImbTNeXXYEadSXnk6BMwC/yDTjJd9X2358xfMcf+CNfVKsEUKIJ7YGrPq
w2aBlNfPCCWGnRuwnz2x0RH1kPPxy8nNbzUeMIz5FHtSkxBQeL0Zt+WMzA+oIBEAyEhMmh6hMlDJ
xclcsIRVjJ4DDccAPvYnw9GheOhSh1fqWIBphcxr0CiehbxnDQDyTa8RN5cBbbbLPis5K8zWgr2S
mEvgzvLiAUZwL7VdGc+D0svy2oBtjtsbJPwrtKyDksu1BYg9jiEIYrCEZhK1tfmHRKszXk73Cdyh
UnwAT6QuPn9/9QFmlLZqBFWA/W91oDkpXF846bzd2/tXDYVmHxigh8mBaklD6A6lsd2lPUdNdwoz
wxzlBVnZNZznPF82TEKqBLJdWZ9tfYyZB7kiYjZZAZjH0kyGwHdNesszwnhDO1KXA+412/M4g8Yn
/VRjradD9OZTpYKdvscmCSSFyDqbNeLwQiBp+TJppbJpsnTNYIuLV4RAcuwq1jamvRBfrl7gZFb3
Sb+EAPVsxE9CfWoapumiAMTTAa5IWBz7yXMAMuJtTggVGYE6ZRVErKCmbW9zPfspCw/2w9UfbCCd
+peA8rrf6cyJoGU/iPiy39ejxdvNxV65XYhgfmK+wTVAwEiHdGRTURQA6gF3LI6u20ODQlUYilih
ZtOGWuqEQ40pWgsSRIRaHg6dWgpkJzszZp3DivCagyOkMqxAoxn+McXJ25kqfCaOWD63PtGGm1x5
HMcjEFiA/2vH6UphJEuH8LW9UlR/Ck++GRrBGhs3pf6E4a942qumsJRiTIgPlwyh2L+K24RXjEJD
J4KqS9vDjo8oUOiHPTHhR/LJhxWtMQ2wNXgqaekHkfGnX8Sw2nYyHGD4Usw/54wRwL+WaGFQRnAs
oKpzUCOFTlg1Ju/6ymXPYNQY7/4gExBDFH6DRcbunNGXRfWtNw32QSk2Djbh1vf+VN3NFtTBDXJl
UnafPw3+F2pQQIvzYHvRmZqV7EM+w33pTraMWnr6urh14Ud9Z9YaOopR83LNN+o9QqgfB2is4Hyd
LK5zNwk34pRP4BnR8qRqSEEFCSS2OXyZd8H0lvziHVwyqzDQ/kTJdUoGTTonQ1OIsWcKZoFMYlE0
71H/27clhXubYMXYPKJJMQ4O+8I27JGoF8In7FfcFEpNkz5z89yq3jOpKV7CBr9x6ynafSesluuB
LdKGfmZG0cRsAVcNkbZN4cXuJX5P3PQ5J8z+ucvUsUw+tv6GZiMpKV/EOptmc586ww/99M3c0HdV
z6xTtE9ddtD4Sxjg4JmbWLp1iUwcDhmwyIXSu5Lx24sOo0Wyt1BiDUXSwQE0vNWJaZ4fNR7mFnD9
08f0WJFzeYQDikWGtYapS7aZoGG4K6WnZxuwgwkYTR96d3BB2LUWaIz5MQDV6AL8yLN26K7gad5C
iak9PSEWhCc9e6jC2znBXkgImoJAVBrbVz4pH+SAf9HFLhRSzTwPYroPnQGkh+fnJ1o2VzxB2DNs
h30gTTVM+OTib8ZFbZXMqQGDDo4KBeqqHMs/YM2+GcgLsxUEaKOQ9YRPoQdoCUz0QX7hndOrMu83
jthUDbai7dw9O3SYaqXrRgwYaa/vLI/BEuAsL6/XRxuGOp4ThDkW4+NYlkZswYLZIuDNMDM08g2s
I+QIiSA7f7fIOa6UqKTVyUt2dgtyc0NrT/tAeYKGHkPTaPzy6iZCIdoHGR7Ags8Gji0tQP2AMZGR
tqGdlQ04C/KYlXlH2NkEII/6BXnWNG6MA8yHLzXiaVcTUzB2a9KP9Ksp1FOwSLN5l6tYfChgGbeE
3c1INx2hQusVJCOkphTsUAvt21nH2RH83Eb7XcsFDSjXLZFtGXjsGWJaxmmLZrzmiFq4QNIa8Am8
fMmp49kBZ6Kxg5P79I2oa0yGKBRsLb+YsuBbZOTkIjegITYTbRToGZ/gMlFWNuW2WM98SJnIW4wb
Y1NucnP8mA7rRyKRipbwnYjfTGT1rm6ivgyR6VzuywPvtTop4V6/KzMKyBZuCuP4e/+nBCj4AOcG
SHUju+snILhA2kmCfTFx6S9U7e96EuoB5Mg8q8NxV/5lTce8TQSB06urZsEXI8R+7cBXmfaJQ8r+
cASUOFQwmLc5xdV8LzHakZI7P9w7tDQm9eh3L9ur0EPbOsmSw34huVZBFEsIvKRwRaekLYYS91VQ
/duxGQZFgMTPHPXfuxew0Bbcqwt30Y0pLRhwh4Nct9cOuvwI0EMdk3GJRhdumpMoJ2jR7WLE7kB1
Mf2EPeKUiR9Gy8JY3rmXAiekolT5G3Pc63sj+7YvM0YGf6nsDXOKmyUvGBsxgiqLN6LHBz2MySCY
rnTyKYWfxqUmUJFYszOR/3/3GWAIYokD+2APudADqcjy2N/he5A66Fa2PSXQftD9K/7RJ4R9h3pn
HlxF0fNl122NxEAkKtPsvl5Vf7gjW3caQFmzHVRqR/uxkXDtr3y+fWuwR64C1aJOmy5qjjt8TU80
sx5UII4+QOTLsK/pUU2lvmFkA/aYdEbGn06BPcmwbRZCLinJsbz0WbTO/c051ys07hRPx831I5Dd
FM5hZivAEqcwXAol7i0IvgshhIUfEtKLXFtA9PrWdp6lXgBZF8taguGHEJEAmg2tPWHhZIWNUysL
LjJfuUHlaQT9ui6S4sDbhogV85WU4WamUmzXvWGak6gV/lBS3s2SJGfufme4QQYrwlj8ar5SPIJ2
cnwEI+8f/RwnuNcoxuuVaSBCIQtMqPT850ImsoojEWWxfnvIX1+Yl1C95Nn7Mo/aWq3RoX2mSCcO
mtWyxibjmengxh98rxA4Nf/CspCEv8b0biju7DdoOINTQM7tI2x6kc/VXMT9eWk1rngEuQFLYe3g
fLqCiwO87o4fCYfDnkvdOjW6+59WHCF9Cn0JwQEGOPpGFyQJ/Q2zLz2ycblR/rvd03cyj8TFdkCF
0TQcK1lQ6TjOo/K3QU8zWsBjXP71IQAJGfo4j3kJ7pF0ptB9RxonEYnVL65g8H+/QG757EvYDjgX
zFfnnkdmuwvAuXBaykVjFgDa25HzOsaxz8Ht5blNmH8ysdi5/hStk/ZO6zElznvCXGScr6CruNGe
A+DgLBx2meNegGAvfv2LPPoPEek49WbE1eTce3jP+od1t1NyJPOG6VPwctUaul4Q/mWXF2TjTiQ0
HGtkBmq+hKkA0PQzX1RF18W39pkNXG4P9W7iEDPZTGnqnB6+DHxrhV6hMWq6TeoVVRvPnQGHzVzl
uvhimVTrrB1bSD6N12kFcoDKK9NY7xSLoSomBM3dDe95X82YwmhqsvcNp1XEYkizqgM4zevddxJg
VE5/eCHhg87Cmiz71DvFtFGFRu37Rbo0rlnCDny+mp2f5zOnPu1kru6mMyIP7l7yVrIkg2HKNeuZ
Xa35elQfCJXII0dIZnF8lCVaIgtY4qL/VHz9IshVxSCzcyCbudVf7282Dx0YnWhgArM7O9Eu885U
0JwvOIndxJBcq/BECC2Y2VzHT5iDi58JLT1ZiyZ4FyY6FX1nwD6L+EJntK058fgLEKXGBRamDlLU
w1KcvCPjLSuvTe4x8Y49MyUoJDkf04Ek7TgHb60S6rlwhAI23SFmlEJo0OTbALUYO767OJ9hhmw8
1HSv3gTW8RI0p7jxrKq4ml8o9bCIInGASKxWZ0498WTdB8hYTo4MuAa+q2mo5uNMmbP3EW6eggnX
VMu9sBYvkGrKcrm+9edS25R3Wyf5KnvpBcSsv8TqH9nIxsGMn0VALX783yGw5McdNU8cFmg5OshD
CJyN+3D2xQrQkg7t0rb4PEwchDlR84X7enfeXn8yRwdbuxL2vdj0AEFPXo4FQPhFYXM4uX0t8Qix
dZv2s3Agk3sJ0r/A2nOUEZyoDU0v21EQMPtVVfPb/K+olnB/qWqpjlylT8Y/mIpbz3+Vk5Y8CXWJ
qx44mX31IV8JlPjV+KTamdxeQ8B1orYgi6nDh2mHl7hRgICpvQMXxwGoQiUIHPoyDg1jPuDT030P
ZvXAad/Z7YFu/tVI7NTNLcEWMUfnoOg53w2QqvG9E6w2DoWXeu4eiA4WFO2BeCjYdg7pECTSV/3s
gDJA8gBcWBfMYsVKuFoXQcXc51sC3ZdFzj5qFtveqvxMs7gVkYLq3+DSMpGV7yCA7SuhUDvgf7Ht
L0IIRKnamx9KAGuF4T0vMm52ciVCP5kmhnSnEqIylVjIhCdHKHaSXveePBs+MJDz/JDGuYUdE8jI
Ud90DPJeDv10zqsf0iH7tBLbT7lhcEwoZxJ26RPUdQrvF83CQeFuq1MPBDMl4j5pSgHWrRi8FbgT
RKua5jHNXKGya5cTreKDDeIa+MzSHesLQFK4RaHcPzC0SKuefb+Fd9fga+xMEtFg+fmuZ1vGM1NY
C/1u/ZgQAoLhQrNB2g8WwqoP4rAnCMiiJgeEYBLuU6PtQTgRKmOSqCW5QmNpKAaauRAf3znyid9A
T3c4AXkM/Rcbf73uDG4KAg2K1o97uINZLqDSJtqt+utq9VFGAKahGdkNL4ChuOKH4gzdVsXeWiF/
ItsUjGqybpOjHwTpSB2PZq/hodWs62dP8p7K4e23bHU5koY4cY/dDmDjgimu+SI6bo/S6wU3zk/I
89XjqKqEX40cdVZ0HxYFEVczSDhNA5pKg9FEjhvDeZyYPPLf12IrA0n4s658bGQoMMl0qM5Cob2I
WF5LiJTJyFkciBLJqwjj7C6mHayXu5BrPpwEARHxdlfhpDzKSR/y3cT2/2GiMxqImctaA+XRCPBN
OEi+OUprEEiYtxuQyX1Rwdpx72fcGAXpjCT5KJk/cYbxk+qWsNH5i/axZ4djtMwHiTqtRNFCuaNu
bvsJ7LHjp9jDDwYs6D5oX7VZ3kpfItYVgdphTVuprAxfb/Aw/vNRsJxT+2ZT+iF8PiTWA9oxrM8G
TQrBMSitE9CuBq6nYOHUUa5e5mM4N9PxwE0M0U0nwFbe07RRZ+mvlPMTQ0YPEXfuJ2umwZ8KKGzW
TThoIR9t6u8U9ebCzAOLEL9Y26fhHplf9dYKZc8/hFUrAIxyZMjgAf3kaW+BG76JuDxTrJ35trGb
OdY3cXgWZ4rciw7K+rDSbAxEkNAUS6y4wQDexAz/4AcAVOvaGDs0g+KDV5elqI6EwEYT2zAaP6JR
n6mANw+ihnxQ+FwXRx4bCWE2tNTWoIdOA4l7G+adeBVt8rPerAND9XEbLcwsR6RgaMc+7Q5iVzFu
CmOaFVMQM/Gv4rD0VgRENNrWzFnmQNG18blYwOAI47IM2swU8lmA6mT4x+mFpRMJpV/fgy31+4M2
C/TWVjJE/rHMELuS5w9CHDhk63ga45ymHZSf0l0zziV2s7bwTj7QTHfgywnojgnSEDub0h/hAiXk
ySxoECZ2anb3w/hUpGJ9WK+5ckAvwpPaUy9gDnzceY4USKQNtqAon26ExcQAYXI07mG4IbQM8ffz
szd9Uv98uedh4N7IHjWbSfMRseloGwoi9CXOmxaDh7A0Cr/Or4EtNoWIClSSd0YjENMMDodAm+y3
kP5Gtmk+4jzFw2f7jnS/l1ZbuavoQrTT0gj75feDqAYtLteEEOhCVPJUBDrc78oZ7jnep2+OdIsv
nQcC2auFhOtC/8f6re0bYSlWJn/M+ar2Pk8eqRYZuSbxAiz9Rv1KMs3Ofe+geceozsIsEOy6s1O/
liOTqK3QGcqAdA4A8VSAridqTZ6LAoCH4Lqc00uDRUlWCaIbMFnnPklN64Yi1QyPvu8XNf5FFs/A
OOSgmQvYkAZWFCRhXBaAvTidRdBqh3SUZAeuMqQvWaxQWLj1E+mRf2L+mhE0fq0k0vkxecoNBTx5
aGnyOKDstwRNtGl0V7Oi8TPbwBAPwskzFNI9v8cGji2cTm9FdVVId80tZpYl1Pzns2zOYXzvgl1d
0/julSQ4RRiabxeIZUiGoqAbc3SAEINIqruLQ8OZH+t3R8g5mGfg29GFRg2fGOQ1yBBEOi1F5mpJ
ev93uWSG6b1xto22QfYlbSWoCbskMbr6MsS0MJfRvUZUAi/w+ndzq22PwE82wm4dJKO0hmKQ7ZTW
54Gvh9/d2F6nZZihFLuL6aOF+JsikqEmbhGDcMR04CIVK3h0llrEJS3+40uXjhFLHKRi12AQW4B/
AqWwTNnt3VzY4HxrykAmL+NnVD8PhtSV3vXeqFST5f5eyRl7MC9xKGp2oBo3S5B/R2+WJ1a99l+U
ZbU6GSX3zCUHWcCeF05CCuMTr75WAJtapx+A9QTl+NwBLjvrAoExh/Sbai/15GRjZRB7tb6cM/nO
pIYPZQ9OhTJuhqwViS+MZ/Sk7ODpvvFaMWdNLZ699oAra1Kf4qVwMFaRjTsTuSZCCSUUZilZhGCL
h1lb9OWPx1QatyCFzIR0ELeYx/rYyXTU4LgFwTRZ7UhznWNjgev8uPrXDFsXf6kByI2aI3cr5WpK
h+RLzeulxFg+CIDYGuNgb6NH+Ky0iQnYaHj4kDBNZWqDKNc+rFWSsayB4TwLVA5+6VQo9O5xXDtC
sGlnjuQv5/nxYhsNuL3GL0bAVvXZUFVjRuZDyo+x7/I41XP6CC7ej+W9RitKFLb2Wf99sVljpbci
ljGNvsEhUmui0Iomv4/4Yt+Ji2cxh3FHx+vdZi5N98pIqL36k/NMOq1aVHZVXnbYgzrEs2oM/0Lz
yRZoLxBVhxxn9mvdiWBurUcD+9ECfvkYGhNfaw/DE3RdiYRec/UGUE/sm9rHANrUthIHInWNo9jI
Z7YnN66wA7dUzlkYfbm+J7p+UZZNTGPUoNFHXSSGN/Y2alGnkgC6TVXBzWfmvNKmCeKhKdYbtQgn
rpPevy2LqT5VlNeOlrEiWEZy5kcRKLwf882fHLgdS1BVL5Uv3icnpZADTnOM3EoTXwme43sSkqvz
vZ+drZGBVc+1EBdy3H5yUJ6n26B8jw7i7OiblwM8bfS05HEiXKlyppSliSDmWUPt6GAgJ1KkB8DN
prTtWGrXZSgaxE0rT1DKUFfPDfXq8AxXtR9PDO47jbVbZ/3n0xiCGdYUKJwN+Gb7rhFhGYMSHgZC
OQRUJooYnckApvbTqs6LMdfVzwtRXJ37J5wmfEoBvK6Ll2uINHUCbVC/u2ovl2vJ18YiROxL6qNN
Zw7nl25ofm874KjRXVxSd14RrryE+jajOZwBTe1GWaZM8pkdNtlH9wgK/L6a7x6brVbAoXKtlnfG
umrGBmXMtGy5Q5VS6zTj4LSYWISZ161Rns4o96Bmm+oF0gH8S3GhO//6h6KNu42ep16oXXrgPu2n
QNUChNfe1calMRfwRRqPgdKDWrUQEjJhUiFTBmxlNowsK9/gJFJUNINyMOAQmt1OI3CEqb86FDqJ
6PgnNlnIOpyvZDXXj/dDUBvEo+8+UUPlNEP6tKzgEH3QHZJ9vUxK7pqmWTDed8Pfk+SVpfStp29c
HxfQBpgMrEUlRruKLLBWPluXagxq61OsSzPFzHVy+Xg+Vdm+CCoE7f/q3WJYebVKAFXm3OQfzIML
DsHTHOxAJ7vthGDMo26eanIyRPKICuRMYKM3t+V7HuXpYI90VQ+0hriyMoV46xx2GyqLKgqcWOq+
K6C1YHZaa6xkIiIXdxYm6jtcuxzeyG8fchVi3cLqb4zDuO70DLwTDKqc8YOYbAX2ZQOLqfdurBja
DYoleAlNwJJayNXBDKgOwRupN0RGnbLT6yBL4DzVQsI8DWAPd1+lklW3mtu9t0hnnTvr3US519im
boXKdIcAWlS60MEp6ZMmGLIIBwa+A4rHw0ViSo1ArFQ6WuT6eK5bb+Vr14VL8VPwUdc0A5k4KRmu
WIxpxdOJYaDIEnRLAlpcHJhYqhsa8e1xH9BRUCMANCdkTJs3jsVFT22zccjh5paEL5Q7n6QeA4J9
BpGserxO1Nbl8eARspy1WVdf4AfDI4wQzX0KvldMuUDtH0GdcpBN2g4c3swf5kRw466sq0ccd/Fg
wGo1xNtWTcy5AbJO91eTdIXmr7gpJa+LxnwMwvPLB/nS8YI1LtEis0Gt+GRksrWe+305UjxD4EYr
e+d2/ykHj96dmHOuEwZ88/LN2nCIxuydP+YoePD49NVz6cChsKXflkST2LQZu+hrV+XeTPHWXHyu
4J1fE0+76sd331Ev7q+Z7CfQyJ4nBc2k8z/r6RHFfcEVjKkcqNKCNWj7qPNkfIwt/VtuoctoWxmd
cZTwd5q0Nu0OmruwtDBz6uH/5lBVhDBL6bTCF85TAioFLFdx9TGGHJx6QokVPb51yyt4JA8Iz7NP
uGiquD9hiV518rIuJVtsoNFSfKaraZvPBxWrcJ+n6G61ZdmxT4jJ4oIM4BhHZASG7APB6Poe7D7G
prOH+khH8X4wgaKbYefyT8kQh3D8fqIpzy+hzZTb7FD7I81Mc6sP/yvRDXvi318HQ1iOiY0Lzpiq
nsleqxjjn8uO0PO32kW4IxU+lz08Cnsa/pKSb0LFzKx8uKNR/CMSi4RU+pZ4fKh6IRXrQQvlyJGI
DLOgeMyt5MTuAhJmthKtGbafHqSwPr55r/nAsic6Z7XabkiSnZTZdgUcNGV7Jc0QZb5uHpRt5dHX
UAUGOPHQr6FcIrpFsNnUcqGN6TKOGTL9RyLY1wqTMVDUofhhB1dxP+FCCdiV9pjjIyKAZLXKXEog
H/mVG7J51yto9a69kL0z8L9eVmOwRrn9ZpCDLmIHXUWRh0PO6aZVl+/4zCLBkeBq6jBIerFxRt7v
EMEWrA2mM27zLHiTQJeI8wRiG+Cak64fb73W6TfhP8Uvb3ttLI3BXPbeQvL6rG8HFFqpcw1yLMJt
sxjiAxI2SJO1R966VSvJEVJVxa2H4/m/0PiG5eiECyV64TZvXWUHcz2tTIoHUEv10rE3aTt3jtZA
9RflPCKQN0PlxTogCXrqfIN9aBkJblchR0wnaLB9G3KoymKVeKuraeRL4OClk+L3UBAROGU8eSIT
qllwFNTV66yNoASqq4ibgNJ7fLas434PaVz5Q4qjF1MbtRuovmdaPC3Ok19Bk2ApTki6Cfh8YqxJ
aSJOgM5zCM7ISI/hZ7PwmfN6I/cE+N/+kVD1TYQwkXopMx9J/6u5SWdxNdD742oM/V228nktoXGu
XcKtUmDMjrnEdJEMtLn3VtcwZbfev/8t2XOfeV9xLJKbWPnZNsjhLJraHMHsfwRDr0L4yx1Y5WgC
HHnCMrYg/9+nr/3SxQ53ikj4jUGN3ZsKWwYDq8aWbMacUQmqS6oAp7xR6pZpWDDT4mO/lHN+aLcT
SflJ8oDOnYrwEYvks4hi2DrJPZ24zU9W3wXHmJqNNk4siIfeyZ2ziK9LOu/uU1qPm586atuYdAvk
lGCHEE1Ha0p2eezRW7N2FvNOCr0B34zM2/Zw+6IK2gP9Wc0U8JPi6kt5t485Nn7eKL3aQJedrWjR
fNGUho/I1v7cSW+DbD+V9AFTw7Cd9Av4x5cbdUOkzjW+TJPrVgMgC01RhhH2kn82vHW1n4IR6tji
h8AI6N+4s8DTfBqcJggLKrD0CSkVYYFo4VN0rIQhQ4c+hN7RmPlRKaBeelZ7E4XKtHcgT+PgVQIw
UB+DZQsUMIrJUJ5tVAwfClU5T+9shiiHS0xPHXRo89iOmsekJVRRLPj6J0yIdSW8t09mP+ID+AD4
MR7O5MsGXUSYuDtjDQiSv1mVIU0Ja+JrnLHdOzTalX/D9w4nD1NohdLza/29QM7riuF1cM1DbyFN
+mLGdJ1wOiNvgbMJqfGFgLmMx6ua2HFRh39/yljg2mG//WFOcd5yjcmToVzKVj8U7ingQu5lF1tr
oi4jHnwqu4VdVU3Kr9m34ebpsCPd8/nO1lCMmiZygyTQ7/KKkccvQGJVYNQO2kg1a69Vqz3dRA6g
DU8yQV6JJeIaT67fx5VxQz9y9BesGFjrqehVyUBGbXAfCmSpkQwvVOSqFoPO0DAiClLROyRYuRb0
m0XaA0tq8A3EFjJ6ejrwhZzAPLtz0UES6buWz/VUsTP4FMXkNvcdAbUse/FPf5gIVSVLIBaaOY/k
GBgeUqvb+4PuQJzymm8itG0gcToVmagnXhz9udYb4llVDbl79wtA5/QAmJhg3nb5/C7sHTxOJhHU
obHSD4BnurgCna2TVE+p1B97kG/Q4sA6LVAbsO17HiYjXw9mFvOcftE6YK3hEM3CkUHVm+7qr+5w
WotgxyzD5xXhhdyjSgwt00y676bHSQRcB3s5vhdbC2OR5eCPUiKmfZNNwFu8lA9/YagyQfI7zsou
yAzDZ36Iz7Ey5NDh5rVKlEQDbP75COvQRq99u+WQhc1HMxCMXJAQ+tIdXG5ImOk1s+qeRxc6kKhP
cyGXPW3e6aTFPXLE5NidxCGZLvujxhGNYNbXxQbRz7h1LgjtLc1Asi9dxM+aruHtiui10QnKf6fg
/JQGJeEOLrezPDnIYTCg8//tj/1jEGRZ4BBxAfQFf3XTFGGu1gOm+KK0b4toQIw8SLfU2hJmRV8Z
P7qMsGCGDsKLLHgZVQsKqR6/93e6eHCsC3ye2fA1MQxH0RKvQl7918sVABAcuE+Za6nl+0zQfIbN
D4zPAwyhZvRWcr4gw86JvpzFlrP1hjm2kPXI1WIxG/0Hh7rT2miarUeZCx6PAA5OMfxYLlGLEmvJ
8sXMLysIYnwkfev3ipluOXigvIA+LQS1nDwQ33nnTOtPX48D49SV1xxOMwCxJaiqq4mK3sNHAvvh
kF+Wdv/8u0+WVSz9TrtoQ3u2Nzq2NwhWwmXRyYURRIN9imdJMIjeCtT/ObBokiihmGvHWNIfmkzO
G/1gwYEjGE+sdXjl2svQaMUOR2rsV32CzSCSG143Z7xl586BWzkU0bNZ10sFnhW0zRa1Uyz27aeM
ACdFRN8byeDG5z39xEeFfoBFXsR/Bx1iavn7CnfpWAUQNBL7NeMskaoRAx4KC41OBzZHc9rvoEkS
RmbmDoyxMCl/95tvfCrWJQByN9DehVZsWyRzVBA1GRsod+n5DubWs29SwZf7MHryfzdbz+tgLaa5
BTKHJb8o++42gfozF6K9CEOQ26PfQbXAmkI2x2XnmApd49M9U8k6kbyuY6wMu2AysnDPMSWCYxqx
CLMXThlrpTxsWRW5wrGhsqgdUevgDkwCq++fL6dmHdFvkzctX4ndIaYGAGWjdRpM+xaojygRt0qZ
enngSyhnSwj0dLExUFnYis2zGuFebPCc/0e9Pxq/KHh7TTWqHvenr1je0Ml2HSXSjKque7OwFheO
jsVVtwHhra/NK7vJpddOwWevELwfqPNbE6s39eMWcwyLiAHca7Dx8mA4AyC35jufZZVCE8EO1lP8
ge6pIpBn0rzMvpTnIq3fmwFCJPuF0f7Gzcjx3xGIa6fdEBL7bOVbgXQm0u3hUQKGC1o2jjc/tRcQ
4ZBx6Pr0etN8PLgy5CLu3AEql+WYrcmCvk3MDR83SonspG4TlDMoFnzoa2d0xin3G9f3b+UVlmRT
oCBC7vu4jRxmHh8m08m6GtW3UnJnSpQ0e3jmWA1FVRIbECW6j4LYLcKVj7aG3lGpOuEYHyG8L2kU
Lgph8CCW7wtwydwBOGpE9S6lmm4oyP2K1TV76bvmI3GtpHJcsHZarD0nlVdc1UT6c86WDoZ2cSwP
oeBvy/JFTWPyrND+3nA7EnRbjUp1B8Wh5FG1fno7s0keQhg/tgeJABpfMYsFz1N2a1FC2owcHv5K
zp9uayVVp96eoq/PgEpMaGauBhIZN7YcyBGaQpN+urN5gXvslrzihey9fvj5J7LGV9TVz7QqHGwS
WOJlo0iNGuP6nQEigwHGkLmsMvZMLDW6Qxl5YdcA6aJLgIK+W/2zwiblsgeq5AOomwcndocqGSf0
2OHxldg43pROhgdhzvMZqaOyEJcdzr41/exSx/9lsqIOyAvL7CbRaetxtASOZ7CddQ6jMN2PPWRl
ThaOJBZwoI/cZUaDj3RHUvAyY+boTIcflRbw9gKI41bQqITMmlBuYadWlyPNUU8mCSZTM8jiboua
QovWWskBiCBwRKAjPVW6Uly1MNdJaNHli5MYygetPySt7hUqDJq63f5mav5/ROjJMcYjpwK6HgP5
ghqNCs4lmbPYOOZSM+rDfQXvycgIyq8lv8SWa+My35WNTxaV+n7oMvevbd84bHj810YzUmT1RfBT
Wfjduk9W8v671LGPpI83wB8WhN3aN8DW/+ml2Tvu667AWJGAk272XDCa7mCtj08/P3ocDaNs3n+1
UxiQtL6pfo9119yL5fRztTLxVyX3fpDmlfhgr4YtSpkiz+iseGrbCb3E1wgFN9OFgYSPAYVd9i3E
p6VpZnUbS9u1nG3pGlOTyhpSzlck2ljhUcSIJ7GMxz3AUyvjyB2gpM+8ZR8UF1GRkeR2hc3FXNBx
BfCeSM+wd1ZopMON2ceE+526PrkRwFwCpSHVejNisdBByygsU0/olcAzvuwuzg4NFgwYeAHRm9pE
PLWj13dZW2HigktqMUQbv+4PnRlVG4j3TRdkb1AnfTgvkFIGUamKyFbz9S5r3IwvaTPm7Yfoq3Ad
Z+eTN4bgSLMprw4JtPxoJkcPkuyq+mDXX2cHivbAHuXhyKBD1bj8McKw4OgDlBdtDmdi7Vgp6H2L
je0xKijqJbSOgMU1tk6VfVJ+i4G1urSTG1ZFjET+Skq5aj2edTU+/Us2ymotKmkPWukYmW6eLlbn
HbJNAoNoEWX8ljR2oZ7i7ML40RXAQoJxw5AQ742sYMMxnq9C7X3L7mYDZBxT6TOKOy+EUsm8mVSk
bjXebAuesV8Wu7HbKcFTeca6gaKV0JAPIkEFQyPfWyxnMqFdApLstoRDL5HGCDTFGv6eI7pssXg6
q+LAUI+ZOGsDoQmVKyByIEeo7PEvyRWrdjc3BoVEmTkiTkMx0rUkJcThwBXTFeKshxHfsl4EWDdB
2q8Ra3xDda4ZUTnmX6nLzKTzbAoPTwlHu7KrXyzV0ztPbT8wMPS1foH+3jntuVYxwvN5NFMGRrM/
Bn5/fqwg4Ta8vwMVt6IAzybwmozKyJY40vVBsnLsqcsvVOhq20K+nt+gTlfvg+5omOa6bC4TM+lS
3xhjHNe9z7O1DGWM2VADbskmfM0FGmasX+nRohxc6BXEMiTk34+lJLdowhzqyoL6lLTYKCWMTtAm
A0bjhnzW8fuKFVCKxk6ZHhtLgJMJ2Js6Lky4mp7rmN69sbjy8cU4i/gBWhfgof3JueKbL4eOZXcs
b9FkY+YrU72RYtEd36RgEUgy7p/3U1aX62AurzNnnM/B8lfaZLQeuCV+YstJoIOBaZU++bed94mG
saS0KGsVgscKX/lS69WQmFiadNsVcMvE+uk5JN+MUql+lI3LG83PZmb7PWvzGFsiK4jZ+2m/c9jQ
aQppKG7IuobjzauJtk/dpAkMYAqQZixh1Bdik0XyppCK3LY/CtGpBDqIETcBYUFPVXjD7hrQkjrV
MINqotcbKwt0qmArPF4yHssjJ1mMowZlmMqo+73F/pO/JV/nhj8h2XYo37K0tTn704E6LW96t9Lp
r3lUW//NZ0z1VRG6xdr56JDdZ8yRwTWOmEoMTBkB/+9lCyG1dzjiROzeAr5JAQIAFIfijcMiBQdW
8yiBfbxqslBNM2qHE6W8o6tpi9R7kIGwiEjEIiyvimcMVY31BEypGbP8OJoFmXRZGx0p6wWtKzpF
JNIDIRkAo0dI1PtDgZjXDHzR6dqtW5OJFe1hM82KGbonCg0/iTh9KygQc4NENgi2KO5lJJElyshc
NaI9MSrB7LOfztm5zz+fi1zsdKLA5huMSdzZazF2sheND97eM8b/CXGpIYW2hUsByOasRlv78hN5
svTmiDD2W+a2NCKdyc6I51Qnmm3jnZnfQu7LMpeMSNDhy1L6rKJJyxFH9H1g81sQdyExlUWwfizM
ECV7aGimkt4UBLLbkyeJ0kURn8GjXGJ2hOPjQb6aPsguwZdhVLDJdWUD8W4sdK5ED5SjwlWh4qHk
uZDrgNVeUunlvL1FGEw/dL8hBVHcS5oiQrUq2r7WcbLK6OZ858On0HQYGA1utiE1/A+TVgfonmV5
u0o9f2+00tNOa9StWcriXZ2QfsM3R7wzsluxz+thMmodorrvKumKg9/HyAfFbQuvYQs6KPPTpkv4
o+mrTUHBXg==
`pragma protect end_protected
