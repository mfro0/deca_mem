// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
H9nzWV9nxjl/FlIX6jNT/qHIWm4sdy5d7XAC+VnDNQW0WW8Mbg+LFBPIjgtKoZXu
onqN1DqZOtVZB1753cQ7HarjCkdmMZH/DF4gooiK84YxMGHJg0ECxLt88+c9bAFO
olh0N9Kk/u445HIkt7MRyyDZ9FYgoZ+hC19RP+XDB7+2XbvBGVgZ4A==
//pragma protect end_key_block
//pragma protect digest_block
BzmNQuLYRafE85coelI6mDEjb4Q=
//pragma protect end_digest_block
//pragma protect data_block
QUpOHSVUuYT+ZbifP0UpRpg87TeN+ftOZ1TIxKzz7RcRjw7ZISOU4Z2zfBJr1fCt
XqPzJ8FcMgcWIh5sPIdxyrn309aHyutiqshMCGGof4lHN2MQCb0nn4yBBg6InWw3
cog0lp5TjTc3wmdQs9cxg3TEkA31Kwkjj3eqSLZo08okdqLQDQMvm3sPSCXfXlwU
ffRN2C6VCL/uRnUsuuPA7G/0Y8ipJCXv5NNx9QLlEHz+oZFHnKJuKtIvYvvo843t
3gEWgrwrws+azNgW+/g4XXJTwu2qGQPKfRrkRfbmCCZzIbD0RXIK0Civ3fHDIqH+
WwbTGLu7rMwUpRoIu5GDD3OrtKh+Sk3w+k3xHKWByKpXRj/mdjbwwV/uyx9d3BaK
7LuOF2228sgtu2kZ1fOLnipa7JVlStVe3ZFHKJSAhGe4D78IKqappKfOzL0vSNUY
CdzOHrnzIKJtGLBPTyaQrsS4erPoryfAtugbU4X6yHI1AebQkHUQTCb7StcGA6Cm
5ut+dkGgI53YuzWqihntB1s3okEWN4KroQl7JOvqwL4Nca31SpZd1aE6mXWXRTpA
DU/ZsFlrt4qZqNP+1uWszpUf023mAcVQ/gYObprqEaD6Sv7QtSGjxNJ7MjlWz7MR
ulzsqNEqYZNqZjAcRg9cKffIPBZcCso3F2RcUZfZStblw7meYxrVuvXBaGRlDuzT
cf29/4m2WCnwrM1xEzBXI0N1eu5LqgL0mWbqL3axXQ1tpbUxiRuHXtZ2zOZxSW5B
sRmy6KHi9Kvt3hE6UMoBlk9oSzY5aa9HaCJH7ZykizGLQpOalbVYW0kuCKA3ZyFu
zMYTHL6nvkGE68YseDYMEa8p2HVL0//GaIF0f4a/VXm8fRTsv6SvWtlVwlgSuBeN
qtBIS+/E++fmVLNS/i7wRN7cpb4dF/NgJxCY55UwnbFyqVmewD9A7TpGbyx2Oc0j
HPSRA7oFvLEoeNFnAohoYcBdmW2TLqbZwAZt9HBwinANwidOOnpHzlnPPHBA5ElC
borQU2H+eCtgSrGvoMbzpnWPAZfD2ZaFnh3iVXlFbU8/fDNyBiIbFO9cb44VRerd
EghWUeehIiA/qVOPpQKxaPu1W7BOm+XsNaLTQwEXeil9nKS3xSPiNzLmQVFARKVq
0lRaoXWsGuP9TgOJOmP6WItR95nBmlgu/mkGTzpXlCrjGX4RfxVr8F9AreK6qplO
gFgQ12UOXsw0LM73vfBa3MHmEOX2rxQkGjrtqOdWxiyjLYbzpdJ/u+NUcjScLuNV
j421a/INKRearyKoxOHrDde3jy6esbvlq+GcCWjIzi+QPW6ALiFGWES5uxqi+8ed
AjTXa0/IzmSczb6FrRzYr2r1DgXORc40WP3CTna1/qQNpRRajZ+ZiY1R2JFhC3qe
05BZ+/qv8jyOdaRd0yK/E5Iza53dtSFXjLWZV9gJaKbwot8I1i8zd0fY7wZlDo9I
vilkMm48YgRFPmw5N9dkCPunP6/xEKZS5mJ6XDNYFinTgfWBkBCE0lLYVPMJWPeJ
Jyq+kYe8DAsSOkd5aQzmBfb9CiSjDRg+vqq47S/WRWpo3b4QDFredPc0SYFsxorl
DSjqBo/TszZqejoaqZVqW+fwRTmjICP4Ynj8VbLEKYEFn9Pc2wOrzXFXyCEdzYJ7
Ge4ZQ8tYS92P97y4fhUQ20vusv/thZuJlCwtlB1EiQu4wx2n4R9oU2ts6USlRWw+
UVaotW6FreyjyoZ6oL3BZpwgrA9VjxyX+LyVcIlj853+nmR8sxAqfSERhGUDvV/P
uNxK/+RMKnqPL92EU/favNdfGNkFe2lrxdvsov+hhv8BbUB15E3nBBx3XwmQ7FH9
wrahoZ0owwSZuwYmrZeMG7yTH2TQ5XFtN0MYTgPqc5L8gzfGNPjJZYWWx23Act3X
RkxYyFbtkO3dLhTbljF20BG5G4Dm5+b2DriXzlQ17yY7ebYBlSAT9WCHZaCYyvnD
SeDmBnKX9lFVgBvbgibQqVeCZ6eaTmoaLcBhLApwCmk5fo4C5WkkP8Okvj5kPwhB
i4vmeIcrJLAhZHlSD5n391lM8witcrJetFcX4e7D2aCciuHhEAUlXQpif/UyMCkU
cZ23LQwu/5v5VrjHneiJmroKFUzXYq5O8W/SmtoeHazgraczAmHqbEKy7DJ/3sBA
mav6w4k9sHgfoC7o/A9r2wzgqAJYEiydWQcDCo3dVsSVqAUN88i49Nga7Cr630/1
pDAHUwV9SdPohWoXtKPXC08cqQaxYv3wiRJaAP+9DMPakNS+raXVIvZReC0BsAyr
FH7+pMUJWbrK2LxUvUwjuYkc0YH1GLAA0gA0+daGjBU2lRw5XtfoAn8/SwdnRa0C
Hh/IDt4U/tBxGcui0Sm9ZM9BJTFwFMZT2e3qq4XcqcmbCyeXmwcVq+8Bfjz9u4MP
IPcUnRfG6w/O6VSLb7B30ppHWp2cTAVuBG1EiFMRR4E+lXNUbApXdZhemuTiidep
8zSRGd/L7G3YmjkVxiC3jySJO1369eLCeo3RUQLk4DTxewLApag8TrckKCVKdg1Q
u9oEDtVKriK4SKVoUXqKjzAT8MI3sn3laABh7AQZ6GbuHhor1XTyS/Do8Mg1d4Ge
cFhukudnKPzLvJ1cx4lCDqI+O48K6LshSxB/FY00RiarcD5l4pNkQDd4U1/GcFWM
FqNqCjGVeoir9Pq6vtP7woiu9bADZL3ZdRR5XrxJTQWSz+0UtME3+T/9XGqnxflp
jbki7OB3GhTxUD6IKx1S8Z83XBluRwnGIxIJk/+nv8+H7RUarANZPfFAf7BnUMf0
8TSsjygFqEeixTmt9kSSvo8dbFeSEaViS/6+JIusoInTJ8g14ytnaUagMjhvZISG
wjoKQsMgcf8fVZgGRm4Y5QlQ4ZHmJLoQSsRiNst2TDwp4XEEPPjz3qgkwXHSJ+SO
SwY+ukjq5q56Fq3hRtXKyEHi1b+mkQEhq86psI5XGwFL5tQtfwNn2hCC9G51u6Bd
0wnJ6O/J68m6M/9V5c3YwCib/SHxWGQv/8tPHs7XkXsJnVZmrwfke6Pvq4qmH7TN
5xGe9NrtCBbWEJJ9Aa8v1yBVCQ4J3mdDh0hcSBsOhyDeEf8RjkvUgDHFU2Hvufbb
UvawzRQ3blHBSY80tCJeISWDcdDGIpr/p+eP/+sRiJFwqWVWmLQbWnnkK8bQW+sk
YNJlqxkaFlV2y8H2a7W1GqcSyv5HgDVNhXQJB2QglvhYEoqlk58vlAaQWzmZFAWt
Ac2nm0kMlbDPM5RQ3VQAVQfa4t9zjvm99PefvwzCykCr68RdJm0OBhFwe1TRuogs
jQROABknws1sChxdvjEGG1pWIbDB/6WGhaIERg6M5DMHBpFU8sw0i9yFKUTo5lkk
uAnhXdsEgoyN2iLuuMhCrSr8XfOOMSOgZFDAJJGH7B/aCC7ifpYZ6icMr/72Sw2v
bcJKkH/TlP3zjiY4txyoKov37yS+i6tqVLhz9CIvSU+Q2uRUdWHjLOQ+qdUJLnxB
TRXc7VpnpGeQBF+RiRT96OUINh4M/HgFo4eHoLVXHN6zsNXhs7HbsorORYuRPzKw
E5KaRLV6zrGHZs3UJ5VqnpTIF3jIN845X5lr36wqa6UmnpLTsqUs6Vj/BC5MXSr6
FND4s+OTNHg23RLUY+yymfpo/TRroKA9mHCGQJrqeTVn82zH1gLNdP2ZmQAwguze
JUllM3ZMTaNZRu0PrNLG9SLsG/T/wsNDwhgzAOUXUkB7HJnaxFMCh6znLt+yGOsa
K3rUKLZvzine0hSE66aMADbYboXMHSdtx3ZXvKqZC2Inh+1CSYZgrGS9yTcmLJ9M
kzx+YnUC9PBblucPc2mZlNtbJ6PyD2UY0VzqNZIxrQGRiGpR89TxRF0HkHLKZOfX
7+4D+c52ba0ZvhNF2+iq5fH0L/vPJiHS2ENgGavAuYFOtlEGC/b6CJuK6tENnXfT
DiqFNlZP0j+sYYHM5hBonHR5amKTN6uEKnPuTisjHmuUunqhFvW7qTONqu/KbRJw
ouJpiVqtQ7xfLchxmvj9/1wYOCpNQ8D8NGVFThDqcIyMGbJgX+m2I1IiIq5SK/wk
6NAY+obuwtrBrUS6EMYn1wmjp6GnLn7fIzGA5CcTqhS6GZVz8B7MA6qr5OhfilQv
KzzZ0eujebFXZSnT5b9M9EWdUNQf5uEUw7ysaqDHqtsuAo3G7BEYyAHYzyTrB1iv
eU9hcWRnkQOLNjZH7h5QWnIrKzDZAfsOZTSDPH/kfb61S/l7GNHq6cZ0FbzzvxTV
3c8mYJ7QLZZpohNYbnI2Hsy5d5wnDyNzgSyyP/FmYh2WTIf6S5Qzi9PGJ2RnDxQJ
omQPohQqOwjGcHcGRpEgsJ8L0tbAocQwOsp3uQw5lBMn8Hb8+5yEbcmoAnVFi5e7
twQoeyDSR+NW6C7Gn210yavCL85mrFsqAJZS0nv2l6xxHlqma+sp3CScpFxIldm6
ejkD27+xqIpDBAL1wT+g5Whl22ZI3NKEOD5zXWE/rnfdf7UgMmqzxqWR+2esDTAx
lsRoKRm5D92j2KsPULScg1hCTi4ANECkUhCrfPNidE5S/OKsuoSaW4npyMN8V0vi
RLzAR0hAcK3EGcByw8n6+koThFeHCJCVTLeuudeow0KVIDK0PCfERq4nLQYoiY/N
VsWPh81MMKxFAh+s5CkK6UQD4KFAh3ChSSYNmvyo9r8VN4P/7l1lfBKAYMYSv76l
F5ug7useOhgTCAhL8xsIKCAJbwhNf2WCrxyO+MpigyrRRBQVfdyyxkcy10d8QjUv
8z9etIpU8W2Djj8wLte2BK4F6fj2RLDuSeT3AY2y/yC8nuGvq0SB9hkae1OxoJ0n
V5FffdLNYS2lIofBfA8p7u0qf8Zd3alN1kTeenVG+s0VFaNUI6FM+lLo+CgTqxGd
0ZDDNEoXKmiVvXH9RMQpuw+2oCJJBHrEJiPwATzNwa/HX+K0WYMwUQqyl0FIJWfG
LmGwFTrCiUFhIWfHxzMX3wFxBpq4NPGOXhmJLqz2BHOzAk6NNgSsPSwu9x2JA4CK
dXGdGEN3uHTBZKPy0ZgRo9umv4H/2pIZTtyqFpdJSFR/WDDpI0XQl/5x2u/K46L8
dt8oOBXWLETlyULjZPBemG9SDLUUvAxsXWJQmHeGHiJGXRgu6YQpyW4rdFHiAAC9
49Jb6gVAEYXVEYud+uuyuwfO1Um+v4R0kvLVryv0zhaYW8aS4qZlpJcC1mFv9CMH
GfDQBSgJEK0r8HLPpJTtM6L6SBGjW0Zbmx50ze5ECG6xviqMI9IpI0yAfYWKqiYc
KsdfUZrxRRdpzMsDUDJ5nywYD7nsj4JJtMGq7RjMGUdSWGeeNWbEIYFQa+3FkknY
goRC2YJLguJFKTy5GKu8u+xoT+SvNpXhlJ4hIX+pQLHsmLcL/ONVXCaY49TDazVP
DyrLgfG3Bl69bqb/Q2d4cjK84Uy6H2vrA7wHWywy4b6PE7O7NjQ7w81VW9zuZQhu
nyMwj1GPa3w956pAf+tq4D2ZGae2yZkqhAdd3ONLeIq49pKtPL2gsE2FJTZxPiQh
cTadRMnn/o6jZEUZFxq0cEZs+ZXgS2IE7A2Ghe3AnRBIYkcv0OH6EssqjEl91OgB
PcfDEiubnsFE/bCL86fQpnvroL7K0RN38x54GAnB/axNL7b4sXme1tm4js3Rnhya
LdgBacYVWUq8tNZ5FAqOceCoBDB74+qX3EcoZgYBKaVLzHgOd7AaZ8AkDDZiH8xo
4oda3b5SWrj1sgStv/4JwmuzTfjYxnKb/pNOFsog4IQBnAijXfOJWS44b7EimGYn
CBovFwNGIL6tq/JWTMer37+FVbUm5tTpuUESde0M8shUQ8SYq9AYgu3vP+Hvpz/s
BWa9pKafr7XCppyYUcK8D+46poshZ5KkBQytLhs16gYQE0koXEwbwSAxUCxw5+/3
KlW7LVBWBI64jWzvn4gGdPSiAaez9IDzjqZljbjs72VyTZHOLDnXuPSsQc0gF08L
xGrbIXItTyb9dI+2gou0WXQ5/R8a8oDtLUuoTL8jaS7RjmoZRbJ5c2bAl6uBnSGW
ox3kI3cXK7bAEI+nXgOEeQNPPtPv8AOAMm/2teFkMBmpEDVcixEj4O43b89+NIiU
fJ2E4esozYWpGCZ5n/J3XSNkLjvScnDs37etTAB3uutEVqEHd3Y+wCF0nvFIA9t5
rE6XLLXDOAbhpexuAzOsrQEjjEOm2BOPFH166EVFXwMO+anje7LBmPF/5IEBbPsQ
7ttN9hGzcuE8xuA5nMx0L5h4EqhUg7A0h/C9Er89JdKAVC7wxBAI+ASGpkrE8cdV
YbF2PUirHrUCddcMJM8aissN3e1RV2xpUGYmRxP4EtKbCjzwxxFfOrWol2GrzUEm
otkASI4V0+waOiSJF4w9gDXD0CS7FR2KE1KwXCND1dTR7OBixYWQ7UcRZqBE6q92
7iF2TNgUjNdRYV5b0inlN5tGDIbLlzIgBAykLdiIgcGOaFNdlVGuH9KvmHAittsp
NOSYQz+vryhbKkuaFdmPDq5V13FNCcSKmQbppKcmXJL52x1oP6uZN5KiNgg+lDGC
tBaPJ8CCspBj34AcJuw/l9ewpXqABh8Ts1gYSKQR5ZjzEimMusq3YIHsrU84R+MT
Cj5GD+az47AnOsibqNOTm1D/qeksiqgtOKdrMNJyA/a5+UYfriOnHpG6HJJpfo9F
GBUWxI8KwZ6/xlQoiTTC3h6Gai3694Gn1oC8Dr/XFdjzWzs9+7GDSbWEFmYyCMFx
gS35us5hxLpRgE3WiyM21H4R96R/tNnH8ddl2PlbqHL1NZwyg1g7jevMmqZ7pjiS
k8jaL6NOqrCq8BeoLW2ZCPA5SBI/BLXNH+92HoroG2hzvzwWbdtyybF5U7ZtbJBy
kLCRAkjEmP/fjnRla9aSGEUp+V/P3Q/xe8rlYuW1MjTxEeZVBKlRSE7ny2IF6zVz
DQ9M5gBK+tf13D7peALZIxZkyJwPfq8Li9Im4uvO1WN3UAdWrHVHRgsloL9XVYTs
pJTsL6JzJg526fazrFwafxxaVcuua5cevWTa5jUkrSaAQCokhHqumwJzGO9NJWnR
wLru6KTx/aBExzDxb9jQ8b/lbvk7uFyzkpl3FwTXp2P5wCt62pgT2pypZ5thLbG0
gC5LbdHUx4PzGm8A8WpOb+oQBsAjCdhr7SJkB+fw0plalx/unTbUQpK7c81WMIlo
8B2S2dFJ4/3Am+fRkUO6rqAEiYsCqCJpylYvPlQkc7sM2Z8h4Lubr8deRYDyYPFz
0PpLI5Vdm3UqXCop16TQ07hi7Yx4QMwEXWzZd94dQCaa059gxSMoFyRAzsmN3C9u
pe5TOafA9bBYBfYnXCE5Jnchy/UQ/BrDyBkHI6qpsJN3G1SwlTy+6k6Xmu5SBSvG
K+Tddf41FFPSIigLyth27Y8vQ8/MqJhtuSj1MUS08sGYlVc5P0MptcJmZTcGEtCt
JsI+O4Xl6cG34h9NQmVyzQqbzN04xtHTl2ncVWSpq63n8GVJNwCkpIdZRUklvMFn
qxRbuOssIKJpVgnJ+lyFg4f1i06dfIPXl1298XtOxUoJtY6fVnB2xglTA3THodvR
d62sV/CtoYH7pKaFP6cCA/brzGBv5NbW5rRYsoPSDYb2yz0qzv3RXRt5fEMR6Upi
xtjL84aHOyaB2p1oY2OF/NKZET6Phbd2WjL/DeLvlwCV1Gm6xSvLRWdLOtAHLKTx
8jV8v9PuGsCOL45F/btZ934oxN33Dtw+IGtML0IQ2dS8nFrGZB82zqybBeFF7QIq
6bG6eVDqHNL4WLSKntW6AsYMDTcX8Oh2c9RSRd7dkohWrmXsuNIb4E6XUdxZQW/S
pnAt7VNDkaihr9iMHLFx22q4ClIIGUHxtbDNNtcoqI2FTTYgZzJcuxnEsrnJMKK0
NKeQQEnh7sK0q2veTJuWb+m1T+3rl6MJZs6oFbeOfKCe8axXzU2JPshw4E+wXZCD
rfN1FhaKTtm9N9diWPeJ6rLkPw1PjtIaDSiJzUB+0CjOO+qkkuUlk2RzqJTYMP6a
VpxeoGrND9nctqoj2G7+1DP8D0AvQBZSg2TkhI+z+X8GM7KzfADaDFiF9t3gRJGk
a4JfHsL84S4RiHgW93bOPNcrQ3HnWLxrrwNmFXRCmOcFSmjLcrxxazzyOT4G7EzW
liG0penGnzeGfRjvc/0HT2wD5wzQasO+nUveB+Cd5KhcMqeruBJMg9x24eCTGAy6
u0ZNUsvrkbr9zQTc4CKvElRQJ0+nFRVnbElyaU4x9eI8ZyzJMwH2i9nzIpZI4enr
d+Gx3lVz3CKMlgrMe4rJyEGZXwcP7We/rRWqpcIoLdKBSNl+m/SSexfV6l98W55F
3f9Sb68zV9m+lDWE1Kw2pd9ygkh51VbigZ+KDsLAr8Wrr2f1in9VnkCq6Ig7ohMe
hMrAuB6DWXHyy5oK9qfbSljoo+HCrHkMkpixqqN5JrzzYq3PDYVoTkH0FcuYmi3Z
rAzkhtOLBoAAanXBpQ38xSIBgzlsTcIXOAtYE6dR6rDK+LuhGFhyVPDZcMmZS8my
LlU8kvLHKwdIEXGEOtlIOg5mcQG34XkCTGfBS9m2N/Uc5/H14mnpRmgkEZYHFcBv
jDVj5jVZRE0r12GZixEwdDv5g9hqrgQFS1C2b1TrIXh4ad1mfbSy9FibNljFGFpG
1rhE7fkw73jTZP1GTC25I7ArsApR4CIulrDhpp6CRejoSlKlsxv/cqwo1CQlmy24
YJYxn4D+fKr+d//u3pALWMdqelA/dA9ZnS+ReMy+ePJYfIpPm+bXctmAsvC6zrOP
1XfNj5OkfQjbf1M1RpepCwHP/MG7nVMzXx6yyin34hL5iojzkFhwzuW3rZHi6Avu
TOjtn1BCU+w6THUqp9jKOD/WHJVGr5s/kNF3BsjMgV5/tDLmImHx9mx3UtIWN06Z
f2uZuCPCIpSFpgetfoaKoaU/xOCwCTGuQZ8EfDQhsGy7/4YYWchzZPOmEzbPK2tD
5JcWSOrNdytd4o1aYkcos1Tld/aSbv65t2TARCI+N9ndpsHnzntMqb30dmZEqB12
Pt6fS898Gt3wY0dC4uTBmypH0sB6jFWlwAENpCNtEAETIe/VIDlCwEqJsn4+OLVr
f9Rqvs//fZ1FqAdZjHufqlv2Kd43aaBBjtyUWGnDK2+TM4mXhQk6zIrV9nnrchgl
Bj4CDf1jc7Om6VNASVBdbQBhn6EOS0t7erh5/9HqwHjjuQUUEEhPBV5SlmrYxZat
SfIRJPtmyVMvrN8U8K6QqigYNEoP2h/D+MDlve5lKFVCBAngRvhQAqYkcZmy5Pca
Go+rWOhbLnsu+d8M2QlPvXaq7ZL9miH7uKJdUe1KNWasryxVyTnqdX217YgSZ0XL
X1Mlv7xxFvBIMwYy5XmTG4LKrUCcyhdsVvkFfFfJZRa0iMO7XwPQvnGPcPQg6q3p
y65+7CxQDyvy7jbGLvT++BH1HaoxQLTgZqB9FOd197dxO0ERS5PSvTrIez/08giJ
XWsTTNCbaKoFd8dwXa5A77akrkZ+uiv9cHYny72PEbSwbcD6OViM2YOu1iNtVqeW
kBcQ1gD5nMYeEa9b4vmOAxIDyx0+la96vF2Dw7aZAt/vGihdwyBtd89oG/SWMhWw
5fyBCIXwNqEAITwYpqlirHroj2jWZjf0qgX1SvW3fnEuj59qdRVHXDCrWRFL7otn
xBuITaLeXz4vjGJrWceJedawlJsxcvBwButIJQxq1l6P847uQ5nurRXQdaiuiRgP
RNuswsPJbkIexJHBUcDJhjNRx+pSJw1AzX5m6yfdDSU78+xOuUT0eMp6TWtA8cH1
W7DubEsHGAqs5/SVg3PeEWrsE85FO3iLCdEld4+GkSznqvzz/13oe2DNrXbYsi6y
/pmdRgnNsduqciDKykVIfebMFOdQNIxGluvArdfKG4EH0hwLhGMcQa+cJXYwCFIF
+bK/VS6EeuogGpxAoa7W/qlDF8kprD+oeW3nLKzf5Cc5zbSgo5n+6VcgmvyJ73Y6
SFs6yBF2b1BIEYZp1l3EzvPNbK5vnod52Dw2spGXyhwJxPU31njVfVO4xuMtbEJa
4PkjtHOsWytpgCcfNCS7jgGuLgKrF+/SlYX0fMWqqZ80rOgRlSL8oYTm+dV0ihYi
Qefmeq7XWa9anV+sGHatm98PgG5uibHtCcRAQlS7tYjyVSKp0ikSqIhFw/RejkEQ
v3EYdY8nXy+zLYEyIL5U6/fylWJs4+pW31XasF5uBRI5+An3v822wEFWeOqOk2Ho
VNnzqPeMTE4UH+ZeXSDZhHt+F+QwzlF7DBThDCSuWAwqFkjpBe4UXgmtjieS3iha
ekDpyO4V8dQK42rh/a2s/KmgUOUBn4CJ8JhHMRZYpQgTFV0iHC5dRmESbeH6yfVK
XnZCTKQMi0fQKaBltofMtZQvUMarj8NuQ3kecI9usAYhl8jL0sk2jFrnV+7hnX4f
v+ZbMTQfznpTPtmc2D3oWmokrXMeEYyIZdBMrFpmL3eXUpgfMgwxT75HahL2+K/9
gK1bQZr0rqf5MBlXxp2L7r8KMUYSg9TmufhAkVsrt1QbMANbuo5/rnyq5BvBT7h+
2NTOBQ3kZa5Ha3X94/7UijMPoVdLqB+ukYCYVUGu2Vd5SrbQ16hsUN2w4QsrWpIp
Hihbl1n8dlk7uMA3SVdNQ9I+DEWAtS+SolTrS3lA44t7N326D+rPnvkYyiI9wvvN
xwbd/FZMyRWpFruaHUJvwCjA+Ap2dgtzV/pmornobysubcVg7/8iIvwp+Bav9ag3
/LE58DodtdqpfT43ruv881gibXHkI8Oxa2csKG1knwRMjzfp4rwSv3s+oiGFGco/
pl2ynSUlTih0HsN85VayPVB/uPKEPwuvtfexvgZGsxq3tfOgB2VCP2hslPgkADzz
ewS1jwIgt/XVidkANYYvc/kdnz2x2+YZw5Ly2YlWFZE90Pgq2T46gXo46dl/79li
nO69y8XiNbpE5l6jRLZaLFjnVSb2r81+0e5Ie6L0HajORX4Jbd6jdKGN/FqKDhX2
FyF0nUWgnyXGBLKB9jiXADV1TneWoN2zyF4vjDJ9nbtE/YMmBeeP+7Di2mjtI0yV
niowUb45R86eOFux1Ia8U5GYM8Fn2m5zwKpl7Nb0G0yCleqPDY4owf2xVSODfZ5K
AGojH3MpKKE3rAg8/B/I5prrYvHuGIxePsGmWwII7A2iq2BfxpJ/RIPl8G2ubOKI
38uqrGphLhzSzZN8Mek/k7sfblHGfcwLh33WRMvd1iKEBBBJkVh6zlC9HgwcJE06
1ffKV/3ttoiFR53tF7h7MIkVmgXiMm162jHuejJhFiMuf7ywROw8sQ5yIgiu7XCI
6UQDG3y/pA2zAzJkj3mUE/hhSL9hW1NFje4Fk6TFkufyoeWZdvyopxfies2LLRaj
ztLqtkgtl1O5SP+UGyRoUzQV7znUJ2hG9M3EUBKsGDJ1e6zNdj8Ryss2W9ps9Ydf
GJy4PtS2lXhyd4jjgQq3gtb3XfZJaW9tzAslaLymYveImu8CJUEZdsGLo/ix3ycs
h0v3bpi12Wt4CZxScj81rOlYqm/G18ZKsifs9eSFE6J+u2b8zAS4X3THgYIES7M8
OvCT7C76YNhSwLC0qoFkbGhANQTxPdCqLhz98TxMeOHJK5yU/GjnULVS2Ki1r1cs
vC3+Fi5obix7BIos1gFarMhr30Cxwlse/x3mrmVyJn2z402GUiM3032Rf7/3o7fR
4JUgMeD/DNqaBapWay8i3wrORbieffjH0a2NehGqJtfgzcQx6PClNa/Q9Bki8Yv/
WV4ivmGudTOQWoYNTfFrSbVomSyFHw6VEigTPCd9+l69HfRXrt1CYxVt9CbyDEb3
NRfhP7LxNy3hVlnZckFKc3ODLX0PKzoNKBIhB3d+D+McnzWInp9Lr5tFFQUqt9Og
oCJpa8it9bVw2FDiv3I0DOfH4ixj5a3R6WAr0Q+CsQo9FYKOCW09NLLlCA2BtvRB
5ePUJWQogz+JrQ/KSSgb1/yZILvclhyC+BMTo4DWj+AFYE07q7XJc1kCkw2MyyLv
WjNEltcqP7ipb9wCgpiP9siBil+Kb9ZujuVOzgjMoCWdENmDAXFlJIq8vWzDsb4H
G1EXh2Ggv7uDRAUm56KrySKjDn2UTMv4+jJjrF8v8efoAmkPb2kLbz8/C1P07T5u
lN6R61YlorxfHNuT8XWqwu8F3LoXTucn39aIjGm17uZgi+pmllaln6rkl4Zf62At
XS7MxVPiiJvBn8Lb2wyidz8HDMSH4HrIn/LUvS/hQ+iD3BgMGLP5QqvshHXMMvxr
cJDezgQ7cq8XlE3dON6/v3ZyPqOotnUbBUJjDFmR1umtGbauou3nnfUBOwHVganf
7wq4gpYlJM77dsMtVodWhnc+P9LpSVTEXWXNdtUw7PjT4Y9EVNUeLev3Xh33j11k
i0AzZveXlJeA+qCaRf9J2VHIdXntLp8s05rVSSWbxpDqlsqMoUOihFggmzeE4Dsi
z1r59Hv5wwO848F1iOxY5Pt0Of3LJadR7SA6gqtkYs2k6136u/W+nJkjcGycQee2
/DRuBVVuuOm9yj3n7SJwuBipToz9xLiFJvdyccNOv+73fCi5UMSjq2sECPAb56eP
bcwrv0ybDsRwCkBJa2k1LX54WrMYwL2N0/5/d9geqfIyCobzeb7hG2g8OdFqiYjX
iJOnKThnvcFlePRfLMVe+XhrjPFD8PO3akiIwiKaON7iTWCZ45TQaU1jPBVuYW/j
gvUoRyNYSI4fXV7a9jTJvFY5ENLZ2DQubAoUriok/newrMXJun9M318N45yuipaj
cQkGSuPnfHKPoh3OfcIw/LPgrygYFp31LOY3MiEfhdgOHWpndo5yFsKydvasXZ2D
S1poMi0Exiy4K5JenhQKGnOxnNIRAlF5fq0JkVKK4jb+mruI3z8FMR/vVqxuSgSY
jksEkmOLa8XP44eTZPViUCCuHbaCq92iNO7EIi4vH3aMxsM68l4X51V4KOq6Zoen
qgRQ80VVJVuTqz+0sMu1VlMjtjlI+agoNTcz/0e1yCR8IjgZkgxIHfxLgQmfvn4a
dnr7JFkcyI1IUUIORTN9D432J8XQB8ibxsQ7wLBqa1p5FeE2L9tmfqsAeL+0AXK6
O4/NppOfof4kkD+g4t+LkBib+DEJ+ZDnpLXQvwCZrabl9f/E2yfuZPYQEFeo0ZKk
cBdJ1LQaGrxbsqXyFKxE6OdyXpVR34lqDuXfEpaKucrpVVFiYckKutqUmW95VGhn
D1cClMRdFKDxriyxaymNBpsRTxGQatTPH4lR6FxlvLlCiSVOz7s1zyQc2aznQevB
LwAnlXRxUaE/Oha3IsfQR/ERHclKuW+xHB0HIopqSY56eIjSm2Y/45O+ksLY9m8G
7rm1XnnupN4ItQEfy1LNbIna0yFUwmU+kBwPSqeKVgZFrRMR9MmBxF8tsSAjfrGb
e35y3Oka0wLqs1dt3j7J09VVcdnus2Uw83hAjodK53ZNKWWLW0VJbWmWg5atLw5D
0c24BzMLJlNXVfk3RKLFGYQcf7LRA38m7zJBaQxBwosHrgxhETylmbFxZIxOX2zp
XYGmIV3xoykkeIXd5wOgM7M22w/+Cer3kJK+WZcC7JEvXDaOExcP4NbUFQG/737Q
C+F/woE9FidcH54355qXkHwnDvVyQH1x3/F3VIEBDrQv+Yj3hDsdeMNiVFwWdQuz
x+vQkZxNYtiH+YmNiVmivgYbSZtNf/1noqc57aFrPs4ATqJOU7aZAHLytOyMwstz
t0vcftzKxH28l5xWmxlCLpwtSttLYJ0bOk+KRTxPYnnch941QLYvZqyKGJqDjpYL
tkkSeGbP/94QbKRkUoc6uX3PAr/v52HUq2brkbzH0F4j5XQkumznu4EF0fIsDojM
3U5Tgb2tZMi7BqxsY5vPCa1d57k4gYil0lviLtKOT7sfPcqryv4l4vuLiTpiD+cj
lu3RQ9o3qhifgci0SpRxTAhXEVEKjuMleLNU9EYIlQDnBYyNjtkhNr0kk3J7V7+T
yWEKgl+ZV/h1nmqOkxlkfMl3AQRgdDxEc6PV3H/EZKVksyqLx0s/4+DWKtuj30+s
QZyIkDIIXkNKrnZ0j7vs8dS2pVbogdGMw3WbrAc/k2EaPvcdBd8/+QAp5xyze+34
fzltetEYMDMNcosp6PXjtxE0yeia2ntn2D28mxULp9y+suKSEIyzvyZBIzY6yyz3
4KLV5Jqf9rbP0zgEy+NjgM92xrxDCKNwnPXaHcJANC1jyMK1K6GzpY50TWnwLhWI
PI9ioDOpYOZVNHBC6l2OxqmNtVMA5ScHwEcQAAkj/E+JZrNrPDKQ2agm/Pbi8lUk
GP+Wc2h0IwVsiC30GogGGFblbObyVIiibRoSUulllwzlRww9edimZNBZsKrl8M2t
xRbwnHJb2WDzmYP94aDwXhQSMZaC+Jjh26/jJRZDh2/Er4+KwhUnSv2XEIoZpM1p
gY48ylCDnlhc5szGLeE+Uyh4ybtgXJQnqQF8OYO2TrkrCcw/S+jXaXTUFe1M0eCL
ftfVP74D+LBsqmi80LXdl7dz78O1F1FwBoD7trm82N5/W2T5DTunEVk/h4KIlgd2
4JAZ0icQWFdBihrSnIVkpAJ6Kx06iJOmDW1pRASk5jIjTUSZ6zqGSkhMjDwL7iwz
O/N6Sjn9wViFaMlHStg2iVPquLXL8fFeoqqFqRwv913tYhFpJyJs95Scbqo1QkVn
/58ZxevwP/zdQjTAM7hey0rI0DNQ5IvScOU485ikCxOhM7440Aghr0isVYP+mSrJ
kP0q3Czg+XDYwpPhxCUypu1xgZLhtjOYA8V0ZojQIH0HWoRynTVHOO9akOBBQx2q
E6yZWny/Ia9vnkW65Ko5x5n5JgHVbTj6lyZ/tZKkdQ+B8ayV3qr10cpQA5aD9kUK
I3+Nx4zFqimGfSoq4fICKDQw/fRgsr8G4Aq/V4CiHZo2dvAz17TsQeWsEZ7vrRWD
20SWRYS6RSAgr6573JkxG1QRFmSMbE4D1dJx6pzSa598wwnQzpKyUvEVQNKEKTlf
xpEK7mMsB0d8vF3aYP3C1rFCjmUvDl9I9hqGNlL7FryrFcTNLnWQBGYozPYcR/+d
25ttkB+WiexthnToCxj5rJyq6lKW3nodUWoxZGjU6OxrwHQ/dGxZL5yvGGutoF/s
mAzVDaoRBAr0cGFa8pVtVN3T5kfnoKCMR16V6bv/tKomxYwCGN68wfpxhJsrEwTJ
h6/eZfSw8LHURlLvAuNyN7JVUvAex52q3k7EoLA70BN22i/V1jdg3XxFMbe3yDyh
eL47JvMGG07jBAm+czRa1dQQHXg8eWMDoiPMnfPNJQalT2cjywXs50fFyYqukBuA
LXPfave9MRt7J1IQ7BrFBc8ct/B2/an0j2l1A6yXrcDcsuWIYE5nWjajY9EcMBcN
YjYmROAQuF1g0TJEOcDtJ06UiB/qIT9o1Oft/EKjkqDmkyWwXN23N9YUgR836Uu/
kZ6LhCL/2JsvqgZSS+iAixN7tzz/GU6sm9BCL7dkBcDDJaF29DArvVtbjPgyAmM1
CLSv0IZ7FwvONFg6Saz5CIqKzLQ4dgOKHIyIiTN8WBVTPxnJ7oO+sp7cTNsRaoMW
CJQRWlYbbobVfFq67abitbIk5CWBq6kvK3xcV1UeHR+mcJQr2zqWcoEj+8IoNYLR
lnyrDmygRjhd79+JeIaEKxRu7ebtTbyL7GYPVGme4haYF6O3muGTERyScr4xUtEF
TXEhtGcJEv1Aacj4WK+xHPOa9LaM8jzWsYTOgqvsgOe5Tm5g3feDSBGsdlOtiLV8
4HBgFGKx2VIxqHM8IpoGU71yR06nNaWT2AZJZkYlQ6eyWgt5AuQadjY9HXDtEZfd
Awnhjs7Az2A5x/1aMVtRjExV2yE5ge1toFvNKKDYPNNoW/13bmU3MwHb9IYJbTcz
sMPi4gv+GP4Hl3vP93/Z/72WJ2pMUCCB/WQhxLJ2hZqvohOv0WdW2CrfodncATI0
c7Ilsf7F4JbUc+ANQ3K/jIdbPOthMdGK58nt8L/ZcwL0avZj6CqfE6/NBdXLYwG6
ZV2WdFBuN0ZbvRzCkpfOxqJR0LI+vsE4lE6krv++KawTuegJInAPT7RuUkubAgJo
a8dEomSO8sAieP8aV5VPpCsenugRah/QM0wxiDxKf01Plc85cdt2Uwyh0KpjHYFg
KDqUy86nl5pt43+Wqrb453rM48aMJiD/ElLfPqUeoKZm2bH2BmurDF9NvPFAACil
Y7LncZfWE5umGhSuy1UuaEALc8iIbh8OQ+3pYVTuMaxbVm0tRRtyxe8ASvoH+gPp
bRx0mMLFILLrb9duFDYAzSjiGoZPzNsPEZASRrT1Serauf0/VyQwvNp/ofvO4Aga
8F00P1EnpkGTtx+QydTtQZjSD20OIaTGRncRdHelEdsZuvx2R9ADFpnocNiz+kBm
l1ELnwZWX6+PpO6A3C2ea0LCEVK3Qz/FhoR4Dc4mH7gNXHXFjCR1KwI4v35IEZey
tiF6ep7jb8vsBONTFbMJDruOvEOfSh9hyXir98R6F6P8zKBEq87HNMklrVQwBDcz
G/zMzxE9/g858vJ/MAUd3WvjgKVjRlYzViSMRA/y78Q01AUCGh/Ah4IiRqNHBOp4
aKJX5+OH8mzgEUV9Hd8Qua8wq/yHeqCzLNNSDMOh7TMIRRNR7ilUC/AHbPkoozr1
1qyRiQ2+B+8zczzHxM09dJlmXrvP4Q4ese0XXVV9ocj30edPcUsS67859tGlgSvd
MFrlnznxarmafyJA7EXZJPj05z7SRuhL1CluD+wzZt+rZ9BXHaIgDnw18vpUKET+
z5PTAQNBnxojpVqXc3SYmJWUZh+p5LxwXUTKJEql1wWu9OHWSpFOoO/qE6VrOJ5D
PoLQOpDDfkI/R6kGynXHHK+vxL7+5hfyyr9/HU4pBA0lx4pfPPr20bkjRqOrfxok
rQWafmkHrTuQe3kWldc8d+yPt5jEKhLf10WYFXJt8K2psUn7GJG4vJthW4l5+YNW
WYnKdRG7bT4GjO0D2TmuC2cE0ORmrH5lLoiGRgCl4BjgaZJwr3bjIDBhU9WPPaFf
Ky1ksraXxDW6JKxGEJoEWmKIkf/DanRmtQfv7PsVwHa4ya/+ynWib0ByUyjjFxV6
ncVvbbTqRw4+2uCd9skc7jSFTYp1yiFP+kgWLrSrTfpNfu9LQoDQRuc1OdBV9wib
RcFatndSH9zmsykcSE/q3njJiMYQ58pSr5lQxsSIYsPYScn5+ubNI5BkRFQuhCxH
vABBnpaNt5LndLGvjnYlLSuhX93KIt+1kva8Xb+dYXNVAGZ109FkZd8Vow9ZIzjk
6bOKZP6VAHdOlfTncMbCf3G9ROhp6ljZre+ye3CPiwCcq6jNxJhuDrmRFP8w/jqX
qEDLNvxHYyIdYiQA/lyrRVZmnlchx/EfwAxEj6/0mW49yLH9fXWBf+PlPwbYSLdX
1HSwPtmhjVBfmvKtemY7vSx0Rr/IiKNqN3mEKYIZ2/+DsIxCW3IQeTULjPo18Sny
zRZPFAXwCWN3Mbq6p6rkpFWv5Eag30Ax99wjLyUeuG/MgqAXeDaH01C4RG7D1mIQ
sotGj02TKPf0EWOo9iBfc4VdNBfVTipQPeKMN/l2bmTL4evmptmFtBoBIk4sGNfJ
TFqSKNZS3JAcDsYBFn7iahEj+0eUBDJTgCgNBucHsKpLzoky0zIYkXh0OjizdxSF
1LkR/L6XGiumVWczLFTSMa/nd4Cduk6ZUoGVdLO20VFxqAuBzeLw6GSWMY3MLC/7
4csd60cnDCEIGcpZK2m3WrfK49nM32WQiSbgMZQS9TmCDxO2EjTmAi+zKre2l6m7
OdRqpT1fjUvxNUNwfm+IBcwrThwd2tdzGA9J6oJ5MhSJDurRBjumvbEv5PKFxZVd
pIxJ5zcLrY5U4T96XPBZNYBqUO89S8ssT0S2KyhkrEGP3mXoldRY069F2blRDIfm
SqzqLJNGIpsKn1zB5BjH8RGsPINttsUlh8CfiF5eGfSy69birba7Vdv5liObsQ+N
OcsipIeeixqQUL2ohDJiK/OGQ9vxxJewEdXoa+MiN55ySBh4Kl63boMu8jEVUGD8
p3wWLEYTRINSpo1RBkP1Le4UG6wud6n3HSbSgmyOrEG1KMM5fXPqdljVutqh54jG
EtMPaNFdq0y34Ez/yTptwv7xZtX+Oklv6PLbPFmq0bg7exAKOtAH1uxkuzI8KIQ6
qZJwdCx1TsiwITuRsNtVRlmVdswasHRqSr0ieFemjkPSLMGavF4RAu+9hEb6ifHp
NrZKin1VjnYTIpzgeC9TatjwTn60jiLtyJUXQh83dHVI2DJZM44spaKapkYDp0N8
7ljtvyfVTe668Opej0qZSi+SFI14OFdKYAu1VXm+ICvdrwnQu4DM7dxvc/t2Sln7
aqy6xnQZ7SK/LIKe24dpvy2KtBnwVWiDUW9mvYK93MTraRd43Pnhe5AOa/vyYXFa
eDYXyv9xCtBWt5yHLpGI5CYZjMgnAHGR/DR8vijkhWnW6JUSIrCXvytCcvYSMY+s
100WmN4aoeWHSQWn2bCnuLPJCkI6kYfmJRyLkLWSGq0SV/0EnzxT6Vzzuu2E17QL
o2/s/lP3YH6YuhanHsiwt694UxE6+SgAo6vtyHKRhnW8UUV82BRmuC3NkS4v6wAV
HBt3F2hB/zSJIr/AsC/enbCa5obngBUeBqNSw6hq6rXlCjcvGxIj1sDQwqxDjIaP
1I9EKyf/fn2CPGE7MY6AHOuN1AxtLiqfVAY6I62quh9aPIitGNTK13cDMOISFmld
hY5Z7J42eJzmZvTLlDYBJ6vqY+nb0pPtXN6KRrWWZKOr1wjeG5xaOMn5K+CHUgy0
eN4e+4yEVVxg/ENiLx+w6yLEhJ2YfWbb2NCym7ZUNyISpySafSpl7FwncLyP5z+f
rSLes324Tcm9eNmJ/4esTihp9AU7Tq4GTjYG0RP/zYPX7908UWmMmhub97YBhVJt
Uk8z/4rFAvhBrO99Ll33Gkv96+YaM4+PB6N7qnoEwamsQKUdW+Qchmg4Nyk8pxP6
syaLNmQ+CsvKzAJ2X1xa/+UkJe00tDCRteyppDdWBZG8WtQuAHTl1t2uVqp61rtT
bh428QEDTQ8KP3YvrEQKO+CTbktD8KkSjwlb6ohSOKHq8wQnrbau7bXoN3Cssd2d
qV0qqRO+5rjCGbbEorteilB9huCBPu5HcmiPyTK2Ha08iy0hCi7TV3u+HDeR0TdY
FCrMAAPiIkG+Aiu2avACQ/q+FPps2GQDeF5/Qs+p5+x4nNGr128RNGfKSENQAV0d
nGbEFlh5XNaMroPMJVCg869rx0TuFEb+JiGhuN7M2Nn+wsuswwdG9KfKUtU9TX9I
9z0YzdmF6BY1pxxYVXvgsrv3yi6VzTX9UpEnaWp8ltPJI/68VUXfaCcOdt+17ouh
odQTuhFlqXNjI0LZ6EiX9NRDdnU3foLAcehS/APVI2Z5/9eXcFkyQzAUtFAREQLu
h/YQOmqkHD2MAuDyJdZHV2dfqcYhtUKMtmkLeBsomhR2k6Z9atAywo7NazT6xhLj
wzjt8Q6A8rzbGOdzj5yEndNF1CzVWP6M0E+ZMER9xuz68hUJub87vbqyBQGoo5Ys
7pJWXSnr3hRXPrPSihh8kSJ7fND635l0929lvJqPJexoQ5DBe5yIROS07jljsyUK
ndczdYeTivV65K5CezHtZ5q/2fpsWs4yigAH/XDqhWy8Q2qAPu4gelfTFvaKCcdE
Ubq7GlbS9GpwSmKt4FYqEArN70eJstn+hLG1LwaLsZ5Mfeqr3BCavPRzS+Sz6/Gg
Jg2AbrH/Vg4uMnJu0lINTCVP8XUXU50g+P+vM2HDhBY2zDFuXeDGiFPzyZxIZKTW
XrHkS4HKTAoQ6bHr7USZU0xPKeX5RH7rIDDVL0Y363RudN/FEoSXCVK6DPeyHSSW
Beb4EmdUEL/C3h4LEZdpkT01FiLLE0UwJLMUB6JVwgOFQP47+wakJ4+MAfXzvNjy
JDya6okng/ktKgfQh61/Aztm7ODA81i9ICqdNi7pcY4ahBrGl64YW20uK4l+62aX
WPAHXKWDWWYeBQkptlgqFzJvjds6HodtTXQje25ExCV36L2VZYbkOmKn+oMTXuvH
7MortHGPwGSLs8teCPHJZeBk7NXtts4LQu+wdCRCduPCxQkfyT8enmFaZyCdF4oR
/1XLpgo4R+HoZRh1uaUkA6y5FNyWBkSzPKWaHZbyOc8LXAt1Zspp6EntdIp1YPvu
AqYsYOQMA1Y7gnMfQU81N7bUaHcXlsjipq8b8EYH2o7TM0RL8xCe41ar4YiRltSW
6g+5CC6vS7DGcc/1/ClvLfpMXhDAQtCtS+S/ySp7K140SbPvBnRzlIImdpDo1dvj
z0+JGxaWJD4qhNF2qfnaXGvcE1hBm8JMQSvne59pLxuoq7fVgsj2nyX7NYUm6bfy
Mi3nq8GiwSaW1hWXbAOauEqAxcNFJZE/tpNVQbN0lXkVCj1iaIKpUNF3ezjs3qAP
Q+NDB+4szhS/lawlb3zksfONxjcPsedgMP9Vf7Ahp+9+g4pPATAlIojjFxD6A2Gi
9LFZ7MCRyJC/3nJHLJZp6jbThdVTPlKOrQIU6CQ5iuPCw5ne9r3YlcrZ1CpQS5Tf
d94F+WRJVY51Fp6MaDNbmHnpD1R5Iu2n+hryE+QEaEKMMQ1wqYYui7oH3u+FH+GZ
FUA5cv9MUnvIJPHelbpTg4ZKUOSeoiRpDylYqHocQi+l0tvEMMAsY4g3XO0+EOUY
MEIDsLALxLAvRQc8eBbWw8zH6D12aNnvs2f2gGkx+oQJrnF7PMI+uSbDtUL1UCiP
Zi4it1Q5GAEPWJugLgqw+uRM44Li3iia4C9A1JNzKB8hp+NzXcKAXdeMWqxX2mZI
82ofVzR5lFvAlQYtWHG/iKSaeU1zCnaP4PYOi7AMtNZUlPf56Z/8s816At7/3IZo
98DbQV9o7eVyPJr0boLPHveBde2i43uiQblTUVQVybGhzi18U37mgYTkEn1G6dsm
VDMfk1epfRwiBbvjg0AntVra+pXQd+aRBk2Ou0wXW9s6cNRzzOExqZ4A5QKO16kh
ogRRE/1DRKxIVLty7J7+VdcPyb7tDM4bX51HOlOcYlAFPI3kSs+ph9tMWj0WvEgK
agTgPRDT8T8h1+HuZkfNc+7BAn4dkLG6jcMHHDVYXVcopeljZcr9gIdjiYOIPQnC
GYK+zxdPkRko6KtNd9BQRzYvxKmWlaPjEsN9L3CPrYeWq/bvK5KHMJXUzBR2E8vI
9aC/LIIPhArTBXvSxoAdu1E7g41kqu3zIMjBNQp/TE+KaFFp/hau46U+A05fH1sO
4isZ5Oss15GzwS+bM062mkywPsB2g64NuSChhTAzqhsn9VDIIcXhxzVwQ9LjOMBV
3NXnwj96hNIDCXTVqDckuIUgHUPXa+2ZpOqs4hSijbLIaMtuHKLyjoGdZXheUvFj
hhN0ow5JvMlnMB09E9rg6BDp1gP6TGnJgKVLhpsEKGnIvslnXkS6lQ1AkV1BmJUS
gHXfS/zIDFMCVk3y3ys3nXC+6hgLgrO4HD/IsKuzOLD1OzU5WrN5OPnyFR7xyKFJ
wDNlu5QUwICWJw2R4OVpS+r5pGBsvc8WxGU4mXASLBpb57VuC9CcND4O02WLRGME
9tSCvNB25QH2s5wAg+3d5IzHvU2zYQ3lNFkd22X23UJRR6dyuSnxq2pCehXIHG/d
/ryxoLm4SZnU46tCh8FstXPiH7WE2N5GgYU5NaLlCDWzl2nPygz2+ANZnHFH/YQP
CKuMeNdydS5/pSDvGK7CxJAYaIRnSUUoAkaXynjerZW7hlqkCFA0SuAWmtpPmZ6l
fMsIedqAhr2XTEBz2USI/uBOZnpDYDJJO7vROfelkVb6Tp6r2N444mwTHVqP7TWg
8JJHMYgjvTk6lKE5w62sRsjl0nkTU/Db8r9dBvfW6gxhMAFLdiJ7/iGjowW5l5se
Ju1heSk6IBpmJm9v1QcX+zQgJo4kLA/S+sXMH4fejzAfqQtUu41DYby/K1j87FcU
HKffj/eVTSt+VYBDWAL3HLF/+CQFRTnM+LavX0o5Sy9Uw+4pDoejJA7NhvQSt8HM
WpQJlMCyhw7SOn0Uqb+kHO77H6ni894zw01iKHkX7glIFXxeCQoXe844hQVlLYyG
Tje3aVzt9EJnZ9p0OctU4vtbSr3/7zbOI9zezpvK2ZtpffbZY1eJaPbfH5jFL1rL
J8VQ3AI6jAczS/E0eCIAgAgjWlbyvFX4UT0/l1y+lH381T7cv5ozxkMg8f4rkXx9
9FDrk2zCllYcLUem3qNqmQwEybaYvDjex+646n+/F9i1Y8igcfT7MCC/nW+EkHqX
QaV86hTrphnvoxKSeTHinAI1MjXdTvbm+h3gxp27raxJS+uPUESlnmSe7hi4gJC1
llhoVDlzx2LOIJQ/Bh0iUrZoDBveCFAmjc0yinH/wjT3ReSvQ16r9/tfazIv6eUy
69NOniCEkwPbgIlRJfr55SCWvjW/Y89hAJ0Q2PqXH3oqdIUzFtCpWOr66EESxQzP
QyhXO8oyWnRKha1pgNO3FCux6p2BnPXyRiZ6NWrCwAo/d0WyNhL5ewrPoEywwXuo
OWP2TF8LWj7AxqygXFMhFgvzmPeGnvhh0gFOOMY8HhvbqxOlgTlzkoBvF5j0xDaa
VknGivCnlRwNDd73IMGWQm275sDTmPuApEQjy78VZCeoynClSSverysrS5KWxjJH
MDEmX+U1MMgBkt8NDdqqBqsX3KnjovX9ktKnVMNCJ/A/7oA84C7OkuoX0yLXFMV6
lH4m95JHVk60zBqalkeszDsVQNeXVKXSECMG5mMqDcA6m18BtFcwlJnh7n51ymxD
H98DHCQcvRlnchDOAGzmcMyuNxq4twCjG33g7kkF+6D4MaSiUBMdyI2oIuPYuFxu
5AW4yUsToFWUDqe3YEh5Hl0MPQ2szlTh1Kr59LcPLw2ApiSTl7HVNvAhhvqdtXbl
Np1OU4PbOgFb1+9WBrRWD88Wew038QjzaTKN2HPp4o5EbNzMChRRcBrR48NcwgcI
n4FZY9pKdec7p/L9/kY4jJHuJT9WXelTeSoEG/7jN4ftW+8MQbfGwrswldNxUyZl
qwez1Pl5tOMDmR01YTPjTEMlauwFp8OfcRB67vBBPAwIUxr5k45WTB2U8BxG+PhI
N20IgLp9JC5qCVto885XR5y2PW1kt1H1w7G1hrJtYpc0I7nTG4XT57xDEgIHmueC
3olR3Z0PD60y0Jk93PSHcQAUCJ5viDUByRW/oLSSrx+NEF7qQyH23GoIIxj+8KXp
1Jotp5YWocgHWIYz3Cov9kUmhGXywUQa1NCkGhSYY9knatxtF05Cwhlu+INHOLMk
lmsXrZDj6t7JcGq4CIUf93geWFlbo547uspV7gZl52jVIpiYD4TJZHB0jUWt9rLb
91hACz8ToIF08LUa2EZnF9FboTiiSdl7esGwP4Y7nQKrvYlXVE1tycHPBASkGMMa
UavL+s9JiZZXMTXS+mEzm9oW9thAns22WBgHwKsptl55eta9Jg/0Sz4AU6zh8jem
j8RutognfN8OfUnrMtMilE7WyatWzbS15CDWDsZ/EldRgpZl7Iz/vseeacR8phcP
1/jdXUkoNHgtJMS2++I4o6k7kzoKTTf5xZXviJLFZlOU79BcIhnIA7DkjElugqBT
Xe/J5vIfTDHIljF9Yj64iEMXD/otRSF0M8vDl9WX2vJ9TMqcRQcycE3sxOgFlYfW
1XCoDWad+326OwUARLLaJJPRKewwLtOfDnTbToiIx+fLSrwC4k9HfG5kW/OqFFFy
du0NmAaFpYky3SLDkm/fWoojtw1hsDVM2Kdc7E1QcPZZLzLPotoZb6pj1QvG24j2
N7WTXimxzIGskwpmIaGRwOmZS4t6jQzF8BpLe3TlnJPQp2yUJBo+xEshAMvrLdjN
y/YZWGuN4zHSMe912avKUPtjHGN1kT4lz4Buk+KOMWdhN9WTMZfhc8Y3x48HmRhd
LQDsMxs2fktF4EjAmPY871jl+Ojoa4Do9d2yeCR+XbddCYisRD9Z9WZfl/n0Of34
ApFkvhAOqC1YIjeQqBu0Yqgr3rvEFpneG90Xm9kE6fPMm5muSALXG2avFK1rzlwY
7YLz0rDaOd5e0hx8yqIKpbx+Ykenn5cJpTNHuWqHbWiukl+NhK44lTi3J84OgPUP
EBB6EAiCtmAXERpdj2MyWfmJbxA7LD/Lfw0lSTfGpGaWBTQONL3q9a4sHPeo6lM+
NWODuF/IdG+IRpj9EyXCiJ3oRQYNvjzxEKYj0+/3ct8TbIhgs7IsjE1niFwaD3WN
u3F0u7NfOamqit24CtXU/6U491lvYIf6OwcrpuKMkgBvSFOcDIaeXnpC/qSyUYsk
33IiRsqNTGVMyoy2rPWKkFcF8cXGIsQi87QtO670aYjRde90FpMc+4/Xc2Op8bTz
2qhXajrRto1o92UZ18cq6i4CqFxkAD8LkjXL9uvIOcmYgzdL8Nw+kVsLRCs8lWpV
inQVKkBeZwH8zpc64w476ux9bDDIpkqmMny3ByVZU9JZogm8ufMGIt/+XdX0Jchc
u003deuafhR3GUV0EphZwQnDRM7EHQHUBzbwhysBqOtLl8M/JNFTChS13HhlISmc
ZvG/nSBctiIrT/fHFnf+NH/qifLkBWyoN4EliR4qNnxtOpJyidgX14CQuxDLaAQ2
LzbQ0PiMNKxbTyCbBrp5FRcLmQo8uTBS85XhdA1gsIq1NZYUlRGzbMtzFhBf3uMv
I8TMTFEQ9v1Q4LNVhZNFqQbfmpYYb4VgbTVzg50YlRhI4rM5EszkNUWv0d3Nz5Yf
IHid9JK/b2RppQqwMXxWM+B0Q5Nf+EuAJwQXodkwCcwm76kU+htXVHz59ZvObOAz
IsvOhHYit7w/5mCFpC5CG3ryTPPBS5SbArQDcPR32rmrzkf+OF8v2HfTM8doMfC4
2rIlc2+Azc+pF/uAlkkatsID4oZO8RzNLW4uwA3fEDJC84hIuwxkgHCIhs3ylfTr
3OClaEQMlE50LoscpClvOLGlaEV5Ld7c4mC9EmSmLVT9mfW8702sHLXJrBrXNLWI
VVAqlPoK5qLgQa+Eno6rPHw/4ulahGZXH4e8p+YRZwC1W/kFk5nw1X24oDcjLTEt
Ob4T0tmM2ALhUavB0Ytp7z1RbyyS12AkHbpISB5Tp4U3fajrr/QZr0ZyVbSt6qOt
m5KMatRBbwC2GQbJeFdgoBD9CW/mT3jbUVqxlOrs40N+MIZT4OdVmcf4UIkprV7p
fzvSara5jlYKc0MrOzZUAy2ktLip9awvGmZrbZ6bdZS5zddnctbJpuOl7StDS5Jo
gQkgrm3EsODqjxquqC9+ENbA1vG+sFvlHGaURv4QeR4Qg2/5lJp7syjgeflo2Onm
96cdQE5pxXXBnKqIKRApRQ4TrvgnNY+0EUmtjyRO7E5ZTavjx9TlOS9NqOwiuODe
JJ7pBF6/Wr9Q+Ft7+3/gMu6prHn8LIUhfUIaZ7CDoHqRB28rNZE9Ks5zJgekY6os
ov0VCkwrHYSUWnWqdbGmAXnQAQ/913mdkrN1txfIBEYcTlbEEUX7l7Jw54dOSLgY
VOa4ygJ90ySYWYA02C2YfBTJVZ/SCzuCks3tLMhD1VIQiJZcbEz0/LGNJeJdNrcZ
o7ivQGIui3tkrKbfZKakadnAidUlyYhWWSqcSw/1EDi3YgVJ0moEV+YXaC2fx9IB
J4/MqCSFXjWz0ZguvvhxWlWT8nC/RJE6wDIm3A+jHddVccgtscwIqg5I83KVHrN0
WJdRCh7y1m04vOR1az11/wA7hQx0OiZ0NLnXvsI+VNlraHIJe7nAGl/pMvOshZ3S
x3DjdRHJZjdGPO68l9F+x88utPnYxqz/IglNkGRY+E6ZoZ7mteOl9vK7wpDQBDDt
8JrcLRxejHxluiIosd2+hThi7Ge5G2KjkKec886J/jIq1O7L5jIqn6iu94vjnkKS
PD5bQ/9dTGz4pUyN9ODscQA831NA2f2yYqiF3KJtUwXsZL84r8NocWErmjfAsYIc
bxZpsDJSjHJRE5ViCd8T+j3hnGAYk32XTF3Ux7gEy7FTqDPNZQuupTrLkp3zQprJ
xRM1PLriiLIy07Qapa4t1rIE9/rxZ4w/+Qheu8NxP0IVepUZrlaf9ssH+qWVh420
Vy5OcbUmIVamSATBUlNILhHrf2BlsN5EIe1pkLSa4gSy0EdcMgbJeBfoSH/Zcc3H
KmAq7YUXlMlb/xMAsxy6CEzaD3EpZIEKycFofXDKqhpLySBUWgYqsKl2wkvBy8up
S8NL40zB5u7KrNMe77nghkXthzzKT2+YSOzDs1Q5MOYRA8hSK+YGZw0E5gIW6Ykc
dpt8jVSwaHjG4iqx8LE7a45V8cPIGGZgqMdgqnK3hHKdy0GAmLWtzKz9dgO+2Txo
10vSOehFcbxlxr4eyxcF+TIRAKKp/nS2idhz0T/gbxpoOcKhwN9wH3tr2SlLUgD6
xq68/nu+pLLmy0a68yVCO1of+agyrOPxoVElSZOmOr4vJ4VOFuZE2zr1QCnw9LzD
EOHv+VZk8nxH/XUjwqNdAGKnr5u1T4GREsZqv7dP1/XgBpSTkBQQbOSaTAazUCqY
uEwPIBplaPUAejQYuYb/TpjhRHnPGoKMZljEKxBZ5szDJVchHh0/qs4g46Xo282T
K6+WTiBiqxAZ+OnP2xHa/8bSKVofTmAtS3XQTy+fF3Vim+k4l5kcWE3vBSNkbXoO
7S0zy8YTBC6cTSdRYLP6ipQ90YXSF9+g84fRZ34kA8HyGF2zyM6BKasUVaPmJCCR
dlS4mudTlHVdYvL99an9EdpXHS1vQfsZjRuGlB1WmxZu0Aw48H13kse2xr8EVX8K
RiFDRtv48K1Pfp0/IxX9h3FXNqDhW0R0jUwQsMRkxNN/g4iYVOV1w8bfikteq6X/
qaA6sPIP7LZRLgqcjGv8z0RTJnL9ES1v/gHEM0kLu5IL9OrYU34p0G+se44MKCpE
XJ9FPC7yosT54nhF6fhdUuxLNgrflRinPs39Bik1nPK+lZ+Tvfrju1nBr9pHeRPX
CUJYhqcZU1FrjNNneRGC47LKmY4W2l5/rdCGDsJpj7YKFK27ElLQjsf0cUKRGc4i
Koaa/vW6BaDpPgC9YeFdFjtdxlXVn/iJwldBPTrL9TKTvtOoY4CbWcH2QETi69vE
5VT6ZX7zORFCUo5KIzwjNZIEyp1x1zvztX+nSaMDI7eILqr89FaeFqeeLeAND+zk
1dx85luAUYf4VHV6rP51bXCIiqR6QNot51/zvCCEL+W02onAa5z+HMJfzma+2tHr
t7hQzkx2G1dO9kZYG/5D3F0zG7bAS20QrGheFaIpkP6YVa38Lkf4ZD2yr1EFHo/D
wY8MrDxalmEa4GbLnRnXpdD/SqgfPStF4I/c8rljT5ezA3NjjkzX/MYWgt2yBx8z
BPtXohJyKgKVVnUZ7xLKDLmDm8m5UFjQr9M0zdoCSNF3sWphp6w343CRG/ScRIQe
nFgDplODFz0DU00f8ZAVD/VPMgqhfANKGX9ukTxqUfgGITjVDWMBEUOQhZ+v7iNR
avnn8owX3fhj6DXd6OTk1krsyOSDMlgUUYMAmuRnfMAke76WCzpljxwdXkMfC/Ha
letousnePpppRvnEIEEvzAf4cQEmG8lHEwlgneNPbmBywZyLgwVF+qR3aK/W/Z02
EKJ1nsu9dtz3zaIIFFcNG1bTIegGxrpP9bF+NVzE3yO21D7o0xJfvOXTYR1WtrUL
L8BMjGF4foxLKxH1tPmsygPh4Z1Lu2ZzvhvNSsyzCcCJEGW633qXZbmqYJVf+9mw
/4HGN+eEQXnITSrjOrA9K9w8A89eKsfQdWpc+O8hg17A3Bt91xcuWNM45WnHUpZK
aq6kN5SXyVFfy7y5oLRGwsfGKCqcljq2o4/3syB0nLyyTPFfj66W42TGeeforiVJ
bgGc1ZySRrsfkMObd0W5SMm0kDTPopB/9XgunwuNvhrjIo+CtlkiufkUvZ/jMEwW
TPNGmfNjalQeKOCuOIHAQZ85GINKbScG0W2h4OIRIn0DYfre+IKhd92fGsgYORB4
6PYdkWclqu0GyBf2d+i423+TZwxTB2cde7qNjhAm3XvhjcUe2fL/VZyMmKPG0fn/
wxd7nzY5jRNAkHLMoSQg/JU+GpRw8mtfOOP2o5j307vPKxy6+G01UlvDEpb6/8ak
2OfLX6/EywUoBMVA5ZiU38M1hOxDrztERGN6vg3ZAiSXhOezcLMlfKMDyJXtDukr
B2zq4OLEdV4hriQDhrMn4702p1fKmCzUCj94sdkPMxCvOmd7inZNQ/7+b23ggAVj
iMyPG+XTlJAh0LMRv0cKw/mm32OOt0cxtoUP+0c+BfvpB4oA8m8ufX93Fv6RuhE3
ObMVKt2VBDvnB+E1VHI9AyvjCcmRDuZvfiqUej8zNVuAulqItRznVzI6qc5Vmh04
dO2x4BLbBaUqLHZwSaD9bIC0NCVp/Ltn86LlOrPKaPRxS7WZtn9s1+RESTbkHz2w
g4ZCH4I2gwsWfEGI6BytaTLdfQTXKIrvBjCMvdyVPJ/1R7SxLp5xMF3NtLucikXP
TqL9Dz0I0Dc0NTQtNooRwNsNcV6xZTsIjnIPmIn1uri48UqhLjWaHJ+X8cdz7Pe5
eupSm7YhQrTfVILej6JxRub3QtHcvUSVfZ1dih1jiWqkgY91iIufIBzh5c0qVrpC
l5zKVxBreRDGKxUZK0o+C/XmBxwo0Cwf1yzmeHoOzC5Q54V5LQcmbiZE4wu6L1Ch
9gMCko5V4fcHZ7srq8r0eShQOOcuDJEAP+RR7B3OcgKNGv3XzfTm1ekNtQ3aEG0b
8xv+OYh9Xdsu5S/+jVDSPb8UvoODnHQ3BWLCpjODgf1dI+2M1EC8hlFC6yK7bUtx
iKeQYqRm/r1vPvROY90pVRDuP60PZXUadKJ3xzzwh6ETK/33hUpnWrv8Jc9r664O
q1b1YHI2s86zFMnvY7PufEApDwGLhpAut3/ZXzgwjj4AHGB0+tLBTd3OXL7lSJk9
XUftVLEe7+9I61I9V2516AfpFuB0lNQXDxxsAJ995OLLCunH3mAmJtRd9xfAoovP
wkijcuWtIKhuK4VnGkw2OS5XDwkcFqKXEBoAU5AsrVggV9Jtsbyfe6T0U61D5Bn6
tqJujocemlj0Vn0kabB6ZCR+rzjzjEvHd0ZFf3p3QYSEfK6CQqOgswNmhA2XNViQ
930yZTqrl0XIWBxREyh7VeJ94Q28nv2ATpVgY5YJR+Kp9vwwmMh3NtZdCAW64cu5
s81PtrA0/ilgn+EIFDsynenfV//2MEAqPLUnC3rNNDDtV12AgDfCkq2RhHGGj0Vy
OxkwEJaoOkgpeTzh8553JD6RB9qWcQaxOvRGa2TA743/SNZcUGiTbAWSFAd7vszl
kiIMHbn+Hpk9E3Zpodsv6ZYh8o3zepqJ48F8tQdwI+wKQgbLwWL0LYpHQ6jhnbgB
rnqZIJ6HUybB06eGMAGFSSOhxb8moaBf7apW1gg0l6GoD3PQfYPTTVfEyM8BI30L
vG6+x+3LoYygrbiWxEIjK2hcLU85g9UNlj9Js0KSUQyXnAtPquhpBKmLKh13WHTJ
oU+GAgySqyL/r1v1occXKC2s/IMN665XsgFLjBePKMkBvLZRUTeLVlM3CXTJemm/
BQCJ1FeFP6T6SzVyvON/d6Z8sddj9lpxbPr96H3ahYs/A6NhnVRkbogODLUZ6a76
VKd6i9LFQGC/Ht2VHiyRK2YtXDLYZgJjHAdpj3iNqHajHyMUeo76jhxAd7SIpis0
9IQmessbhliysPQ4pM918V+LKTqxS3JsGx+iCfl2/LdSVARHOFb+SbR5m5GXBYZC
u2ROzjVwrlx9zZBZPWXCXMUEDRUz5gZppTqWx9buCivu32havWunZRuMjwaK1i9/
0zzBbYbcAv3zwsmIzOwYjNwzloxJt+z5sQOAVRXk7J3aJcO6ALMKGKVgtpWrlK2V
FQfjK4Ys9zJhV6rnv4rv3D1ScmDQUY+TnrkEbu9NM94g1AhK5ZN6g7J3q+Spvuv3
alU0zjkf0TrdUUJ1uMtQMpWBDQD6n1Egv+BYlf99LP/mcnqquOYfFbD50oHmRBh/
TLOlwuvPDQObamCi5G+lSwOghHZuzZEbnVR3LUfe2qjCi7JAfN2647IsTHBs4Zta
xKBav5xr+GqHR+ohjG8siaL0fPf95d3sjRvjHbZ8HSXANqib3VRThlIscx2cXXSV
r4mkD+W0JmApeBtixheaML6Hhn2EU0icm7SQkLmhHEtLtkgKKeFxy+bYZnX10vUs
38jowbgpaQee9CHAU2QurXgidj8ACMrGD8Q6jlQKSBWR8ZCIouyPLXRBpG2HWoRt
fn8Ad5MSUoYp4zJxCUyO3Q86r2ObF1N3lMnV0e2T8REd0FBhnJT/3xle+J0qwvkW
WxiiU366e7wjKfRO+KJF0H9vmzagR5Urm58GDXIFl+/vijYvCIxZE9VVujOA5IQQ
ftg+alrojXtnBqoRhbRtQqSl0y9wVhb95QiRBAT66wgoaaFhBBxskEZ5G/6QVeaJ
CMyU83/gVxIPTDxXXH4HNLRnQAjlhLCN6SexKcWz/8a9oEV7QHRYRi5g+YpBE6mG
EtfsIMdsFfujaYxvWdCwGLTrFk2F5HCuo7YRYJZk4poEXu5Q4QJIDCOT+H8jU+gI
Ax2so/9MathIcw8U3DfxLXy8zs4iUBcfl1cfJZO8LA447RttNqHOh1U9DRswqJRi
mhQk1sRPvsrUDwE+rjxrQjmsKYN/5ZfZRqeiVMdpwTUdaV68CHB9c9vIa+ru7jJ2
8Yl33pOk6S11CyhiISbofMEt28pn7ONP7Q+yloJcIj3VegheaUbhkHkCgetTZAWY
6nsjqxQqczh3ui0asT6bxG6T1ciRvjS5rrnkJGuHLXmTIfS3An4ay0SjvjmHwcAO
vmuDbDT2QemYvU9VV4gfwib5q5BhEMA2sIUsfQlqL2jubE2tkjb+OSrX+wnRpmLA
pktQ1r42Zs9XB/JI19xAPF7tNTRLeqEif7N24+YBseCoeq4M5/xn0kavsHVmFTPY
Q5ejK0YTF2gQ8RS2YsqM4Z9aLZHa7fFzRw5M9lKFdjIQ9mkBV8Xw+pLbiTejGbj1
dGCcL813H7vq2VYRkUNJ1ckLaY3EcxI15DeiN0s7YmnvvUa9Xi/fx3UcFoBNQFz0
yrMpUMLLCXtyyoR1obERAaCfGDYGRYJJc2UWrykVEMM7HB4508MeGvNkuYDp8GuR
E/355tiiqcK8gZmxdKEdq+BYmBtnijk1ZEDkMNK3wMGj1WViy7J8sdntz8M4FgBa
n1LR9G56TO/mUw07wtDR3tuS4x2gkRei+ZH5DkK0YdBU8Am/XNsLAU1Jy8qo2vNr
ucOaYLVVk+CFGx+0pqeTKFEK7Smm6u7NTuEsG4gh0BK2iSyDqSZK+EvZFgrqcy+X
UbCMO+2KZXCKi8Plfu83xG/dgkvtKPfEgKuR7evICrykUrqas1GDb4E+mDHobZGd
QH1CQinqYIUHRBlstIUHqSlWC3R/lKJroH0VFJwnkCwXysoKdv8nFTEnIXXgyCXU
3kyVlZw6Eu7xc4/3BaAbAPRBN/WEKB285fwJtbfH9RHsmYuogSicB898NfCZ6lya
hXZTmGBtHpwwv6mIR9sjhPF5PSUeFEQsPS3eYf3MzSUafWnHAOsyMYWq2wGThZZv
BYiR1v1C2Qg3JyZvDnY3aW7nBiPrBeotBWiXnmJzzFyyO14JgTDndQPNvvm5fqMA
AlPJ3aElioFsk8/QFSnZqLXkxqhQ/PMqDmFiN6NMgWUW5vKe+C66VIp49lOpp7bC
7Xfznn/3WcChYTa79/aZDSS7oy1jPnDVIyuQJ6aBSzaQO72AWdx0Mr+AdU5NZO6Z
qxzTyagx75EnYeCzSGBnM/Sj9sMeFigWeOtwaLQi01evPxhVVHjRkICQ1MP1Fol5
YwCYb/I7ErE07qG+LOlNCw9FscGghJdf89ncRwWQVG3B+iWhu1bt76k0DB0poxGj
SNkN3h4hjjH5HSY0qa7WT30+x25AUcf/D9OPKaimrgZJafWQbDY8ERG33+m/DfoD
n+m9HYAMMRQyi7uvQkLTusr4J3gK8hcJKTd3ZlXzKXYnetWzBXZff5irkUD28X+t
vCIzLXso2VySsnwjC035sGvxAaXVvKTUR+nh3qr3cBg4XXxNKD0YjnK4vcaeYVVF
F2aK9QjsmE21PqDKMhh/Bd9lfq2jYjcvSSWDnST18jbBemjFf5AvNRTpvrsuu2nz
BNr+HbuPuXqLol4uBFLTugThrw5Emc8j9keE04Fzh3FrsFjj6QkZ/CQeRCMOqo/W
10muiZN5KFfEFh2qMVcqq8WAGbZOVUngrzy7bRfrKQxvqaMXeztZBPMX9Q+zZAZf
/1VdamwL/xW1WPMXjoiIVlJRQgRdhxNWjdvZVTmjA6pEZC/KpDqLYkkgro4EhLLL
dsVRH/CT1VfRvO4v0rZuDq2BscGp+LHLpRtkWnT/x2y0cDJ/qmrNb2XOTRC+dfjR
90aGj/jklp3ikdOcoTqTyuIiKuS5RMVAQNZx4W0fk9pM6RrHjFe++9eGCPB1mivj
dCRZy6simvOeYfN5gQ+Pu/Z760PAPO3JL8CSJUbAwIA7BmE2/PQAE17m2+okn6ZD
2Xff3fDixMOufDn81Yd6k1r/Qlpt8iz0B2FaDDi5Is1E8DsBcNToOM5F9iPRnGVj
A9msTGS4zgWXBd8mhioAAPeTUHGj89jLAMb+FCILT6fIRalTKtxQSqD1aCV8ZJAl
lt/ZhdgbGSqxI83kbYcRX/EvIJWLq9VYSKkmKDWrz9il5/8gplrVlg+LfvwW+ORv
r4ZCGJr5BeKbQonxe9tlAtfZM4a2uDSnGJF8AbKMsqNeCdniwH5GK9lFEBgt5Fdo
K/+UM56sqfeWtcthF1RchZid1R1mK4q65SpfEHvkaZVewoTswlD/JCGDNMzZ5n7O
kXIea55w2wu3CJQZH+tMptaDQtWHh/t0+w4qjV9kH9BBHOEUaZrEtmiRqgSpmI8P
EwrOW4Lel6if46Z/6qJd193L9MsLrcvVN3Ab/zsecJg0S51UuPrj2QaP58sDV0Za
KWV+U4wWMqfScqHAAv9NduVS60Y8bfYuSHLdOodeW81dBhBhx3k5uDyad9FJoXtA
YAQGcP6cpPBA/WXXcF/pOx6JoFoJpPVtuoLuwTlzrJWNQaUX1mZgzm3YzOs5ld3j
iCLZEmSnZEwSp67BFaoSaLIVIUCDsBZdhsiVV0bNz+h0UcYyN40iFYPIDKOCdfSS
tPNrR9ZB2gFVuPZHaAdE7itSQ2I5PGXiABdR0JHJxaN7LWqxLj55X3p1mrhWETdM
+s/lhqA1T7GjUOfTGtGQjNMGgtMYI+z35VHaWBGS5zsF17oqmnO9qccTLg2CY40C
U2R16DWHW88obba8Nxf0UhXX/6kWy1HXAzz275XV2u/WspeXwK1sbWMXp1OO/fl6
2oSHQhzJ9FXxtEdwjdlSKiQy8t9OrtRMfh1jEjh16zQ4avMBKjaPzFFE7oQ6S8Ce
uwgxgdou3jTIknIxijG4c0Tesfl/jXFkVg/v8NI0zWO++VKwtQG2pazPShckjFeP
fPY/0u08bOnpBVFrOJy8CLmSQVXllNs0bJ4K4yieSI92/5DjIEA2ftnT5fcaTOc2
JkyHTNgRsSe6+7wJQb0N3mFIMwDYPKODKnOpgqjiauKrcIObizRHu2ukDjdc6Nj8
OlHZRgn0+mSAIrrzLFFyNZdVGEdJE0dSi6rq6MPCrnIJKYtfCHWvjw3fKhZie3+E
ZlCkKl/ceknTQH/AOlZDvslcdHTqQsTQPuop8JtU8A+VfOaZ05koN1h1f+H6fRrn
cqGJ815WHkfeUvjqdbuphhrdKQl1xiQZjhpYhEmwuGTQdyT6tsXqMHLy1oH8QPRi
PCtt/sqA0pVdFv4xYwvkvbBUKtKAj7cMC/SmarjtvQEDvuawCzZi2DCtpxRAjpAH
R7bSHKYmPX3V/d88sQmY/iVgwst64FY9k5GZXTjCl/BORf7Gw0uDUNZ3dlaNXuBm
RsZhyXlmes/ZObc9MXlvS4JS6FJwOKcjklP0mU56aB5qHqJ0Teu0mLRcR4YG7zTA
Djf46AHsM239gr1IDyjbgFi6xP6J513x94lRSQW+2wV5OEeSI/Vinj8OOelxJs6g
2LFGumA8fyu9E+aS90Ldp3DOu/vTbYfpyk5t8byPLHIFitXBrpphR0mNzppQ5O8W
gtTPCBBXGPCTtTETIF5CXSziiMhKI/8pmYAdNeGzGuOAvCLGdHspefGnEnlzLOhC
kbuFAbWi9s9cU4oqo9hnE9fgggDPZkSDgFP9+tPguLaGAhGZkGYuQiTVvoyE1DI4
pEbmcImDU/7GdrS9oV4p9gXfdll7lhLxbGOzNwlgfE766IypGZ1UiIqZDXXAT1eb
7yfciAF53OC8Q0uPznJqBfOPcHj2pijb9Zm0xxoaltFYqUvlbDgEdpBoNQNA+D4L
5a2yGCojrAAdmwZtKkG1PD8suytmLiXaCiGZKysVNkZdIE8KiZnnd8SHjhP26b3G
7J0XFOe4Mx0xBxwrr8B6VHK5bTzOhpwkJebPpZkzSoXPodsS68qvOCRC5o7uZ8sE
66ct/F8lo2xZtDYmIip8S2Q0trIxSivJ0iZlPYNQ8Kxa2LsneoNi/pdb7ddZdK+6
VzwD2FhISrFePyBEJEBHlGzpwXqr1mUhUcek258I7RLEdtq60bAophRKV1riug6D
F/fcJ81C65FcmWTiJC/BoMwYYPQL5Qgjw+vbZCM0lxjdqgdZhHP5RpJH15EBOAZF
Ghe2ChSV1hRDQuvXvxv1rADY9+Gqmz9biWZEsObZ2oHAmVMKvOluqxrr72lzzFYd
GSXbm7Xf4BVq0gDJuArcvUo8HOpWq8pEtGGdsR3Mcryqk0z8nL+h95mokHPUKjCz
Ohkdbi2aHIQMI361OV1jCesNFKZ2O5Jhqgkir0DBoG2Ez+0jPzqGWULYaMMBcmnA
+OFwCllhXUN3apqmmkoUXZyGvTijzaF7/5qLo6/QInnjEjkkNeIMHUD2GSB5XxiP
wUCm6a734V3xBfjvtj1WeuRCu3ImqmS+FM+CFjvk+URz2NLBTfn7g4RNkSowIay8
GG9Xdl+3PfucFlE2HVq9G6AHX5642Ja+XRHiJ9LBIq7+LYKzDbizxe/68KZGGM4A
sZF6OE0wVF4Sc7D+cQ+IvJPMPJOk36O4LRiCUtPdR24fwcP9WjRY8/UDmBESZFVz
uY55Yi3dbmTLT1lwjDD2bmVBjBpzBUqY6A+JzsFXHN4108QW6thc2H6yWVyK888G
t1dN1+zC5V5hbiXXt/8Yr6W7sBCDFZ/Gwm3SndTcso7hfxGb5D/VGQAXS+1EM+Xe
GFB7/9hjYxsrv1DCDe7s4U8Aa8FlRFololEqT90UJ6vtG1uQIzpb+cNUw6k85uPm
ZGfXowVj7SB6Ifvs1K1qABga0ggiac1R/xtaGvkQq+PE5TI3eSu4jiDCPgRJt+jX
Mrwuun/gdFI9bh+1I3gq/j19m+y77OTHvQjt2fwHQ8YK1GslO+7tkq4usl/3u2lB
UNssWcW4sDxT7X62FNQsjG9LQojxep98X5++BHeX2BmV8g9H2tKHKOGyEzh/Bx3w
BIcCk2xzFDGdqIo93zkTQnEFyB5Um0HW3UUSQpuYvp+lyY69iNbxf0zculhl44qw
N50HUE5PumftkHkNqc1w6xKWglNj8FhLpyrWC29C/TQrausocA3fcBEVXyaZcnDX
rXhvtReevhiKjoCje1u0fifA/b6avRKMBeBeTLfo5CWDftCz3NNzXzvh4rIesW+7
w61FsV16EE9of+EJfnxGnNqCeAwIU0iLefh9pkZbHT3tYMGDWhHHjgqGGGAKxO9b
gkiWrhw7YFIGLKVFnlaovV7YvcsT5McQEwYqJ0/O1zf3lzI+6WkdupLY+gwKqc/K
m1TbwBQVGU7asvCnrmNwzpc4vNpUxdHFmVZxmm0h5omowVT/9YlkB3bSi7sANp40
ubpc3nv/v2XaBkW95+QnoIcVzzOrMPXnFX6yn1YD6lLBnBs67UAHBYNHLd3Be928
LEI5i6pcjU1xil+67EHgE0XC8PJHLx6E7I62G9p06ecA0RoZ9yS/nn5HdOqWZPef
9Z8DmoTjv05GfpaaVUtr9AfIExswQsGI2zhhTFIbn7MZ/XpgWlY/qyAVmz6m+O/k
DyOXjhutZ25x7pLiaMKP/41SzPG3hV2l1UQJMrvM29ksfDzwoJwHHmA1Ni32V5uq
Ii74TCou1y6vMkg/q4NUNwJH2/ur12fUIDWELBZgxxOGscGcQmIJxQWSc5r7FwcJ
fbJRf8SY251YHC7wMwAK9Cwcd5QPhda8dRmbr/3gktJztGLOpHEnACeGMCVxJ7fu
4tNKbJdbDOyS0LMDO1UmCwrcGCOwXpjiWrTvhlyBHR4ppCUaSpgQ9T28K+2O2R6e
wNFZCbncZiCEJ78IcWys8g8MWE2ZC3JLO7Vy/Vf+QroF9FIR/37/h0ImQR//jzMt
TKLSfpP1X+KigkYW6VrCZSf54sU/hfWrsee5L9wyNBeQFpV15Eo8vYd5aYGx0acA
kjv+aHvrPk69k8yyaesd9kkroop9b9R04RsZUdHBRE483Xue4zvoEbJKsqiv7j2V
krqCWo34XhezDeRbOEs5CvozeaRfFhcgWHF9zf7P3bIGUh+l/SIW1n/IzTsUYIOw
b7k0p5aAHsB06FzIpSxlMf15Nb3gUGhXIS6LuR5g/8Jh0a260tEJQsL766bGIkzo
yQZiVjfMEB76hkOvBqv8yq/iehUULxTYezdbo/R+veEm/qBPfjsO8KqCjoi/cbFj
etk4FCWGddXL0jlpXM8EugKcp3Sh+bX6Bn2TpgtMhRSO99PtdfESiJB2xKRzlW5h
QkxtUvR1TZAAVPEewGeBuNF2zxl/Qbl/VP8+/SFakGAPZOxE8fQtStAlGFz9XFjZ
oAxZrw53OsqWFfZ4SbpG2xIol4RpNswx0P26vovBUPh7pk6xWFH71idaQqvST47J
m7B1cgYjzWerDa1qCsoQqAYNQDkQrcu7ll1VF9HmboM1guoWmOE1pejlfrsKGY9f
Bgw2BFwK75I86A9C6OU0TXxDD2+GBO6tPrSECN1WmwheL2PiZ87v5jN673VFDMTG
aHWzRIdtvqGJlKtzMnamACc0P+FHh8pZYHy8yW63ukRrL5uDDzKxDIqy+lJboo+m
qRau5R/UHZkVlJ5eHZg5ceGwWl3QAhKeJiZfcncKDH1tFw5eqvcRxQJO+CJrbFeF
xIQrRnfObk5lORLnkbOAIyCr798WEBpr32cbOBuJJao9wnvdOWJE25SQvlgwIKbp
fjbg4JEHKDjqdDFNu9SLxhenIx02BvSb38GL4TH6Ub3iRQmadYZ5nAuRL7601k9P
UkoAdH5I32jI+3RB0mHoAZ8gvVfGfnXefOX3BmhPL/qCJvCkgCuom2rXAg9JmOoO
ijIHTnkzP8Wb4aQ2SxaQ3asFi+xjqfp9gt22qdjcAQpcLsnZaMQHF6pSdkPqeEo3
/UYSUvVxM2X5dxT5CtXbkl5O6nllirURN2MNQVY5ZLlzqF/hVh+SeEVbLcdFCcgR
+ugGCxoLf88dLUlNb3k90WuYD2djJgHHpO7L2iHpDFFKL0bPOFcrzAgVSjieIvUk
NFqGK6NrgJRWjmDB+6zeAgVvrsFVp1DIVmaNP1MlLrAe8IoIZN6YYIw3jHM7J2Cm
K/jfgwyN3UMCRrS+nYmIgd5STyH5Ay42JsdA5vvLO9O2spn9rNTKE/+GAz80hGGr
v5/T72W9LghYFNL225JebB1WizYv2j4DizQHbEpnDyT1zGNZmSw6GKR6do5/OEu3
GbqB7R40HLIYSChd0DwRelJjFhO5DXMDAw6bsmoWSM3G5yet5R+cI8b+SrbSMZIS
/YDfpauIGBfUa+VCJ5C5FdJaHBOXXsqTjj3VjT/NDsjZGH/un6Ena1TW5nrmryqt
WpimBxC+yvXDZFJ4jNrmHl/jp/CfHB79n771p7aED1UHwwI5GoHkitptQGicDafQ
kHK8ISt2PBZUBDSIpnJyx4wvbmt/OioZnhy9b4cEZaS0DsaAIFjhMEoTjBUYx3KK
sSwolfNa/XYYC7PneRUqwsVpLvdNI/OAenfZqr4v393AWeyx5NJREDIBgRAgWr3+
VH9p3CDXPKbHORi4cztb5GnrRo0/zSX/ScM1DY41/I7b3Bs7nTX9kTTQfS4gT7zk
0vPSsaV7lUV8MKUZGX3js7/aIlAN3rOTH/NtOJKAV++X/RVFYCttVjYVnRRBSpWY
I9cACq/JGbxqaxRLP5hZqfC+A93G0qpgLHBsC54g+brbUibLEcrMSNC0kxLJDwI0
x8qOobW5Xg087seupGZZeQg7YVCrdqWTz+91ce7xK53hAUxRel8pxuwUkxDT2YW6
SKbFuxa7nQtla/e9nvwcB0oBIfUbbI9OrqthqhiOpQ5TIjMlai22GXMJMsNGkaJB
sAXXvZh66acw3Mhj3X0/ME/fUOcZKIG6FMbaIXnzxfkBvLgRBDw22TS0vBdE+RY8
G0TONYeUU/Zrlin0sDfbYMrFKWlKzW7NvEKyeCGapFx0WHpBCky2Q/1WTcV8ROEo
qJeCZfEe9neWDboWNLaIJnM50zH6PxaJpVYZs1rfqIwxmxXQZMyR2FO3Yevjo4BP
GR/+YA48i7khifsVrpStijvTIAyJU87IAVX8XFt5+uRP2EKhj5yJHTdSDCQQ9qnu
LzFDib54RyyjICBCbf9fjogVdrF0eUajdGFmlQ2FjHrQBPZZR2Nb4Ru8JNS6ZqYm
4sAUqXgiCp+jnre/Nf+LpMBWKht9JCr8SSNQuvSDlgAWyuAr7WPYUJvglvviy/pn
retTBL6y03U8cDVfOqWjQ9ZMwqq2yGZCgLWt2jf+TcuadJlkXgEHti9OFnICUOu8
LY074SRmljrZrOoQBlb50IUqiBUJwsCty+ruIeIaeCDnGZhDf/QAWUUbSnwyl/T7
KfnPHvmonsGZ6Ay5JC7I0zbbgaVdUMF3I6IqDcwj6/D8p0czxmgIiJ5UGfjk1UDn
aVEjF0wbluSHBdJBkSrHxIRia56lor6tCXLXXD51b2MdbfdsZkbBHubJqSbLoTqa
nsR1jcoKZ2Wg4J6AiVFl2lDiscDqDk6nIGgWCAGANMCts3bibUMs5tHrLLWMwry4
FBZHsBM/WJzKcHqpNYutxWB6u/KQRPaCJ64xuqKW384G0aOo1bW320+WtTaANpfJ
U3v/qy5gdmmGizIP51ZqVQ==
//pragma protect end_data_block
//pragma protect digest_block
rKuzmLgB9na+M5123FbqQxpKTGE=
//pragma protect end_digest_block
//pragma protect end_protected
