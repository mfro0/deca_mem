// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
a9j0tC0vIbS9e7OLB6jjUfMuwWRapEc3OVqiJLJrEpF7YySDli5oFIs1haZyVuPdMcBkuEewFtfT
/kwsv31lvgFiVGrfom4sV58h5ZnuxykLfnyV12j4+TccMuUooMYPJz+u8+bp4v6XAhYMsPXvw9+x
SKCDGEOstVdzmDBF2ijOxoqDHmR13vbhl2SlgCdXDPJZAylLrOSiNrgzc7fjDjkRsu0D9/DQiMBy
w82+8d2DRxd9smH0zxuD19ixm3U1pu3V73KUH99WMn4co4Y4Gun/aZjd3t8VrgFF9RoNHp1K45Hk
WyBoY+qMSXluPM774LsXKPCg2UtXO5gFitB6cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30032)
1PtHYMaW/QCRigHEpcTIMxBj9plpEwRSQHVMOda39+7ZqLV4vUkZbO1vIky7ii+FGebVdm/tg/2z
EQKLJMO1LZ2L5YY1MjeEyhKGA2o298QoSS2i9+O9mYyGz1XeFQD8G5pxYZ+EYhyNcVhY6KB64XYx
6QwI+MbG1RuMK4PWaxsgLO+vmXwU2BQzgjo081nArfR7gGy49n+CcV82xDLRsSpBT+NKpmF9hsuE
gerrnkFzYdEAX5jNegziJtLgsiiY9il+Co6AwEpS179FUtzXUSA58M6gZsg157BZTQwxUt9njERb
//99ViH2Xo1v80p+ZpFnPrTR+K/7fXJ9AAiehOvU0hyW3dtFucRKpq88KYvqyY3aYPFLTenMUn6u
QXzouzs2vebQ6307Y3NKt7BnO75Dyu87L03S+lK0CAR9PsIfLHhHOg7eNsPTNKzg6voda2PhCcbQ
Cn5rRxj7gFQJVpO3Yg5JLLkMtwB+iewbrfPjhD9z86HWVrJeTUXIyJ7DWl0WkDtO3FMeIkW/l1BC
rC3s+WsUISV5dtGcBj6NYABZ2w6Yu88owl3pv3u+dXHWNWAq9CNpFsnPMAgegwtCfDxoL5rRoYVh
8TrzQFG81021JXu0hH8z5Y0rPQi/J57KEuKswdAHB9yJHENaDzTd7QAL4JKu1f6HzujvHZUfleYi
Cq7TbfpBRZ0EVLpbi4ZJSf3PEOknv+QNkH4c3uGfHuW+ZHjTSHm52zwMKlYpdtqJHZzTrnmZ7Jvf
arfPANrIMrOZINkU6MtMQtnDcJ2y+K00cZv+BWDZacV0f6oCsjKl4LjWHEu0FD48GN8gg6+qfwsf
2O34ElTUWSJPlqGsQ9IuxZI92MrkHtsArftJqzfiUmqWO9mWy+oSvOs/WgzLo2swBoVxvxWQo8+X
1t1b+SyVjZnbODCbouCDt/UsM76VOWssP6qJg9Lzu+9v8K8VQ1ubzGh+tAUiEQ68+gXX65rabz4Y
8TU/+AVctGuwUfGPVB6nfwdmkgbKOGxGI6BT43CVD2NacW9utyB6ddXcKTaXkSvVF95Ar+XkbQ6t
47oAcB9HH3KGUZyOdYgTFDP61JrXGpq5pKxNvfgRa1x4jepLEZAcfJy4GdWglK6nFnAcFhSNT6Au
HLkD/QY8kYvQw0+8DOaKVKPpSacseEeJHNY+FcG/bttNUdPU6ntHJnyBtNqpYIa9KphGXMqvalP1
Lpt+IUd+kU7Yvl5Q/cbNirYboWSYqmny5TeGzKlWa6GhYOWs/ZWHF6trRXAJ+BnoZbks7ZHJO7n3
z4NAKpjme4MqC6xxT+fBiGpGE/TFNzZsv8ccQ4/gCLh3gctX0Sx219GkaneYSG4wWIg5QO9GzEkK
//JFhjemQYPuAUD8yXRcl4bWWQEnw9vCyzld5FJ1vnE0dJfq2Vu3O4y92lsVpanqJT8Zpu8f1ign
WRZ0xbxy4eOvgNK/d4Ps8nTlVDkXEHWtjAxhQn+At+jMumtCFkviwIzwVSG+ms4xCnwXzrBQ3ReF
ojFETyu5V+wCU8pmJukYSNXn8nqqJRMza5Rt0S36s+6wudAubxI3TlBfnlGB4DZ3RgcdlQDX/+GB
JypmfARCV7/iI9CcxNJP580tX1S/f3OiEOGEo86OJonWgRX9so1bC58DCGv6lKmt5DLuGkDm/qvw
jGlCAPSJ2BncjETUODy7QSCS0FR9z4DQomoPoyVdtAOog2c1X0/izrPA8ojOzjKYVJM9UVGNnYvB
qY+N87Juvqtcvyh+8+dlT48DG7pxSMsH1aDqSIPDRhIyA/pWJh+mvJcdI2tdtqGqO73HFbGdE8Qf
nlJ5kkhDzjfQIF44FjbDyz6+wgxkeM9JCSrel2jmLwkb7mfEioBQXEt7BjlTrTMsahXx3EfgTsqw
XmZLDijFuS5H3QRGme4PHMymaqgW5xTHcvKorWjgbOW9uwa5RjWP4Ez0/dBuLnt74ik5IcFmXdD8
3VYrkRdCC1Br0NnsXNTkSMEunBYqFwuD6J4pHLjFHwCg31JT0ZS+uhGq76W5hE6mlijDxOkKSCZF
2UJKo9OXsZy5dR8q8bTHinn9yUHMLImJYfd/0BpRD4HUFpTk1MvRQkQoDe9apDMWBYLwFO+n6zOH
gmFRU6gal6zLtNi3Y1eLamDDACpxWwUNBPxND6ifti8f9Hs6M8+CO/q/W6vXQpsNRoo1mYZhUJBA
xve8AvU1IRyUZPqmRRKN/zs+aDsGN5dPJMv1kyeAitpMH7Xes8egjHJnZIRPLpPmD3BVdq0LaEk6
cSH9LNTE555W2jk3WncLA3xvSeZk+5qY7m1A41wtfLSzqs+3JgGtlwTw1stCxcBBIxcCzIWrTOSR
6CHJ+H+rctnvWb6QDVU/CdeTokTGWnkeDUSMjBz85x04HqqQ8YXQR5SLtpTsfNqrNwqiuois6vr6
dbuiCqL0W5oJYlvefwCT1LE6xbysJ5SlHMDf0ew9MPVO1pSW8dl8vxvkBEmUXzm9QkIAMctvtQmd
NJnf063QFmku73e9KfS+XlF/YN7tBhfxZ1WiOXmRM7wV8Q+asEkwhqxFeSdJwR49eA0dFAPwOdcR
W5bekNirbewCt1U8cGPcYw+sl3SBNaCTv6sx/FTZLw5uD5VQ+2O4yF2i4alzpZXT25k/oOTPqZkn
SV97Bfz4JwKFyC521UPHdvqAKwXeaCzbXci11vmY+P8DtZ9Dh4roIeIZMfRYpXWomUAMtlAqZJmo
wW1r3zXxCd+z4GWz22O/OMs+32MUSTqFG0BIRdmwryg3avhTS+mB7ydD0Dl6zg3PpKQv1Nsa4A12
FArmEb42Mlo0bPHKVv293ErP7tTuCE2tAjwDqtC3EKFmoaD8xfPjBHPTNIYjH44761R5xu1v9Ccd
744bh4ikcdwb00xsB+tcb1tm9PepPJxcWA2hRz/NkanJyid2r9OBYJf8uX+nrg4bE7fbbCfv7OY+
SCxTreeBlgQKkCYe3Fr612EZeC4sXH17NWVdJ4U9H+gCY1UVN9MGfPkRoenqInzmo7gRfTis6koc
33vGJ2tZQMI5rqgWyZMv9ehf4VYXg44z2SKWV+ol6gT4MphXuQ1ITOTszT6TF1QWodDW5Ozxvbtc
LICIAtzXzbDZgwyF4I2zGr66FmkSDT5+IeUqSrKkP15pzYHWOyYal4ZBaQMu1mqr2OuFhPUXMgK/
eYME8mOIGXM3EDm3nsHUaZQMIzq66IdmDbQYjPD6n8eQIfzyueL867gP9nsSt4hMK732dYX3iZt3
ZJnkqwyIOWDFgQk+wN3pCkutw+dTtUTE2rnfuo1wp9FiuBabjvDVX7zKxJjcRCnhg2hGgn9ojMFs
RQ1vVQIpqPKEFR1i+lT5NhlVIQju9as2DkO7wjFuK7MHKoKgQHUYfzh6Lr6EjhSQUgpbR5yvAuZ9
/f5AMbiltsKz3JUKdMvpJHC07w7w1mTn+rX/wZEY+tJkdbbC1qkr3wze8M+lPN6Q++uJVPoNdD/u
blvkEwIQRMwmqptpswtNjjDyDAAukI8p9NkY9MB+FajmEcc4LSTsDDteF+v4lNDjXRYcXKvWJDOB
gnnBsbfTlkqVwbZRxJcQJcrOZp9910mOUR7LiNicJMAt492LiXlslYymNv1qLB7yZ/8HoPRcjcZS
LRup1G7maaibDiwxEMevh20udrBWQFbdEkjcUa7wgFchdLLD+rWUNNt+W16mddkDqPFApaolXT6F
2A+mQhykhV/12NsqHaq6N+AjvS5p59QBmj6LmGn3z/LpBpvuErZnFDy1ESx3LVsdW0fn5Kuz+r52
EhGohNFGPHV8elITIakqKEmGbEsQ8dsdU6oakD90h6anTg35vArhS2ELMAR7/2obcioNYm2IVFeS
6riiIE3F+V1SVBmoh3sSg0zYzpEiO5P4TwHjcUWQWsmMAZYz8hdvKGFBx+7mime+ypn3L/93ZvIF
k9X4jnn7Y3TiarT2979bMgRkcRKA3+qBjNTFLgchlK5ZFLTbuP1TMadOhugyP0LU2I6+haNRjDcv
ikkc9QXj8mR5NyGERfdnZeaHFiTtyPKXnqk75uORNr7hlA06K5+qU+dEVTlC7/f/YQ9uuKL/B7HO
P1QXbCN1+nEEfngzjPavSj8UnRUtXN1eoEzi2vrJM2T8ZB92jRbKf/dmYgmMg/TtckMJXVq7VfRz
NFSd28/U3+cH/3DqurgeP13TMNZGcVxA95v5+bNPC/DrTD2vi5cSvrSsngfuoRXo+BSCUlhtGTnm
gGWXYf4oEvlwqDVE3hTJ+2XKn5j+Wp6UT/S6U20d4gz82P6LW4rJuZFb+E2gNN2AhC7ZL5NnUrqz
LTCovC933a2riYOAIiH3Nh1BtWSzAtQoeU7HyKe5RY3eIT8ENA3veaB1bPkuxfF5LqBYEKNUHdiW
wigQpKhIwg0Q/R6kVWE0w/k9HbosrtYeigGgyVpQ4wIfTzdu2o1Ue9AeMa5z30KTfN7ziBYLSPhr
cJ9hIGwN45nV+m9Wg/kkflX/7U1SzZxk6bABWCq9X9WGQlo8SEE2CA87fwpgrBM52e4hqBx2UQl3
DyqCGFemrBS0dukRsFL0xD47ljDXp64O2kMXYs7boigIs0vX7rAYzHc8e2x92iLXXNFhKvK9+g7t
oRXh8V15K7umkUKN1BzeXJ8x6rjrHErcptlRCGdvav/+pV8XGGG/wnHdKex5qqJZv05q76Vm8cF4
aR7GUnKjv7Q6X3WKxf8Cg0Ifx0+N0s5mY6swFJcrOnxLYwM4oPZ23vvOJeEuYOdzmLuHwKV59X6/
/Y8/eo+BwNUBePd1HXSZ1TuaWQPQioXQItL6cybKlm2mDb/7oqc3aNONgKLVQArAzcrDKyEY6n6F
qi+V0Enp4+nvvhBEjcurryxhULEF5f7zjSWbBmkMMRr4/b10OhBac15q+uiKKH11eDgMXraSCge1
b+eFqlggClUywtr6YiTWOf2fVmW94jWHgGnTq26PVMwcbR4THE6t67VfYhQ/j2x/vow4xlVHZsqf
moU44ptAVxAxfP3Llv/ictOCbIVTF+17Gkrdeh3XnDcNFt91wiJUSZxgLGYalWUTX2uuGtv4wUK7
depNpDrVObaDfz0/S4/aw2mzELdE3xgYeh+OCKvcjrwo2aN45Ks2COAONdYJoZbi8PzeR1rolVvy
uyZstByk7pizxlw7QxzilBMuKs4FnKbPotmmaubnaqB6GCiqaRnCeS1wHfCcIVAmtWLYB75IppGy
BGc5u2bwG7VZEgYvEXtuBL2hi3WBhonIk+azytun0UdVDS7VLdniugP3UyV50coHrWdZk1GRaR5U
AZhwZHLXzuiR4RqbMmWqXZOVe1625ESGw5c7zVsMck5ninOXLpN2Em3PsMQ6A9fUaC0C90ArXs3W
rBQdrShfz3s5ZM0AvHWiJD6uYjHxG2hna1KjtmkGGLFKb5gBGjiCRRmfGYyE9FKKRxxfDunfIhg5
d/MtsphUPMyntTeZ7DV3zyQFSnr7RwNbQktd7+/UbrIRQSkc9R6l6SqzEdphsl5PU8aXXjohpF0E
CRO5t6fYLuVuxRT3fbFmG/dX1n+zgmE6SylQVfV5gQ3JB1jPaLI9Ytlwl/4BMbop6+LkW8sh3zK2
hMpHRrQNxoGYb9kt5Ls+S8nR8YKbJqRgls6hJCOV/r3QdoJrnteyhes8W66KhtekCpAGDYg8zUS/
cJFQiSD9S4QhU6HM3sNipKYX5Q1SEf1ttoNfVfNn2jQrQor438KdC7u5LV0Q2EYK/dfpobdc2lTI
+j5OLzAGr9Z03Z6ABmd31HHiXBbcsww3Zbg8uBDiyuRK1gW5/ESrTq4Xrj8FNG5XcHUb4ChqZYRz
UJVVwSCJad3eK81IwbCXEPL8hMrtinVmRtDZqqGpuUfwOXi9rNPWK2pDxC7Ua5B6MYwVWG4QRkKF
aMEGt2MNo1uP+hAE04WOpOv1XGXVWB+SsnIMwNUCib2eBGAxnwdgX6Oi35N2QRtfT4bUcsAojkzy
EzGRr7NgGEKkmq8g1yuLMggHi6H4XgU7ENGC2fCBXG3qaBu/CoXEzjzVHyPGY59jXtCXtWDBsADJ
W1UXGJFod1t91g7iy9Ubhs8CsYLkpYtdHrHCyzyd9s0c71KGFluniRni3ZI2/M6sukQxpdgmtGcm
0lgBsqEAEKnZjRLTRmgENGESqRLHT9EASTr15VspOnQm3nGoU2iUmqE3EEQwkZ2i4yjY5dk8WKsq
CFlOckbR1DqVbLhSH/isYodpYY7hVa/O/mOO1iv60ipVSEONZ+s4+7R2xHD6Ic9YvSlvHmdhv0Sp
Yen/xyonqAJrVA61pwj7yDoK97rvDISZJt8K5r3QJIKZkjBMCY6W7MtoBurb6SIVD+SnObznpK1o
7AaMpt+Qti/iSFhqKT1x4ufSv5jb6QBDhK3O8QMqa12W4gOqcIqkw8APsEzef6aIk5mFGX7GsD7l
TeXMhGVpkGUCAxFLtZ1WCx2ylfkF0vFv+pMaO/7ioXjU36sJisNMdBNJQrlxeEBnCtDGpQzMEU0p
4H/W31CoC/gw9N6DX73fXJzbi1oyHJ4Kd3aRZfXRhotydmPUjdmGv6YnXXaOmt//aP361tI+s+/y
Sacc26RVwZM+ItdeolsgFQpsutHpfcAXy/IQWCOXSNOPJwPSX4MAjK2y2rfsJozDOufqz+VD4+Si
1f9AjNTvW607CMDnr9Qw/LOQuDEmu2Zk2yn65fPZiYHP1h6lSz+z4tsjSDsrEQ7IrhqNLq0sEaH0
QhS5AU73DfAoRSLd6oEot5bHNNOB33j1NZHJ/Xruz/idbVjkiwsqwbqCSlN8cfXIhfCFiu6xp5j+
oHV5VpKFBpJC682HvCMLUrcwnCuOdTnG4avG+xqrmcCI5KhJoQDzxCT8II0VgZBHkEvhl31lF2ly
FvLgjgleMQivtVhX77iUxkSLU/NfejDkosjnAZ4Tu9VBmgWShQtCNknJ38/gUS7OvI76bjL+au6g
zfaGJsT0RYfnJJPz/eb0RXzi0F9MdF9HwioGECpuU+fZGjC4K95yjo+pq35MAMhG4yjAJLF+Mj7i
2hVAEcYCgbKllKbc5Ekj9/PdTOeukTYFchZ5dmzyJ8ULAr4ZXva1iOSLzYdd5MiIqqkEXeA8no7f
NJ3qp6pLkGxhvp+8WsLSM2kIW9cf+Uhlr2XK5lWkxja9LaFTqUy78VwzREpy+gM2K4LbzLzRZY26
Nuuup1gYIbPjrXh4WDSmQvXG55zVUNUZeVLnsm7xmxfz1EpfZxDE/guJnTQkEP95VdDSE2g9Ziw4
DyPvf4VJuys0FauVy2V989XIcQSvhG4QhYQNQ51PgXkK2DHSkDrs9oqU8vKvGcQqTzUl8kW+BY/u
aoA6wGqh3nalP0qSoxzZj86lbdplHG18+DLVGwgqY0rODrkNIat35eEkTswiLyYret+oG+zOecgG
kkUvSoN0BY4xjJdq5cBjRsnMylSTt8SxtOv6lhOgyF2CgOgl7hiNIu6YpdBZhXS/ZoNzj/0a8hk9
kJMbKoTXaV3xJPFdxdJWZyRKi8ErkrKLGBy99xyNUp0zxXcriudG8oGCh7Azh68F/9s1Y5H9+MNe
8YlJrHavIr4/Xs2xgJIVl4+OoZTaVe4+bAkuRc8HDOI3qR+pD+ixXqsClDjGy3UASUbrc4DLDv3/
k4J8huxZDbFUNXSz01zVsATbn1NVge2488dhNI9Nm75Zia/ex6UpJsbijTZTeSx8PcZYi78uWkUx
J2NPurOGUdtOOwXmqWVfwhhjA/+AW5PLhdiT5xptsjg0mAKagEIajPEpGBpiNrQ619jY3iv2vxQt
JaS/Dp/dUJuFrN0g7LcdaL8EiUjPyXia6bNJe2XYeBI8Dyv+/zseCuwWqt9rRsIp0yJo3ZWp6Pjj
2FwoV6+i8gnWD+Upm7b6FL65X0/3MIpeAQrJYZljhbTL39QaIhaPjlSjMzBQlBLt73eSjw1NSJ+7
lQvdUAD7nUW6rW9/WQO9RHyZhvTKkgraWLA2cUtHNmfw7h1ami7MRwP4s0jjw8QY+rqC46wKUnG6
yGozzirne3zszQ5X+oMmMBmGyjOrY6sIVIe4QdnAj7cfNpEFfKUgtI9+hDjUb7QMjX8ZNusTlxq9
oJfmfbrXHWrONH7OnOAOBqM1sJvKwUgk0trC9YFO8PK/FJzvGP7Cf6RA+WDy68yoNkWEAs9OflW9
6Uduc8zKcNO6vsIbI6CmN8jqQPZf4VrylSccvsqnGeBnPAshLtCfjveP9kg5NQuSKwh6NLRjnKUK
edCnIF4O/hbEHS+50yzxMVqxXUyEXRr+Q7OzIrra+fCJA6/U/tEJo2WgV0i1OTXg1N+TZ7ByCGHi
ieX7shpYKzYowF2nMzrcy4K8zpGn250WWVdDbJUU3wlpxYGX6khJNIv1u0/SXJuxsxmBml7x+vCa
0so/F7MPH6/H6xV785OggY2CJPZAdaNHkfssX2IFM6HzOvRHJz1rOik3tZ1uSpYB3yhyfQ4Oa0Oe
txpd8mpWUu/K3FJZkCPIw6Yu+XUnxZ/klFzsnTrWRGIEHnbKgWP6dW2OkB2I7dVT0kkdoeYN6xfl
v4rf0Gxv2wldN/JkCHdnWxFvpFaxSweH5myYz3i3xNoL7oaIA1YExI2R0faUrPF1VM+3NE+XPQI5
HpwlvNyd+TsDSwdv4PFdv2U3JLNen2W374XsAEREknMisbA4MZLSipMD1hWpSx9B2ZS+z4lQZ+sB
ML71zUcS2TVwWnaf13dF+d6mI8twTp3A3HKV/dpAzRtJ4JiGr44O5FSfVldqnEFRN7k1tYOf0PLG
xHuhfvxS/9lFtCDd3/59GnFBeYIYNYPeW1YNihEKg/+27DExkT1Ll0fMEaWrwebljxTHNRhXQnCW
JvtDEoBiZ466pcQsP6pRsP+gxexuwLffsFviAk2+OjLCXQXmbRtIZ60qyaa7ibOdp4O6mAgOnbDa
qof4vu3mVUyc2P9fNdiuoQ9X+EO+G0OnhOWYhEfnfBhMcpRNAKG5lEcK6IBW/Re5lji3AfjtMgCD
QzM4R3VlWMNjQ6RkeqAXBUHFZSKQx2ozNhvv6a2glbNXfSXWu6w7+gAqUhxAOKHdseUXmWzmDvtr
3FQKbqymi7zn7/Zqc+gQiGluc0xCXEnuXJIWBY/3+wkYqBA5BPhIzFeFRWy0eI3v4v/OGdtfP4hz
YctmGxSc0TvzNvHTVQ/u3RbXYubayDjybVXdgGaDmESNx4DBhk7K+3Iy2Zf3pD6HAbllzOoIXxSu
8PVwcN6P2kpL6OGKLY+78zvqrLElW5DAuEqqqtlRcsqf0cWCb9TvN1PvByBF+iFKv4EEzRKO2Bsg
yvSUIbIHtYMMb3dUGDephl1cYMrUWSAICaOcsq3hpNkcrfrQ4q/IB0+orOGmHfscyqhVadwDQrGN
TakkcpO4cfRiHsegFSXeWE7hjvEURyVTlKK2uiUjwauS863H0FeLTmfSozTQmDi+BozGUaPAPBrJ
yqASUNz1E3c4zEGpxr7U+YztTKLedeJOliQsQXntXxIGTN+/zPgkqas6Juy3ZZDWBm2WTntwwPXp
BXHLoPthW96/oy4QgyM/3TXbyFjGqHK0GBgcwE7qeB4v3dOlGnFT0J4ZTeav7vJoPoh86b5UXVMg
cXhXa6eQO6LpIY1cSJqbpf/xA1GtNd6Nq/O2+NT3rnfDqbzpQFMAlJpHUgT+pe1PkSmfJUbxTKCO
lPzLKgzREq3uIjd7q8ue/7y9FrDW+lkna5T/lyqQhJq2I9XEzjxPHv1eXuYTxi/TRuypKwTNNPCe
UXP1hHQJMfXtaBjBgpAJLVpV4Ah3LHNeNlzW61f5VsTkgz/d6L6Nbgv3wujza0WewY5Wr1S7FDIH
hNUNOyjg5JxW1ITq4MT1IvUQ0u42TDdca5dmkzxYMCkIwEP9s26NGslehmEtcUhLXKD7/mMxM+Kg
pRWiQiDEUEu8uIZFOgutMYb5U/+2CAeq0xu0YEtxXVKjdk658Xv++ih/mBzbPMc+7i29GYUC6FYo
U5Jb9c357aFh8EBI2srNgqley8jP2aoh5R2U/DNfaldVRY6l+1nBIaCQzHBygPXgH4oPqxZbVTDT
Y1vNVS/s05xWHnRSx5xYtRvJ+pTEnAgBMkHxfMfWK01/lEx/H8s7J6ppsu1+T9HF5NeZlTR0O5i2
9GngkzJIuSdFVVBTima7JMQVw6vq6Fvkjs9l4tlXfZn68Mjqw+/8aPc7kgvwMApLJopUc5fOOSkg
oYlgxHNZGGWFbmGSHKmQerneiOAVlGfg/FyPYSsDt2qvMm+kTKtxtMhNl9/736sOc4PlnZjxx5+2
o/fwczE0Z/P0HCqdGYKLpe8eeKzlZyDhiNtvkwtDj4XdhG15kNOGf4g+isAFfrh29Gys52PtgA7N
lcf6JHe4Mtwtx34zgDjbiV3ekbpt2ckOlLk2qNdpv9SzPArO7dGBAPfAYH34Fd6Eej0LNmWznNPB
ulEiLP05J6rR1KtLFHTV60ebGuznbwE/jl8mMemjJ+k4Tev4Qgm43rmfK00z5ZzxTa2Ea9EhNXGN
Oygx/I1QtTvzyPLfFtGd0kYc/OvRwvArBkHzXb3i8UPsw5nBwd2eqe14gZcN6NjGysu4O/C5Ppe2
hQGMkHtlr3ZvqirTWZ2AaiXLhN1D0QMUDktyIsbP/6/qtwctE12d/aaO2p99c8lCSJN69AbRgoXm
bD/v11/kG1o4O1jItAjyeZeHBT5DKGikBY5f/sxeETxm7j/k3GHWQfGHu5JbAc9p1MiIEkoKOWDQ
slvYRC9xlwbxXyHU5i83x6Ra8/OYTHP/ar/FBnhCagGW2qxst8aR1f9QRSjJFqcAEjRfAO7goH7o
KvaYR5jrvNAj8f5eMwUVAr0PMNJvdFH8+A+LSF4aJaht6o+Vbl0sf9mf8HtlMOF1A36FIRJkpqcY
1INeFJFJnQ6t+nN23qnb9vQ9HOz18eEL7NbClRm8mm1KU+S9PnoSrErzOYFIXMlf0c+aolvde3B+
+lazwJlL+kgGx0qa3kwM4RNHmORbDEWuNthdAhXDdSWU8XGLuxsPT1wMcoxnTQwXCWWAoJHv1S6a
oWFv0l/5iKMrWQgMYgtlLDr9aoEmqOkRYax/IkR5OuMKdfavzTZL26CZBkwUNbZat7eCaxQxTcFp
cygCCTmdntFz4biq/CeRF8lyarm62YqNlh6UGoimCyB1ctLyiWNtL7a/bAaBuJ6tbhudN0G9emeJ
Jms+w+YAi5zwI6uS6U9sDVj85HcXUkBJq7Zw2Yu3eCdg0vnhTHAVp1BPNcaAzRGmebfxj+9HA4e+
CWFo8G1Q7uoLHOo6FmxGFgSKYEticFGw1G4IcPfODDIn+uE5sCDCP1upJbEi4Xe4aGGJZrL+ZnpJ
LrdzivSRi/9nDsIi853hOBN5YX3x5tvSplbOt376iYFPsPto0rqqFU/tTQwrKfToILzAZjIl2pe/
tHnzhkCZgrVz6zmK+IJw1fdk+AnM212VlcAWBprEk5yFjSACx4gKyt+4T+xFVhz71MjAqEpQFD6l
W2KOE6iglVPCyrUj7aNfssSL10NmTMjQgxtB9/cqyWkDuTggG4K4HbkAPISNgg2ic0p/PDWUUCUZ
dp6kaqhRHJ8SB+WpZqGideAuxG3S4b3WK1HIGyFggvsPxHAwA3sYem3rF9R1uTgE0mexWiwf6CSy
7nVCL6qR+m7tYRmKGkUrlewj8CKhpewh+dIFJ+JYhmPFQ8rExTlLtfv+ng8lH4jpu4RXg7/VTKco
2FOjLqjkyLxhI84tuMktWOdgGAujKYVtG217f37QyvHUsU8pzYoUStjIGyX5/k1biauAVecM1ciV
cxqdFmVh3NIZB6dt6+R/JvTa6KaZWQgqrPtGS3h6bx9BhN3H5HrPBqPkOt4iwEqtqwUisppkZ9N2
78SFZpRRbDZjYlZp+WOBPO0PCuGLu3fMj6ANXwIfL9TPw+nAo28w2OZrGComrI2JzRBqcSX56STQ
Z/blkeMNf/Sti2mDqpSpcJ16LD/25o/KhKguA0nMMXle7RX9J9FiKyBDbRuULk1+VLplEZ+GvpR8
qryEBjjid9COxxZizt4ssQCe4p6hcdywU9HGALiwvuBF6pWbSgSm5hRuL/ri7VPh5udPqPbwCR/q
ebahovIXCjCK74L7OJ1LHkgF9QfSNVa8yIjwXFm2ic0VMOHZ/ei4JKe247ipmDmCKuhykSSTJ4FN
xwbDH7VrgsdTSvwnVtlEVB9YF5NVl1xU6GIkUQkoipPi3RzMLqchujjy1RB9zftiJxQDwpvGQgAU
s5fk/8rV9P84ie1zY02gBUH9/a2KgWwKWFH/N7se7fAlNndwi01+fSme6BSycoQkw6+WgSw5dTqB
LF5S+W/NH57p+FtUPoOL2ZaEuILzH84TWBMXEoHgRZQqgaO2W3XcqIEC0gmq5rBHDyBS6CFrbVkd
qvFaOBbnQLe457Fm304XdcGU1FXcnED7SqNeY2hMgxlR4RjdeQOYvvUl3ZyIqTqqlV2Nd8u+ZYN0
W0oMeL07lJqzn4sWoc/7AbWXQd0sRjAQH0z79YZpN8xcXcDEIvcrw+zxHpBtM6e9dQ5V+epIkC7v
tyAFJbETxUevXeLslR74ehEqqtYdPVw9J7rUiIArbtTB1PKT1bO1OQJOnyo+dNpnY6XPrRHzjJL3
jTT566VrwfxfAgYB42Qfd1xT2Eikzg6e8iApv8PRym34dfD/y/v7tjQwUKCzfuyjx2RhllgnvJyq
Eu4b9x5e5VXhCaGaRkTIB0x8IqX4qQtNoVsG7YOsw2u0wj7BdnrzffPbTUmhUEYTi6luE+JsBlI1
A1rjQQMcXEhGIosDGUhL/jn3NZuS8WIUyqsR7OzsvAOsTL73fDwvschXt49JrgWHKISe7MTb5Cwh
c5DS15+M97e2PzNoSJ5VgEyZPUGhsi5bOzW7yNpYXZMn5Ed0cJ7Up7VnExqhAFZ3oJ9rUs1dcosC
L1pZxkXEMv9wUo3zggxsfEletX7lNk4nTzXr1iImIWhEtq1lLgcijZDRnKbwiQBoVQWqgtNnTEIU
yMfLpC796R3fM8C6sRQDQU1gdo3EVqwsYmjuqj8vn2pXJdRn61Unr6eBF3ddYMT8R60WuxW7CmXV
lrDzRIL7cfr4FdxsJMGTx7Nf5qqjTbYCR38oFTeK9cg7LdGjv4+lqHPFZJM5S/UHMtAJ8+M8kM/7
+JNraeabP+aJnlkUea/Gr6tTPdaZECRavtUShzHZeb8Ejlo0Eo93RYMj1YUFTLPTwlYsGNTHwuF4
vUXIlo4+LJzlM74a3BlbuqbKCGrXaMi7pLw5+3p+rUPVx1mUVIR8znIcQZZtKPWGlkGv2shCMO4H
2r4sArZzt53gDS8zQ81mGiOPl7ZihpmlzWA1FpoV6DexGk0XqBJ9ms667WQHIgl1Gwmx4VdBtuGu
4RBBU+KYJnD7s91OOjue8DW42WN9d+xu0zCdfBaSG5NEqUMs/i0QyCFg/7hQ/0kNMDSD4vynKZWL
53shVkgV4bm9r0pV3r275jpT/uZaXvXUWF4af/Hs95hWcCLwoohVwaUa6yvL87+coRJF6FssrnL8
D2CXI021/JZjrcEkLZk1EclPbl/PJJ4l1zg2vZLuXcCD/XcIeQ8vV9ld/IJgGMkTG/236mW29frp
eMR6Bc2VmQbLoIK9Am8VDuA5VTkYM+jU1aFz3hjPa5A8I4asge5WEWXzRHTZrNV094QTbwR2dg+f
FjkhULHQkvdWjiZa29z0mv1nLdvOKU+omaShDRz59U0P2y5SwsIiYr5kPkwXT2tgp35P8q+vGGBs
WLxYVn7AQkcArW21OO/rWmtNCXs/CD6+JIoLoAOEaFVpO9To1r9tLvtxsPQ3grzVDcChkBszGL+a
Ktg0Ds7qjlSOM6uqV0HmQGqeLaf0sPcEDWf7IVY2cFDCT6QaTbp+xqmc2yFmYYLgPUcG7sjSV9Qv
pshl0Oi4W/TVH7Hz6QOU6I0rmqJgqJ59EyqTxW57AcPQvzEXkFUxMsUTLf3/SteHcMLUX0/CsHux
C+4vgtxabla/85dLtQwf21gd+WSLY1Ubx5RdU23RIRZBbXXzFVUu6M+6y7jUeDnrBFlGlLs4Kmu9
gmncyGQ8npiSTz6oXE1+8qAaekZT+Jz7L2NvhypOZ9ldezbw+uxHUT4QdRwx3Au0J8Mw82qQYn5h
KhFs6nyx7P85i15n1O6+P/jWVClk8USEzwzLwIXfO9aPGt88sruPBjOEmgcuKaeQ3VAQSNV7RItn
kd5Hopsf1eb/E3GqQ/ZtwCDUH+Z/AHciAxF9GgHS499WUo445M7OmzZkePApcnEPrRqJ5dCApwWs
OSFL2iSmOAL/Il312ew5GEffUNToi4ICFXhSlZft3h0q7V2AS0UZqYdjTs9oX3yKXs/4cUh5GSe0
sdep34JBo87ylHrb3Qra9A0s6HPTXUJYs3p/J4MH2p4jR+7cRqtg14qqHEfjzoGCAr4xJM8tfwGt
1w9Y36/kUYiOD0eeCO/74NO/7I7sCtBWw9mV0OH2w105/S2mBQq2dPg0/XB5RjSekaFxlaNTKUIq
wYTr1SUA5g3WeVQGUZxyxNp48uJpvJjfCd4/bHs6zp9ZO6oVE3G6A+SUZTGJApDXVYSfgWncUivm
r8inxWqn23Vg6Zi0KqnLWmRn0/kyXYLMp99QG64nI+azl2VIQHVBvybHAA+pUHFevEqb+GVZatcZ
VWsJgxFlPnmKILE0tD7Q651ubOOY5dtt+rObHwExeYet589kEVccg5pVvaIId1tleCIjkMlRzXqP
RMHRQVwjmTYU+CusUMhYVHB/3txOFHKA35e0fsBlL47xq+nzK0ZnwDO8mu15K6WA8d8pzZ49VfLL
4fx4VHVNEjMUb9Gw4fAK7vgsK7sRoAx2aDqCtOJLSldTGEn0+zEgKnoQ4UJalP9mDpQvWNh+CmIJ
2oJbmLbuDcT31iEI5YUy4T7X2Fq/Zja7nokesSdcpA1yfGkbE5CeovOAj95mv9Pb+8zTeXPVu/Qn
UCady9DH8yN4nWIPCNu6cjWYXiRR03U/apgqJ0A7niMRDADJ2NFmWZO6uTsCctZDwKINpXCiZijS
fLWiB8IO52SgO0YSfFYlh9mE7DJMqTzML7jn9uYWWENnl0EyRLk3VeluZZr6MuZrkXR03qSBv59u
xvWhrLgFAOBkhi7pT88OfBwhMsyMvOYSMvS8xXVhmk8bVau0dBoumJxADITU7X6SGa6KJnt78oqi
YCxlk6MZZhpwPJAexKODo9OiwVr7XVr8nXivej3WbT2abS2p6SXo7aYfp1JLIF48nX7NAr9QgXRj
rP9oHgr7YH4mKTIdC8/tbynqV1mHl/OckPt0vLykOwXpA1nwYKZFgb6BIsBLIN+uTOA4a1Pym7DS
XW3/OYbtqHga7ya6hJApgDk+r8h3py2FDC79SzWgEm+UV0cBwAnbnamB7G84Omw0xezp2by/NAJq
H7V0Wmgs25vn0c2FMltSPar1jOJxiIiIvGH4rbv2uG47i6N+vvB0u0qEIv4dL/gYyM6UfPRvYAHy
1kyhhY6iQ6S6WFXtus04bThpper0kEMLOSJedQ4POSa8A+TJqmqeaor5kWwivFqFbiw1jk4PMJvm
+8GRjHCWfZ18/SRCNXs+c/dK0/I/sBSGQVWhEqDP38jhmATb/NRl3r2uXndE0+nH7JKLhF0tbTc7
MqHz1ld2Iy0z7pUh1EunyL+e6sfRZDKR7RyRja2iXV4Lm7CKTvlLCuWux9G2k+F3spjX61eBfI6/
qMFRP+uRMLncjDqkA8PcaNE8T0rdzqV2lY9nrTvSpBhZ0e5Oqi98Ts9EA+LPfoy4EiPHay1w8Xms
JOKpDwyEzAs3Z4/nhXwAH+1gLgnUkCX9vVFL8aVfUx+tSINSP6i6Z5iuL9CTUiysusyafIMgGQ6U
sghiBgJ6VsbIhW/Li9BAczqMi4vBBLNliFBDDRaAbzQAg0gQcx2/POC4B2v5sHZFfcCjFBJ+5OEj
n/kUeIHVxGJ6j2aiBc9MhDeSjYDSZfHqfI3fxaNHORJ5303rhjKB/IGjP/07rQwDrSikg/CotKnz
rinbT77dYB/QsVE+33DCb5Hcbqph/Emj3w5yJv/KV6zAbPFtf8cK8MgyiUdGSd/se2SIFpaOuXzt
h3WmvNYNWJcUNY9QLdsfaKLlPlQiDQD6As6atif4y95vxYQ8YFgiDHJDrrYqhSTQyBG5k+F8KTmf
CdxLacW+xej7qCoL58tyHgH7UN4A2QQYahGHqhtmPJH6BSoK+XY8WCQ0kLiiL0VhM2HMzClrFuAa
ZPzZY+C/2QfWPaTVKX3cS6OtBkBMqIY7YlPp45124EQee9cVPcOgwxSNAjHJX++FMZYXh6c34TmD
uVOWMfbTzYpCcUve4L53iGOKUb+7Jtsdd55Co8i+/0VuWjqNxHSIYWHHsAxK+5TUoqTjnBevxUmC
uGR63o3YsJGvrMLAAl8TU5JAUJVFRm3BTmpMH3Yw0BJfB3onlJgNkn0VgtGeU4v251FeZ2vkrfnH
6BHnjCpJCkwj4k7lNRgiT1foVKqCKh+6YgnEQoXLmJTqPERMqXfSk6EfTym0bJDhrpWt2OzDuDoh
buHBIT5bfQy4nRtB3TX0H59QdImdJWDSmCgs/4ujWG8DpOEfbDxubxOfIUTxL4wpOYuqln7bxv0z
vZrxvT9eYy1hewKOTO+E85mvtCCFVmbRJVMEdQFffwu3Hnp6GiBGhFnpup2wRtb8EHQ/RRVFI9K3
1e8UcG2xbcEOak3EdPrMTHjHcgN0Bk93dH2DMeACYH9jaWly+8jIpksHbapH7iQ6rQdOlzwDNPm6
CXBsgwxqSJojCy5850c95W9wlJ1P247yIgt3oPMsyNhw9XcTK2nERMyouySpxblTt5swaxJAx0AH
lNWtWp/R5CePlJZ2tf8aqkT5n13qvqdtnzm3aZkYelFTIR2APDoD+srOsq+6yD4UsLNRgPB89fee
OeJTOmFRb8VXQ4XpWgZ7Vtx3OFv8rqFKCuV/XpBpr+Oqkk7DiZuPWAenoTDYa6cVBIhFr+2ED4B0
hfNLjaCs6FdR195eJhyIRYxAKzEK386PGpvQoOKexfP9zhz6u7YKd0fSXFBrpWraSnnBlUUakqST
EVj9qQZpDtVijK5OIxHqOspJV4ABA34oVJVEPAkpoGiNlVjBZgTM93+TLBzf1ENzbD/JVwtLf0Bm
h9zXzbo3wmwP3raLpeJHTBRLuRonk+Dcx2t3lI2HDMrM77P5DGZGsIXaQFc59Ysai3sd/1RNFTBH
un55gBHljii+WScnpBb8BTY+zjYNgWpwtOixqP4dqPJjtCWP/h9p5R5/UTQqoEARVUyrtJacKsGb
YfF0fC1C/bEn5hNYOVe2aKWEpDk5GU25ual0qTX9jh/XcavblaU1fwu4QPsB6TZnnWwNmOxTO31e
xcxj//yR78aM49CU5m0xfhS8iyhx7NXPObUYPKopuexm5d7HLTu2nfQQW2gTWkWMM3bGKvrYQwdA
9vY8DoRTPcIKTgsVxxnwos4qUpaEL/o4G2srAsDGNaexCUwJruoJpWyH9G4SHtWWTt0/qzFVQvoN
xN3YoVs2TUskR1boj6DUeBfWWN0ldMSNWrvPKJyowBa41w2cCn99emzTg7cy+TJzE8yW1vMtjl7L
7TYnBAHz8XXx+LgDYKTAwQTkS5zCq+W6QYvHSvgRwkgLKILlWV72rcnavAtYzVhZkjBWd03bPMf1
0utmNvBl9mKdZl+5XBTX+3bLY1iqKM11bgH4kOPU1AmRPKFyYiVbw0L7TdwS21HFpDHnGcybPagi
9vydKTGli2JzOuXaQmXYN2zk8uGrnG9aRjqHn71hyqJWBxCZacukMZtpyEnhD23yxJeegzs0rbVy
9/rl5Ze4q/RsQUZuAJmUfJ+syJ8qyJR3venbLHsvHSRrC/Eh67Y+2Z+e6INryYGta/B0/bLvYjUk
1JAIowWBrgaVayDTmbdoZytLVeVRCxQLap41SXktm/PSqQMj8b42ovPPN22SZRvyUHC4r/9EiWdO
xuB4nsQqppML4FQHAFi7ZluT7WN0RZx7P/HQzVltK6RWUB5Cn4vK7cAhFPJMf2+Y0xAxycNtxWWC
3sOtmL+vp/PGEsJ6wC0gCfrJ+LBvqf2HqM/JVENkJIgQ9OnMs5kEfB9eVedFvFmlQWHi6DOO+Ikh
LfypO6ncTdVF/PYcdrVHYfRddzo2YlgduO7TgSjor8EA7njcDQaMr8NxJo8N5p5tipbngOi6wa+H
l5YKGu/Yzv5JtQJCAkTWSpivh2uNCVPEwCYoldpMufo2Q4Ht03j/QPoNmYPhSuWxzb6XjnVkR8CB
MDzGK7o1JaGlEJeRbOQWE0O6altNY93fo0lj4G34PnQykDZao8lUGn6vlpObrr73gmHbBnK0RET2
0qVSnBLZrq1a8ikcyAS37qFUX2cc4fmVmUvVGimyri8oQA0YmRZWAxArqTL3lFf9xADIOnD8L6P4
pZ2g7adqX3ZDqLjquCOuPSOUC2Ed+6dmWKkLMvEfvZBsPcaMtZEtv2QlPpdbNrbF87Jju43OewhM
qy78Mtw0U2qcZGQtCKJQrtoqyxbhjWgDMa0MHi2JW1IY98mHvTEbkeoLW8R1aV85iNjmVdAW5eJa
nt5FvPIvdroulMEAqlo7QUEA+aIcTVapnAXxlDkRin3CHfL0fZ/CNCApvXKczXPsJvYN+g8iYcW8
KU4LNIecOv8/tL4YI1V8hQvY66TciT+WrOnkzL8XAVu4Dp7UJQE2z2Odll9wGn9LiupssuZtnUx6
a/vmoWhv2sx3/0+DoXmrM12vfyaXcGL5YxzcuY/Gg+Rx7ecuyIa39hc95nHrw0a8vyv/2/x8DPmm
cW3ZnAVWzKpGXC8ZtA/hFO0gFyaUVQbNoqSrDGMoM3Gs0NA2dxNxZizTtKPblfYvkkJeCQ6jILfb
zNVSfZ8G+35kG9BbtKg3dZvlN940HVK53KqVNtq3rCLfhYCLkr6OPRKvd0ITGx4wQih62p1dQTMH
K60+49lpQfMaccYlu0iXHUg5caMToNBj4gwkuU9DNzChCQrIKUsUvErhebJxAnIbTjRcKKocUJA6
1CRcZIjNIo4SS707z7BYdZZl6yT/VkMLxpQvO5DnV/xrUspshChbIYY2oeT+qk332sb3+gYnpzAo
PJ0oeWlCiQD/hD3umbV+mEagSA04fz0A/NQMOSpOZSbjv926r5FCZD1M+bw1+KcERP/kOzkR3e5l
iZSB0zk5+nSHUHNnPi6X50H63eA3gM1E67L5vsl3OkEeWKt/VM7ss/S6hERnQC5se0zAqdWvyQUI
z3q5MmeJf+rt8PfW6aTQGew0oUFhrlLGjTgdo/Dr5CLJtuY1PZn6wiYsPx/Eo3k3i2pHQ2v2qwJY
GscrK+caRjiuPDDdZG+yWL32Lny7dpsaSYjwLnO6emeo4X0qaRUTKan+/ulhV8mXiMwZgvj1NlTj
hLqtfeshleMt2u8vlKsJllrRevXM+Jkrd8zxfCK5MMPdQgLnXcGBfrWs6n8Wf+aT/wc5XkfKnvN/
CixGXt+763ezTaQj+WW1aRA7jknefIWZ5M9x14bt/sJ8y0EVv0oSktc+ydorM9mW8k/GFsqj3Z+l
RB/fNStzU/wLZD7QELzwPJw3kTT6Ncuo8qG3Y8NTmKUfBHROasRO/c3Hwm4Y7G+p2LZErTyl2c+/
t41SAqU43g1yFY1wdG+VG6I099NmV2yawxx7zNvYZ+wfKkYXOSnT28OaTgb943kAwpr+Z7+eEDhy
UyLcrU8ntv90heMoDa86Vserc8/1L25WXYj+B95NmMEpvZHDZ8YQ//CSbZ8i/rtAaaGfNW5MJ7HF
AWBLwCz8lb0wyG9hiXHPyShRyWFO9i92EXDgYrwH1inziu7xa3I3xRDeb845EgVlW1+k7BnZ6I6a
BosKNMzjKnWTHvI8mFb6HIcETB/qw0KvLgOVTwPC2WOQ+pILvoOQ0MLjX+LKlv5EdaZwDXeX4+12
lqhcZDqCy3oymfr+3NWbSm5mmjkP0lq0kVjbRPUEH9hQdqZ2On3MLiX9OfpNGq4f8S1FwkUr8xdv
1M6zXCK0s6BWkI0t3oXxAEwrAS1S6aDr5kbMXR7CEpdf/YtjcWTbucTjL8B0s0HfndYhRy+du8Gn
BtAzoPfwtkFflTFT6bJuCmRxWa71FvwdP2HszqowWpZI69taI2xilHuNyz+LughsK8xbO5uylE9K
xfq31y3kiu5hxXwMgGcOc4Wytq4tMjpjzIi1/Pl93ctJ6Xxbfih2ag/tZGMHoQHl6Niy3VRjGm8/
ZS6DVVgrbnUJU3SFjA8UCRiHcThQhiCM1q9+V7/680hrXW5U4geysbrrVs+fhzgWOOalakdL2nwa
CuuzujAxajQDaf+lF/no8JPug+Uj6e3LiZtJ2mkF3cRQl1jnovJOZuJPYX4O88eKfb0nPTXsPb5a
vBfMdnTJSxB271xGsUfntYeXR7kh4gdIIRYzhjVTzOrzixLpe24RdVQecrb4hftQKSLJooGG6L/8
r9N2HCZEcLJXl9xYnRCvt4641zf7y6OvSlk6N4zF4ajHulJS1eG5upYVYq6e4BemnkrY1EzjKpu2
BKnGHDCanIJSmXex9NSW7YrHLS7ksPITDvEuXmpTPuojU/Kq2TV3Gfv/CaOJKtL/xC8tqiNAFlMO
apQ4ryN/x2U8KaBg4ZZ6EdmaRIldZrkqlVHjXa9QChlOrX21q2eF/rVrlVenY1P2umga1Ex14q3M
vuY2Kghyr6BYwTdSLNUdBr/N4k+DnnwROYXkyu1jSON1hcJoP9Wk6tAb8nLWqJoXE0zvDPs6EDAU
NQ85zL4ovpRyDIf2DHgdpFtuEEqw+LKq06qi0j8jGu0RZ5ONAMzRPbDBlutIb815LV/O3EGEcfft
Sob0oSkCfE3mbbWMqt+ggKE+vhVhxjUtLytfkE/7fD5tr4NUIBm38jsMyuNFwK+XH+RiXc88QJdR
X6UPCngZJk2GVaSpbQUI0W1a9AUVt6nOsHCPpSw8mSNI/+PIDwsw0z4X4A/9Op9W+D0vlSGll24H
B994Oay4Pu4Mlq5HWVE3qXy4OKjM/uPX4TFPL90795zV5ustP3kDnQuedtRFuDQIOilrbBfTSdbQ
QzP9jzP0BjPMc6rbOJuKP8LQk8aoRbrj2s9njjD4n24F5FXw5UXq/NgHmqADco9A5bZ2rYVzqq5+
AnFzMES+2e0gYfvXvwFW6BIQ6ECmvsSU2stDwuzdPYUpvZnsIJtwUPznrk0auGPSjhN9/BIepgVY
ivg5u6wT8eVhNSo7V9/k6IwYVoFBlHFuwthufe/zgCfeDDTKxG01emyniCNfndk8vXS5hS2mlbwR
PeDXPzFMJOD4ycUsxMqkPUa7O+rIlQg1c/rXU8GtC/0KvLHmcWBBqMu/B+LzGXbEpjFS5OYas1X6
0d9lnh2seHWAAKldeMdqhw6lY6irkeqFO8dXNR7CxeHl8eJkxpHDfsvvP+JTNNhzS0aYelFidiKw
WPVeHu8k4nELi/mqYY3fvc2TPsp/dW1aamIAMjCqP4V3y+pJUXE5JpvdpqaLNdguRD3OkrIEcpgm
MiJBsPBiKhLPltCRSPkJw7QK9bLzFHi0MuOharR09zgOZ3VuYZtAF60R9GDEGvhGhdCmz4ED0DPp
hq58LLkw6jiI4G9wqJb/nCTs7pqi8yvBwwieNLUJAmnN7+lTBgPEKlWxV/7AxIeS7bKsVZ8rZ+bg
OXXqwSq0+97n3OiSefX2GfnTIvSMvct5Vp+jQLO85fYL8Wd5IGuYVTYeaxzYWp+EmcgBNIaEY+QT
55EkGN9rBC2MkPyeOx0IxVTbaxPScXwJ2u5bkvecxCbmHFCmWZn5b2459jwdWRFP76TsmYQdKois
gwmCylbn29T8UXXN7ykaJpHMJ1l1H8D591/DuBFE20N0MsPfjU2Qc8nyMG383WBZ9C8BRVfPnqi9
DG8aVFRCdK8y4XRdTguvcYMpe30efozzmBNr3LahJWrAj+1p/Y+wOzA7Z1ZFjMNjsmJVv7c0J9Xs
4rvSefs5uZ/8dHtbzfQqESq51UT3mn2BACTwHNbQ+PyKgiLmfappICtYUaASbncUzmeAc0VoaaCF
T6FOvXx3t/rLQJBwftVTW5dVVMQkDvLxj+mxEjUXQ1sdG56mrUevSSQRs+gBh1ONpunkhKD1Utvw
0GOYONPwWgu6uZoAh9wQTNCEAa+jFvXZoDFmA4W+hBBwNleD2/FpMlfGwWmvt8tsKLqtqqDMYF/S
P49V241CInXlpjn8oYqJGGFYcRPOb4ChV5PphgOIac8fnMRPAuOUy1BSkYhEy1Y80NUwlH5c/DwH
W51ii6nH31ASyJtx3LimOWGEsgS3m3MvbMFmA/8eeXZVTggNR7XLM9M5g6BVWK3iRexej6eonCHO
9MCfBCXKOdbZ/svl6iKLBs+FdAB/uyBXims93sjWgsPR0plixIIQ9ut9KNBLItV6zGormVYeiJJ0
mGTHPPi92od1uzELvGvxp37nQ+5PEsJ8k3Zfr3XcGSPSUyjJjTEofhA7ejUhUyYPfFEtMiJy8eJw
R41Fw/VX4vCOBXrxbLQVdzQIbYb4WV4mK1mAl1IrBi5MYJJyjmKHO/sZMVkIiq9BZW8aGUu5mD2g
eDfDnMlwswAWNypgs0s1nj8H/fpEUkCR/BK9tUhv+3wlUFFfbR09FFXZkTlqNx9+mLUQv4SYRA0u
pxkPtf/G12301gUWtfzleNPW5H2VklPILTygoB81KtKT+SZ17DVKqwJT96fJO/+57eLF3lAipTGg
CdXzw8oxdU9uEt7yOOrO09ZUROMe3JiqsLxCIKqVdpNtez4x1NPV5GJAV4PDHPiLqmTXgICEn+4w
ReLRrqUAEtctww9qFisNMt//v4vsfZV8tEnIIT7KwKgFJYdY9pKNWUlbkCGccyO09VyR0oUQJ++M
Y9BztYYvBB2P6DWrLB/3e/8yfrmQCxNnLG9vi05tHoRDSMSg5RdUIXlgn84xegvhHnmeeMnEzTpI
zRW5WBagYBRFA7otmvyKShaPBybki62PXwZPdyhczZQOTpJxU0aVh/tLF1tWuBr4tCBeJKUiaazi
SsInzSdmtqcUY9eNFbLHuWbi4qkZz9MNPkBbzx2JePM5Dy5B5GnDnGPvQyQ0/RZpQyTkvpLgQdJQ
niEJSuZa5cXbP/RJP+pbcTdZ04y59xwCRr2m9tLpTCarHb2Zr4ETXns7L7kXj5039GA0B/OAGcpS
qIqEw2kOipXYNJ/yIghJC3KKa1aRrTJX+ARrgh2UYoZXInVlVKnMPXF5EsVnhc3AEFfWvem+WGac
YPIOhyqo+V+RTRjE1dzWVnPeKMqrx42wSAxBiNo86c1eu9KvUqepu14wlP50SabaVZaiiyNh1ZLE
E4eTENb86m+1J1jKHthepw89d1OgqdgGheMHk+nq72FBcYf6XdDUOs8tai1RJOOGVdgZgGqz7Kf3
RPI+e1N3Y6yidvoIRuKqo4ieRMEiXqwMbkEAPge8RQ9k7w123/NPRN/2jPAnPjQfLPiBH1w5/yW2
iLQGzAFHc7gn77EHv1E760JUdAiq8d/G3Tch2wiGu7R6jGaFDhuWQe5jkqn22P1Day0VvbayVzz3
Q/mFpAx9Tguc8/jNXYzydYiRuBfMOnkQCaFli7rvlCTYvIOwkbn7ei1NlhyAG0oFFGcXW6ydKXYj
sm/P5Qo5r852qxd7jGNjQHBNMD9wHZJ+YxW5sOrKtdJa0lDewSF0epcR/gQgI2D0vEtC6QFhRifM
qqTfbBf0tAHLl2iOiTo6F+nqvAoBurcSsXUJNtC8La8jCJY0Wx/lcn5MtWbbR8JEpDMefuhk8U1x
Plzkkz4xctYWmI43snrf3KNbLTbYZh2yqrLheqcWw3yQd8i+trzgGIgBdkWvfo5DM+ZgP6NNqfTF
rV2qRMP30lcbOxsHF15CDZ3FyAk9AtJ0l4Hf7fbYRkGtnVgdQ4z4T5sJo9z59hqcyB3GXBGtpQ18
bzBy7jKi0AGq1Rf1z40WfUcDj6/yCaUr1ZtwbmyrChPIFBNmoioOT+9JYJa6AufTiEqs9zHsV5NV
KKwBqa9dblujSZlGwsQR8aA9dCZVHr7xDWj94QhqT8INrAMnW5/N1IIO3to+X3hEdrF5uoOIaKlZ
n2uv1Es+LaGStkkUABMHn8GW2bxnVKwAsr5q7+OmTpY1XQMn1EpLobFRo2RVBvTLJrz9hGKLhucg
LIcdGvg2qMzHJZZ9qQG7sCWMymqSuvKNI2Nw6K+b4+SUa0Wne73F+Bp5SHlhem/1TupHfYyP6e9S
hVSs4D/9cuZQ5Qolrg55nYJCawfuLM8AeNccOr6cBVKDJRMDlJCWx4cXJKNCvrrQQznr11EWXmHq
LwbDJrhDqlX3ineDOFnL8zrwxH7LqNf7E2KG9BPf6nXMBt96DyvyxC1leAInRNnkwB7T1FvtBHqU
0RPLQ5NOkJhwvmXWplhuOYwdPTKsTfxAwGHdBPcOfP0KV1E8NbocP0+1G2Ltne7metk1c88v4afK
stEGyZsXnMuhqO6cHT/7NEAW4Llo38FjtjMluDUzE1+oZZMEKDswV3Z6FIHuZfdDEDI9fL7912l6
QOyHRm9cyXtGPGGgAnsKDT3Z0ib8RvseSBhX2rbY28v1vACseDPUYsw0YOo9mhZAETBUZFFJ3uQf
wX5YthZnSBoj3UB2gqRQw4yq6v6yKAevDkxw020KlTMvBZ467eqUXk91+8sK1a3z0M54R7hnVmZX
aE7g1acQOc6VVggIIncEYUtmEhnGrVnkogukM0O+3HUhuCcPIXE+iKJI5k9FqoPUDYR73VYGPCJd
HE7uy3TTDA4xdge3Nly4wR5GDiCVG9CGitNprttC1u2ckHrrIHaCauUt1sIaPxWmRPMdlEZb0eKz
CJ/IJnVXjC2xjVnMMKIEErwCf6PiyfBzLXyye81BDByZOf9quijP1ODYFpEG0B7aorBgm9jNPW+X
o8v/RWvdgLzprn5JpLFKuDarjnJk9XvsD+rBToVpFdm5CKCdqQs9kV55kR7hqtgWLNwSnb9t3yQK
HaDyDKNid6F7KXGxlIOULwT+MLSvm59AV45a1FWcJX0f0A0IE8D33bPMElvMXA54l4AZiaM9NeNu
WfIWpIfbSwOUmgtWhrPD+qITwcltIHxFyjdZ986WQlP5leTUZasiRbNJyMEMP98OlHJwixjD20j0
yj1dX57+TRFoKZzxEhE5wt2NvSEpUjZm/GcFXBLLwbkpRcJfj+vYyLkvoqGAhYUDoEe82Nv9uWRv
7gs/jRmERBFAhN3RFoSaFtzzOlFqnxGfyabIKmjGsHEJk5wxoGZ5lrggnjAWGulS8PV/Pnhvw1w/
ZUPsDMkHhXDHURAWPTFaeK0p/NyyVqveIsd/zk/Z7ObPXxud/GcOME6pw396FSLG0uHiKatWL9kj
mKaGkh1lw1sIqLLPwT0Kvsq7KP44nkx0RkzRHTt6c+whUVR5L6tbcnX+RCsyXN1oTeLrWqIoe+kk
a5dJWScFqEAvhguu1E0HQ1OZFUzIRXXOmv79UX2D/1Dxa++ft3cKfmqO2OEELf12hycAEmZiJJHv
MHg5y8q1H0EdTT9AbbNlm5a0Y+lNh31t+vA1pVh1HqS3i3554QmE5B2F4lIk9rMcKSEpLFRQIyoq
b0va8Crgl2s9ynnesIaJOqiBg4VX0TiNVPlroaPp8dJDglNuZSKBuRiECR5sdg9DsQKdybl4FGZ8
obK6aI77Ndloe9zjMdnpPg2vqJJrSfr4fn3j+WPsBTAoVcWcjWiJq/Opt227hvgY0awVSzCsZEbe
0bjQjOrNUEVuU5T2wdgIF0EwI4Op8TIKU70SHirhAQ2O01KeDcJ31zlbiIos6ncpEt8kvPxnnW1F
SAFyD7g8wHHMmwfbKo+TjnrAx+zvoLcP/lEN615Y7mPB+sYRHIeHxUp6oWolXgh8wB1xy+vch6a7
zD2mTJFjyB0q0bhvDN555CEovAZ38tUSXKCvt+gAKhOOB389W95zgbzeqVx5/VGpVoGIgh85I5id
8iE+XR0HzQczXmBhVAlzAg8DOYHtYqzA68ozRqwqL3xM+H4pft9dXSyG+FDpeYL49EN9zGh+l0LK
HnAW3rgj9IXb5gMPrnIt7X6T5geTHa6Jxztk/j0oMSa5e197T5V39hii4YtZdDOFIAf0IqdqoMSZ
KB8PIZzwqAK8va8CyEpT0tS5IZinwOq1nLx008nhRljWadELh3NAWCxRdb20lwRl72QpPlxSE6xS
foVXKeMM/GsoZeYWoV9UubBz/kmlSVYSPDCoaofplx8HRZBRXXRbXeCDlq5GuHrDH5FhPoYj9Nmm
xFbpDN5rgBrgeZ6iVhE+DG0Nvbg2JVSlVR5TIt3r6LPpBQayDqPSBre8mqPnljgi3ib9CsOZX3kN
/pO4T0N/e2dIItWpFHZED9J1Vsrf18O9a2NSGHjZ/qHDpH5ne2d1+3mB9fOGhgIJQPDMSJjb+Lj3
fKs8Z4y8RZaJARTTqNV9HZNr1UzcgpNnoK3CfHt4EJBJKFgJoc3Ftf2zwtrc3ZqYumTpH0Z/HeeL
G55VbpHu/738aDfg6XaajZKARlMi/UVicElDJ1j77kvTra8usVQEJUJYYuND9LWNR0Y4vInli9sU
oqIAHaIBlh81VpRtdri4zQG2ZQq2tch10EFKZU1N97Gt7863X9gELGGdVMB6i1asZ/2SR77TINpY
PYpMywhzNFVMHGqenhADjyA5AA4bs8nssKOG7T89/d6jhkw6QkMllVZlAjEAO16vpccNCf4Vqafg
8DHvqr/kFpT6VBheOuia3zRdv5YxyzVni4v7Ro6ixVvpbIoN/JzX5FT61b+77IwquvDEsvwtkwXf
zXIKATULDf6clRxdDZybIfhNJp2xF/90WSESGve96FvHu4m9ooUEdbyHxAHUNmLaL2dJ3H9KTKMo
eHOPGtSdHT5cfEz1wVPBUwPnr8rAU11eo+sUPGceUHXQExEs+QYcpvuzwkfpLo1HkaM80Ltn/cHb
pLOzo4Y9qIRvYRuxUA64lnKRvt1zSRelP3z1C2qCa0b/mlhuD5QD3X5gd7bvBa1o8Im9p+Z0FhRw
e65MLiyt3LT2teRD0Oia6OENPDdjGoAdU0tCe5bXcOcTumwiJlYtKf9MTvMVp050H9TIHKIqTVr6
3Qb4TqBMAsb4am4LH1WHV4aPP5VgBPBGDQ5Sa5BNPApiwAJjAzUbXzNJ2+vdKzesFxbKP7FH9Zos
oxZ3zz38o0Pn76F/ho+RXqkjiFEFczMdJodcCr0FOAAWWvbDCjGP+TalO3mLDHSCs8DUt/vNCNrc
07QVL4ASvho10PRXq5WWqn59OfyS4qMP3nk5+jSsTEFd0zcGpOIbwQcDu6DaGmjCmMr01gUuc9Aq
jU+77njpkbytBSryhrPcFSHIzNIM9viBMu+9gYVYqm60JWjbvICM4dW+Qe4AOKUYAWXsBzsWXgtl
zh9R9yjLdYOLZ/d7LFEeWffiXrGB1ZbIQk0/xHSkChEoZZTaKb6h7XN0E9lu72bkK60oNYM0rles
l1a1r3vdCQIl1+OO+2TWqzk7w3m2549Ndfo5zIesuHdlzoAFtYswKFzMZtTpRtsAk+RoAi7h17f5
ORsECjNIanvXe/XCy119CcdWFmUMPy2b+sxenvXYBvqWD8daCm6Gph26y6ZSj/b1fCL/QjQqlhnO
XYSJyKA468TMiKpYBDFjAWV5pA0ov+5DUjbkRL7fjY/HW+qkogc9p85H9r9ljs1OnwvSwyQwPyBY
bV6vQ3hHr73Ul1Nlx5xYwvc4pOGy9j5Jyzcm5ct1p+GLMQtd5QWaDN53x/c2CwLTlZ/t8uC9XTal
acBWMWC6/r/IHq0KjTKe5jd2s0jhOcUqcoccWw12m87ohO3RvJQmhHU90l7MYHdOXamhN0ZCTVom
KItOka7/XI25sOdKFfgV0f6xofUbY5zO9wvk6J9UcXnPYBojV74HNd0YtjVsFn/9TQeDCYXd2JAp
ivisf1oLGnfMTx5kM3JacQbumrLf58H6NJ9C9juNrKx1STfnftV5jborgm6IguUr/ZT49zAxktg9
I/WAThVZyJd1OICK+9ltUExI/IibbhaOGsymMkz4I5iIeYxyk1SCEtpght4tEQW0V8SJ/DgMXVyM
pFn5yPhEw+BHiQWRenb2tHPENXz6S3Wn6TWlBs+TQgMBUfPz98ePsTtSXvgiVdcMhGObOmnlyNtp
lwIcTyfEyun5/OJ4irdKwU4c2poknNUQ5AAa6ylmJstF0Z7+1cfIeS2HZyY3S5KkWW0mmdxyFQ84
WljQ3tOvtt0vJYV87Ztxx12uyZbffFJLjbrXASXPSrSXmAV8FGghTq2hyToOF/Vwdr4NszSZpDfy
JFV3ddb1HGA5V/TH55V2846CupPddTvjoY9HcZv8BABVoFGDdNgx594XxDlT5VT5BFJk2jUmtwu9
g09AZJ/SFIHxlE+ZwEd24XpnvaR1/UgP0MOqDCK8MgY0gjf5cax58LjcxnzpnF4K6lq9jDO/edzM
OxjMbZ+oA4MnFK50LTlO3JXTJppU8kBccrCJ+cu176dOrOvzQyyt9vVaPqzw0MYhLYyfWOv0J0l5
Dk9AFWZFrAw9CS/JjdQ1f/fNaqDhiMLNSk1nptAJ+PnZgcI2USpbpSaw9ZVnQbJ9f7LGUhTJUXOW
iudUegEpmoPieUQVLbmdo8fxvjLtVj2bNMHdfjdFU8dWTTj9BUD1PNPFNbS4mVCZEaFTLkblW+y2
TQ3CHnsbgimqL/CURxl2r2KGJhMQD16FkgExDjA6qhYBovkyrjp4jmY4eBdN5ndHmuOzoZtZPHep
icS1Y6SXN8JfuiOJPmvuOesBc9KBHf7JkUwsv+inbcvZsB2zOEZuFIFbfs8gT1gBOWU1PqCuGUT6
dKYR++ItvzOKCTJTcgFq9vlpTRmdbgEXqkzSGe9GmjoWu5BdkrASqbS8OB+J4QAA2dG+0HdMMf4r
NF5pilcaKJ8qLhpqxpJ0M1D719Js56ghHnT97g8VIqPC/wZMylf0mFRd5ZNF4af5KoJzc56EIMYK
HFT+zjnXLHm05WxuRA+NHn1ntS704SXM8O+aiTBf3kAFHL3WR4e6Go0ENXfuRpxBDjwNuPIUgMn2
wt/+3IqB6+hrMotzKssER+G7tzVyNg7l5fhPgYtJTVi2JKyQQWHbJmmWVpQRKypawqJBVFJpNh9V
UMIMyUhePv4zfCHePv00Xthb/jUlCOCMp9iMCpvPcBCBxQnUFNG43KeXgmhMdMi5xyXAmTumMfG+
YBL4M1HEEmlFRLVbXB5iwb8ov8sVAG5WK2JD2ro4c8Wla8vUfDL2I/1dtiLyGdlGJPGOs3+vsJUy
7sPXIECp2rP5WZ4xKprrLaSZExOcSLEpVlRqnJynXG9kwgyrwkp94PA2zqG7SannSPsAxvNAYW07
jNpyfXkTH4hGOwr4VjyV27PLZgTBZPhPU8xJ/d+ACLA3wMnwdpJ0Hr7q8LqOEOja01+OpujgMrcZ
anolQ+pYYcc3ffAbC+tZhRVIjAj5r6PsRHdCeSmELSPRU+xPPsKEhMdNmgQ8KQk3kbiQszZH3dIa
fq8L41Fs/0qsyazYeOvh8ir+f1EZDe9Ap04nDHynifsHpG11P8064h803elbj1hMFOmzI3oyKMXX
HQ21RKacTO24izyrhvyLZ54W89ycJ6x5MZydbga2yhaE+toDcp5j4BRom9NIjaY4VRnGeo5vBmNc
CFB5wMLCCxFkdLCwyzL9C3bkFPUBHknzmFT8DYOBiitn22fVhlw32gmJ9or2euhgQlwUf+0M3IwQ
iK61bIW5X/LybakOukk0zqT7bowY4EqcK2A4g75BYGVTn74sGena/5YSDQKLJe3OaY4SMw0UHCLL
sYEsFfdxckXXWOeJ2+0a9DgQsg/tCSSpcWAs6+X9XNcP/3KILOuKXSeEyqjRPkWP1V/Y9Wo0OOwv
y1q3nBmChPogt7CjgL1msC8VKYnFtW9ffOFuQoRwxNBjFUbhvNI7/3IjpN3xnPdqhN7ENwO2d5/b
bFbMEe+PtAG/tXHimhN0Q0TxOeUpGG3Q2tlGagbc1/Hml0f6QwZgO92NT27XSjH1gJqdkvsSonKK
YCBRQBTw68oQvO9JppXy0kaS+HHMOK4GnbnQyzoWjQf3X2jsLRAvmti4hgzb93bS3UEcD+72zEX6
1S0CzCHMd92KSj/oDCFnHCLH2yQtwtlneUR8vZ5nHKcE2+WlSBz2MeXGA1EISyM8Nd3zXutE7HGJ
pIdCJuMTf5fwYQNY+mHACboNoyTUwzdvDn1yRi857wTAMVCFq4L8L6FhIHy7WbpLawmrBewuwT4+
VpxbojquDnIuNXOser+Pt9maovkbhWsEKquQVcpawnnTPJFCsakR37YutpX6uu/027lNbs9pZuyk
TlXZHkAcepsUOUIoBgzBS8qhIySsWnJd95LfCJNWupC7RfUu/qxC8mw+aa/7gf/YqP5fsfPbuMRi
slnU94Y9j82DJ9dtkCpvIEpd0cn4UUobQbYCYLRmFmwahsE7HV+iRxIdb04ZS3Hcch5iCzuh/O0p
8Ilc1cDOZSD1EstNjaGV6RhRL4Q9Y71ea9pt11Ixz+LCTuxulAbrsp11iqRiavbKNw7VDbjHJ3kR
EnBuccrK6Yq42h4Btma3nEYLbVgyMt6VKnsKhw2sXKeRiL9eQqKpjJ7AQFpU3C2EoTZK0zYh5DIH
6mm0ScWZ3FNrmkpe754I6BIzvvo31ekkKQVoKGwsubLbw8tgZWycOLiv4QY9ba2v+Nr9df4Pe5H8
UYq/S9+TT0kN3tgg+MjsFZq6kfD3alrNT552+HP03yoHY4zwAsWV3s0Wp7m3WEopNwkmIrso/YJk
4xLmxe7KC3CMdwkmDAvof4Bz0TgSomnXs0gZDgpKLQnhylXif7w8IOZ+1/p9SCupDKlbPk3FM/uL
5L1zSFIDfWOMJYj1b0nwqp5OQbTJexTSLY9jqmAkREVMcckpK+zyKq1/TI+srlVKdZzB9j36HDri
Z57ghUkw9UjonQsFDn0wsnfuKHD9W/O4utw8i3f9MIcOExov91JDgAxYjekQbXHw1TuZ76NNdoaw
H/lBp8lq6ZaSr3L28lAaOjtOJqGDDHcklzRu+QXAvgy6ak6o3+8+F5ZN26wu963NdHGufUs7Wr4l
HaHn90bc9ImAN/6VfCsgymMSfjTJha3r/FIYYZq/eeNGcpESo/g1QM4fsTR3Y+L62y6HMHNiJPS0
1Uk3bAoywNaDTWJMTpSd6OLHqUVGP4sMpwzJ1e+adIvA3cMf4cjZa1+HXUcYSs8ZmKi3SBiAepix
lXdKPn9JJwrPPf204ddFS+R9TF+M9UPTuLzHGBZGQ6BXJKjg7I88ikFA76UoVsNJtr1Kxqog/Gw8
wdQ0KsJBrq6qMiR9gbmyIDvM3t6GsW+I9TgDai9v2tPwTP2iAbh9//Oi31DVeFKOlKha+MF0eUew
CB/p24qqIvMc5hwaEMfHbns3bU2ou6zURaqR3GkFIB9M5dSfsZV/oUSiZfgVhTzw2UaCSznm/hEk
kycAHWDtKGeT2Fh0MqtfIwPmcN8Y/LBkBAB1dJZI8jkhG7TNoK96WU/CO3w/Ef7YgHndnXUgpmc2
PCgs0LBoXbGhhFoYpPVU/qqsaa3losKrS/tsh6/r81KzJAFnrvT+jHbyB+wZwf9ySEPIPwPK+wao
hG2blm2sMQK9RSDD5SxZLtcoXWFUe2pLXWbB1qDYdxbEQTHKddqiY3l/ejjyzA5oYO15YdLOZIpS
TJ2aMwSvYeN32ao4yTgJhU1lCbdwolROgM4WjEOL2pVkEi3JLFl5t0528/J4p92lo+swDXm5qtK/
o3AsXtCBhtgwSZjVNbhx8no1bQdwk495ZGM+WmxdbhiJOXbWUosSePWneRQkcYqBoimR06v2tOpj
mF+YNEaJE9tLC9P8te9JK6M53n1nb4snyZzVHF51RwAskHV7UaifZXiB90FVr7UCYAxHUkT+OhM2
PPKLVrF0cuZwX3yN/n5AFIAWSUBABQ8FQyNY2diQlI9rdWy4N3U7nCMhWOyZNenNOPa5sfCB2y1L
Q32WH2ofGps9iloRaw2d3vlghET+3s+mRnZfytraF/a1WZXuNtCEEAzJ8gU3aEJjljOMMxhJhw9/
meVZfS0quVTpBoMT4QBcWiy1BvP9QTm0vxMbofBa2VBihAYey9joFWp69gBdvfVXBR4U4uVjkNwc
IlUd9KbRiZPY3Ug18kvOonvnC+R4lr9pu72ZdEiPHs/LqfW58NDeXK798FhKnprn/Fw7n2aYtKyA
YVmYsFDPeEenBPYNg/OSuYsCJBzcvfvsVKXsqM357ZrOmj9fjU3wD0IeiuTB2BH+5yPhENLeSfQU
oXHRDXdxAxQ6F/ONDQha9DTMN0n10Jb0g8FTshlPjHpYt1A1pe2wzSTrILoKGJnp7Mgmu2tGH9SQ
gx2kKneHXT4fTxhPF9H3IZT8byFXYf+WNp9uutboQNjnsVM35KxE4bTRniKpTQUiwqufOc5xgKLF
gYPHFdrf+6OMEjt9aswKuyBLSVAzBvL3zUohSzX4CoWnoEPCFiRt4ppLcuvXlVjF4CSAbF+HGVNS
NBxDfL1l0bbzSUh5PUqwniulk8XfaKDoHwFOgVMgzHmul3bIJ9pSMcNsPe25Rb3QVXUsaLI/o1h6
t411BsJHh+KhxNvGV3MZCXak/Mn3tRQZjuOsEPqMCNvtkKGqSUDWECNExPLrfcw6veknONBsAjkb
faKC5coBtm2lIc/UNnOQKPeD15TmWeZdvTGDNJ0x7T3eCV/cf9iptN4HXd9HRDHXrclKpnnkMiDg
hUZKqGqd7yzkKKkgIFIevcU6kuwHeMeq4KrtwP0n3XGpqnY55GxEXqLP4HGWWmm9XtHkW65rJ7VT
GAqos9qukeQzSSOdNp1gleyxf4tz0VGaf7cQcfpSqipLOVCFkpYQDAFohuajc6oIhPvhEpz4yv8S
U3netotTAmItTXYQeIrMOPpCbBjdqV85cqmTox2yio4CgN1ouWGoRjS5w9S6JrcrFXtJ4GLo0abk
V+YRuWNJ+LgXn9yne8mLcMs8S4xjudSvuP6omvg14GQrHmy8Gr/5lrwweysLjxT0qm4i6EgXX+6v
RaK0AQ2d0EnApQjsF06PIWf0K1aoSAtp02m9ST0LpuYvQu2965MV/7dVG6ze2oJtp601+j9jwogA
uaKSIKL3Q0fxHHmER+KHOzNWyGx7uJuiwgThBujtyA0m/WFU0ImftWXfPvzfZKlMcNI73fmFdwQu
1JWmx4jWOgqIPoFCiOhNTPxutX18xgH+A7S1C2Nasj6IB4EPBuFO4F8LBGgw/btgbNMDhFRfC5ES
lrpHec8Y3vpRHIFiu0vvO+02ZsPX9Q/jgp03SPNxvp21LGrurYLIjzlZa2OIFxMFRxlqfs1/AxW0
HH0cU4WklpcEOBuFhG9xKRcJ0LmuI7UCiy1dQlBUHoTSWar+ToblmvwTuNXn3xkqJ7k2cwR85THX
0qXWqKBUKDa9hkWMtoC02o/w5WvJR9zMPYXnQNTAwutfqaigYvsh8R+WbQ1icP3pckmcDhA3RzO3
TIQB2+xK0qySJxazd3PCkHoJHUMhHoidQI0nudElaffg4EppipGyhE2rdRx+6fGsGXUBY1ppb+Gc
zlN0Qmew3yISUM3lMFE5Qt+JuYc9b+NbQqg0ZuAUuQRdgZSyrhSWKAcIjPaczIss4vCPL4Yzvd7P
c6ktSJrLgFcA4SdufODInM1bKu6TrU+nEeYoPAq3DepTPY/ZHgOKKrKs4TOmXJc8b8YiBOxRHg00
SwoXwmIAGC7vsOSMU1D8dAyyfzHhGolPMayJLAdjvdPI5W8KiAJ3nWkVo/LBzXNnTgBLj7rGBUSg
ynuRsKGT+ycLoseZLdraFbNlb4nLXuZM1L2rD9HOD4+mbklYhA0V4pd8b7YyjJnz6mW9LAaYuib3
1Zkd5v/g32l7mwVGsmzbqtwVAx00RpRTt1PjvxQLSNqvAzwCEc9z2qeG7JhbP57ERdMMRXoN8WtP
LPJ8FJSkxOP6m9mFHBWA4nrTuafBNyOKcfyligw7VkSxNS+7n6tm2OAlwdS00fBAKWIT0uLY+Ssb
yoslgMWr66AbjYfHOfEZoevnRmY7GjAGdHSS2HdbUmane0aifGAfesoo88yl17dLUlxClyrKvNeU
81O4v9DS8wp/RDPkRk3mffwVRCieE6UoxzMZNHGb4HoUT6Cs1pUY8yG9qubsiPO9mxWRk0Ulac1A
+A6eiO9dzIh0nSVVjx4ZI47u74Y5z6hsEpB1o3FevflGbhYmmmsFlPuZPj/KnTrzLQKNcpnMK3JV
qd/nEIoJ8QIQORFZMteRBLj3Cetqb7Y3EonVod2WuZlkMq1NKtM2OlobX69jiviVqJn6oVAgWaME
LXIaxn55GQgvbCzEwzupC1EfQ5DQz2EH8UtomrvAS62JiteocNiobwvMNTl0qFYbi35414ZkRBt8
ghmN0hFiVqlPiX21/VxXPZ9BqtgwtThAMqfAUmVfrs5/VEi5pvS9Z+6M7clwBNDD8JA9mSpd24du
vdwND+jdxi0tzEOD6d/aN8SIZWOX9FvdFi7jtDQDFiKC1l20iVUi0DZ1wgTxE82xPyWVTUFpOjQB
PgdIPu/xOoRLNXyF1/tHsQzqJBN8LmPxBQ9GKcTkjWPJSkjMDM6g6MQh6tKaqLCI98cKPUdW3u/d
ON+e6I5eSHK9Kzr3Y/ToCOnqSa+bL27mnPo8YbGmqb2bMsDcS4NQfa0tHdND1Rs/DPcxbbRRnKaZ
V/XA+GtrnxLFyx54bRPMXX9usp+21ib7z8nqDJIhY0uwl5twUG0v9raIufwy6kCk/XtB0y0Qu3xk
3KmffIb/xBj2aYPNmTdpTdo2uXKaRhtOuyD2mEfT0Wpb1OxPtN8zfYCZuSbC2dF3UJ9v/7q++BCB
EKeUi9nVhjRmlVD3pPQxGw3Q3GA0zBAMNRlfG9BLoleNmdrblPOAZ28zm65AI3bX45xSxZt3/f9V
mzh6JAegGyqhRDWka/CKnAeBovaTTJOLerM2PNGgPQ0J1n0AW7lAj3s4GBmnodc7YzWWJOND1Ru2
QUsgV7s8navZdabuYUN913VkWZftL21Whg0ea34dIyVEQZyx2PgSuBX+ZdyB2Y7WGPjzJEcvz67f
VdX+XkRIN89wfqF0CHFKmjxsByB4Lmue+BBoaxg8x7eann+qI35XXZrMPh6bpo42t2nxN0zgwwVf
n+36RxTq9LOjBe4+TR01fKTEyOFgg9qR4Mer0GpNvbExOpTQ+XD63pCUjXsfCrT99iUjllv/BTle
MMmfkyJ12rYkD9X/Utw3F3X6f7bTytrqEOZhhHi85UgjHoD8oVq+j/99x3rUQQvgzSluhM7Jzp5h
8KOFRJhy/qMMTd1Z+DgigJKfpppfgk9jBheuEW8zcVsZctejySOtJZHiIvC+bRDzZYMp8r75kCnB
vqGOyRJAu2+Rxjvt+OyVNfEDdkrSAlbatt4+8y51/a1PC/7LMA/VbXIeEIl0aU/NBwmQMk14djkY
QCJmjI6FbunLqkvn8lryAWjfwrv7nOFLL25yOlx7NhwAkyI6mIjGGYlW/V+g1OCb/96IDLwF3P54
ptxGbcReGHkTHtQ74oJUgdQ0ePk5qynkpiDhVTrHp27F2Ulzk76F+6MioEnIOTlNaigktUOr/lUW
GkPjIECppD72AV9trlFT0otnHmpDNT5kFbMW5uDu9tkjBGEGx9NcDWUYbZL68oWra1Hj6dtNQtgo
lu1D80ndbIUAsuQhQMnT2MQkZUgAD5IqSq8t06zLO5kYUkhLSaBYBe5YFUXvaB/oiu1oDIrApYuI
oJcN6IKH4WbDU3Bzj6AmtpPP29uR4fV7raOCjEISKCawdZFzZ2lP0jxWosHzxFc7a9ondudIYdKU
E8wbdGncYnn03J+jzRZwFB6mPd6Kmc9t5esT3fPsdhhNn28hvqAMS877MYYAC/ac/CDKKVCPZwqi
TGlcYLBpue+lW5XGlweMALFKK1kO8DoBmxqPzp0XyDOKrq5mU6ilwh2UoxSOXDxgyiRI9YJopAsb
5hcVm8OYFwNphgZAo6MfT88rJzXcanTXUcAn1P8Kwv9v3dMDg9CVcZ8aRV72gSw/EuFEwqVw0OK9
XgpUEwoSFauE5W1yaMNk30MtzsfVcwhYQdxgTSh/Clnkok2tp/KLgqzwGEI00vekvqUulpnQJ0Za
jHjhcrjsvEH2XXSOMiM0J5aIAqRETvGOK8sIkRka1SJpIXBgCBs9OIeBYgDI6OMVTkzkbU2ZnwP1
6p9FbKRf6JoDeJHi5vIT1kiW/l5GgvxmqrJedgF6G0AQVVtvEEeEZuVSMatKzPOkQ3uDZv1Ihpvj
CRfrkf6ebM8IR6Vh2Vk5oyqNlCy77OL4na1R9G63ind0BgCYC8lk9zGlPSr+uDtW/1jrkGYzp19N
GE/MunsvKD67JYylBFWh3iLHPYQU4AvNwflj72uCdqZAp8XVc5CDvWdI7rJ0s41Jwu0gILz+K5a8
OmW5v2rRPYeDh8yagyqF/Z4dP9GGoQyrybdU8HCSJk1FCAaEAJpbK7IVyO+REHPtceHn2028/Z0L
jdW23naP0WHTori1DTMa8oPBj49l8TSC9rdHkMUCdopvvryHk87JsY1UQhYH8AJn6LIs45vWHnEn
YLKHLb8q2mIMCsQpocNDacDZUtUzBa3LULTXUQw4Vjas3eo4OdAV/qSYFHpylAgGTvo1BcdL6zw8
B9pz/iazxuMC7WmTE9j+Z194lQnZL6dbtz+isQNKa99KjTxF9cHV0kOsy320FD4PRcZZu4QHpZLI
waiu25ZTwGb9NTKZmWbLQawkgKwJFrhIzncN+UuyelEZrok61ZdWjvoDgr6AzEI7FF5n8eS5fJPU
gvPqsPofoOwa/nuKA/uZrvsBY1qP8KKDpd4hE0b2sLiZWzzyfGbh9P19hco0mEwlP+BDPW21/z8n
lmVm8YpTBd9YoVzsDgzRQY3kg0R4hUrpQNS2QBLkb3oyZy5U23RT17dsUtU2AyP1H6heCWBU2HWj
+ErnIaRw8+eh4faxD2XtzhqboLNpBZW/aXzoR7/sVA4BCj71qhPZJyUoadhprUZ4VlI4dwBNYJBr
DdGL1qQ9fWLc36GvBAMpWJ+5psbFIIhcRe7uZtrcIAxAd6iwArmv/Ht6C3TsSC2GcvGbxFnqb9PV
Lvq10PORC+Tojmq5yjcdPNfKmpvq4k3sJ0d5TXwhxweeRPtloSaiDe6ujB2o+OQp6U8KkfVnCl2z
lp/3ThsL3VXPWuv2JP6JtOxik4MFMy05VneLRdc3MmfHC0/8oAP5YyMUXGH/n1WDh4KaFIKoNFnC
CxZco+VCb+JPJnfxmBMXw3HTNi2XVw6Wcf1qFLEx9p1eJ+hWuvW0K876/+Yk2fU+twZkY5t5Lt8R
pZ8I6seHPLSf3to58IQNxNSh9vTr1XrioPCBdgbLews3/JQdP4eXx71MqPQqeyvH9FE3dFL9ZI56
G1ueZKuVzqm+jASJ+fTmlf9ExdSvIyYcclA99DJIsDUGnBDXY8qgPWqohooZL6LJyHMxhn/xpEJX
9UV8su+m2seTTEuo9O95yXryVZ80h3LyNRXJyL4+q8ifqtFwYoSnEJSG5GavPpNyYE+J3uaJe7zM
GfkrkrU0Vt6OYbeYUHLv6DwgxnGGhLY27Kwisy5xL5T9+JqqJDCJKSuZZT9EuDLz2VE9c4THnkLy
akNmpfzXeZtihgLK783uaPTl9r2sbfKGTDG02u773jD+t9YuXiPpWzupDJDwLzISzZQnCequJioO
zd0rTF8j97Y2jnJyQEcdqY2REsL0b7CEn9fEba1G+0OZc2uzL9DPfpKBYThpVz2CgMqEmEL2f2KL
/wDOPFqWCJZeFwLM1gEOHXRAcd4sRfTqXM1TwdItalRYQYQ/HFITtoynk93Q6UmNR6IRRlUvPA5o
/IE8AMhvecEHAabdXaSXUhRpIgAV0kZHuLztIgmtClsu4Q+CHczje4b0tqh7gcUjc+dXfFEHSdk2
pzOtuc29Hw2MNiusI0zpnVqr3kYlPmdhzA1MLA1qOyHM0cVSxbojjUzR1v/ZE+2hHycpnEuIaV/a
BE1vxzCQjZDHmhR2b18hFGlwc+fZXI2+cbjgcDFJqBHw9IyFX7FudHPru9q6Xj94NWHaIdYcDmE+
q/YzLqgeDhVwFfKSvXMdWWxrtPftUquv2a8dynNG7ODpM+v1nN6q/Akop3SQCtf28c8kukk+KFJ5
WweJs/8j/p3e2rHqEL5jxszI3v6mMNeCZzTT7unlAD9XwdF3AYuN4umfsBmAqPl8qGu8ioGTKoy4
J+UCU3BJU9fghyvKzkz/CezaYli05otGwKNCgqdjHNDg1rDxMUUvfScAlVdSKYTW+gXFxX52f7Fk
PIZPXKJLEAeHGvsK2vZfcq2ij4CtnAtXToxwEkGQCgOUzIWSHARTAz99rytW7skWt7eNRMV22INn
/cssfnBIiKpXAj7yEeL2U3+BOqWaVXc6D3XudV8R4U3zo0CfxwK/rK1l64SAeJ0sfRsfB6zewyYZ
1el39K1PHiQOuWdKif5m6FDMgqHt4vxxGdX/NDGIMYAmbBaHluOLXl9GWJJTcP2ybMANmnZW1Iyg
Yq/CxIZJPQXv+0E4WJupnOd1zBTsFlLmKv4rzpd+BILYQB9VBrGcE7TbIEgZa693OqFxw7XKhJjt
PHhxJvS2GNUJdR1tAYttC3XQj8pWkBCom9Zwb/kFIi6isJNX18pG/JVllFsdcm2/o7SdCLt1IiNP
b3fPVehH9VWU+NMgybm45ze1UNy0iRK5J0wMCCamqW6ii456hlBn/fSBkv65aLIVbBZPt8FTaT2h
r24ZdpO6rLMXZC92griKuI9NthgUYl2csOx1JYk26/WeX0QxTx47RGHcbl6k7gdm/h2ZEyvaVJJ/
/+kwU9xFTQRlPPzahqiMGQkk4L6T0q8b3XTx4i+Ab0LbbqAIa/QE9X4DEouFAolaQWpv46+Klnrx
qS8l6SzHU9SAt9VOHtTFjgshOgFYcrmRpONrXdnoggIV/2QOMCEP6ixw96sKItXgofEl9gyQ5NAf
aG1ESe/GAS3dZ+RheS6bWYBFeRu+92eRzjs0Dcz9F9ZAg9p8gLg2xu7S/mto0F6v9BIoW+GuYGXV
fyAYaLRd211/tdnFbLCrhGjscN4W/ceDPmmYlQsCgXAQhNxzFmhHN4gXSG8F00qefgEtdXvEobg0
gi1HH9X2w4fX7CLAyRFCKLsXCrsV7PsAOSEgCdxbjdH8cGJC8eeVA6lZq+kIL5NRMB+PbLuqwsxW
ZCPHvN2dC16c1vIVcecDVsgxEbMYugfukZB12051Qtv/N5xldqELXawPe7oXaonlDPkJFbJxLXw2
FzZInalDhQJCsxtEmxkh2QTK6WlFGqPdPZQaQ7TO60Jxa68lrxGzU+Gwih441dLBpK3IwchkjueJ
zy+1+yAukHNM2rRfjgAtlXzM9YyiIyWS3+BVjML7RpZiR4+dF8Alb3Irzhz3TYGzhgGRFQASY0au
hTDTULlFB2Me0gmc14mmG8ZoLa0iPoKoCl7nhCHrK0YDVG/eZA77xlkWX8j4egQB4y6SDS/U56Nm
NX5iQ+IjpJvWDssWvLHVkNrgYivUILH2vafXwlMAvOhTLq3rrmcjO83glzMFya10YufBq/LJessi
3xyy++yvAzAXFdQuxD62Tjq1eJbyBFbjvV5RqXMqVEcETXfubXcsqbij+QvT3KlCvkNa2s5xJiAC
RmxxxhJ+epYPHjJw+UR5llw2bDfVpDFwOf72OlU4tsvt/SOYcKqDzbIToaoxLVKlTAA=
`pragma protect end_protected
