// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H>0QXC9N-<80P4E4;NS&B1/7D#4T>WRM=XV9J)!_,+XM#T3_?0S"!+P  
HWN.3&N2+9F'DDZ0V1)H4T;C[0_C[;#O_/N&$RH-G)<D;X1$*7# 3 @  
H:F>/0^TXZUO2.KBC["K"/_)/$[TD2G(K!RTR>=MS6GF+J4N-%N=?YP  
HNEQJ#F5LQY,7<5"<$KX\<_Q@\%$IP85;Q\S/BH<[V0O8GHO'/24*B@  
H-Q!BG]-L>XACGT]VHO2K/:1M&*%Z)3AEHHQW 4DW[!\>P0(%>'R46@  
`pragma protect encoding=(enctype="uuencode",bytes=8672        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@*M3;C[GM@T34+^+N5MU<\M]]6Q2TT5ESL]JG%-Y> C\ 
@YKHT11YR<GHIV\?%1O69)7!51OL?I*?1[3/A7EC\"B@ 
@ G@A%#3=-S%2G.9TLL&F(E,6%-$A?\H;SC,'XJ]!C[X 
@\*G/+H1J;R"S-;DXB0_;[,PTZAH2GREK0JFL BX>JTL 
@)UF0BQ%P\.(O5A7;<GT*\UC)B&J7RFS.0^U22NPVM%0 
@>)%;J,Z5Y5;N2FJ6$FT2>>A^6&/5A]X2+ADOUA'M9\$ 
@G\,VM#1OZ)+\\Q-B(-"S9?)(VMD^E+N]H#9F/)E<43( 
@6(N5N4+_DO_ '#G$Z2@;UCN[+O?"CZ^R?6^QICY7>$P 
@.&!SRG.)I+_(T%CT/!U5,<T)\:.ZL\Y@%9?^= F)ZW( 
@-7#N5DH^X73'MWD#W0"*M>?ERC'VIUFAO**]?S$T>:4 
@IGJB5*LFF]/D4*PN_^(G"@QNNWB8@O<10V/'VC$A&@T 
@_FOPC-R%3MG5G*TE2R_7EV Z^_F::P2G YT OSGH=8\ 
@\6)'TA#/$T@XP2M/_T/9$FA)O3$.;ILP!%)IUUS7<F( 
@3ZGKQ#Q(+_83*O&!H9NBHF=SUN-7!GW@.@<&L*I&,:, 
@.2!L?5,WH-W DV6KF,G27;"==TM'H3U!Y,<I$Z .$<( 
@;QT@B'1925&<IWD?&A<G^*:N ]:\T,8/_EH,+O7;I#P 
@FJH26\O@&_PTN/8V7C30+'@/?GP-7K3;1#Z?4?=@^%T 
@*\[I<Z4KI.W"2@L=FM/88YJ'F7>#\<R(-W_K)=QE3J  
@8 Q]3!">LZBD<T5"PBXP%@S5_K6'.Z2C,< >2PRN@YH 
@)?7?[QOYGN H;$'!U@:8=-PS+A%0C3W2EBUWUDUBHHP 
@(>6M45Z5$B&A3WWQ)Z1T-)&R&RGZU"?INJH/2HU7, 0 
@$B:"=#,<UK_A.Y;VA*A.\A<VO%B69;'@BDF[T38W=D( 
@:/-Q\2=2#6]V8O\=XV(]>-H%A)H<1M?/50"T:CHB+!0 
@P> B,'&%>@\DB_//'\.N"C[R:9ZH+CL6P'9DB*2[Y7( 
@^\5HRUJ!4]3YG'0,K6,$/Q;THQ8$WM1!6#7'ALL;K+0 
@/[(6]WR>H*-84TCZ(/9[3PE]!S^]OEB36*^<@X9@3[\ 
@ZE*VY^0W9'<3PW"[XM0_\_>C0<SJG(&3O.)5&B0:F$H 
@&0$!(RSG@>8M4HNQBS?F/KC;0>X!':?.6&/6.+:W:5H 
@UKDDZ,HMR%P>ZKJS*">COH-D1M(LJ%3"]1$/>D/M&'L 
@/%V\N2?\; C^4[-M]0-6CH[DVURI0HGA@<S@0K?BH*8 
@&,C]DF]&W&-,KJ7[!CD!)%+)Q4$=S6].X:^D:>O$YMP 
@"@G@Y!_8_?CS4Y0^:U'#]@4&X?G>;$K,^ '''F>=4#< 
@MO*EM3GJH)>8O3-PI%;<C2A^5+,SU/ <C3]81^ST/]  
@*R"9VXF+_T#LOQ\498Q4-=P,^/<N@V^JWP$;#%=THO0 
@K!$9&V*M,Z205(#3U$*EB$'\,0/)'!4>M<'[\RD2_NX 
@%-PL:[AV/73\/: KM'Q$(+.@GN'_IQ&^QV8@/PD)9R4 
@"J]/8O4S*Y/^8H&?.'IRS*O9X[9ED)FJCU6@$^R$F9\ 
@025[.!/5F[+#-C4KR-C1I=\%AQ*[%V#B",Y\ >,\<M, 
@M)S0!99PAF#?6%E!MI"I(E1 9Q.@Y-(9B:96299G:1P 
@=B%3;#08?V ?5E%T+\B4VE5C=3?_V*FP"L%*F95,^.( 
@FW%?K2/[V72\SZ-)0,"V7+;B'%:F^MPXM'LFW_Z4N4P 
@8AX8_V(=%R4N;AB/9&4+O(X$E^AR$;[.7C_B;O,CQO( 
@O_3V"4+]#=8\RHU#6'FX)5KS?ZHT.U27(?>IX9=>$,  
@&16KF]7E5FE'*\S.>\#XC?#^Z&,!CC'/_>'N4V:.TP0 
@_S,06U,<, D.J$;(N-WL:E!!7>1[L%F7M5R2FX6("D$ 
@\-W8U_NU(<=0.5A;GI_4*8&T\!]CE7Z<+ 1/J:/^GK  
@IM#3/Y88 9N1;C4 K!YG="LRD910&)*T=]GC@?I17QP 
@ZRME_*!G%A*S* ,A$ROS\B19X*S$J_YBR+OF\%G&ZH< 
@&(Q>6[&0 !#,G.JS,<VHYU2O^;)?5;39X>G+CK.4Z5$ 
@6H4V5::.=FI#79>1C\SY(NO%!!"2FW#Y2#1/[7@!D]@ 
@P/?=&QBS&^A6,;-*%H,PVG%GC[-%%%)&O0Y.BJ?HG5T 
@;%I9-D,N$"Q*9/837>,!,2\L+\=D,)?#0/]#D)K:O2P 
@WP=.TU*_BWXWAY>@(AN-5_"C:$=FWC?Z)QMIXX)>.', 
@FDK@L3#_+=>\-T$W\75!TLPI+1NY1QX"HJ%\<'LA:7\ 
@D+VD>MM,:?7(Q^H^RKA8E'()DW8LYA&_=CYE'[)Z,DP 
@!*B!N43OPY\TNRY15185ECIS6Q&SNL$=_9](M[X_!L< 
@?0#)>L>$ UZ44[>*5E+/44L^"*7T6@R1D&N\+_)(<OT 
@,N(B!J^ZN7'/X=\2OV(RO"USW>W5G3!/#O3FTTN6Y[L 
@%E!H\(GP: A*L??X0.0:)_0T) J59',EA^VE<+Z?'XL 
@UA.\8$%[0 P 3<#<-&_ D7W#<L;=D@2=Q6-TK20<J;H 
@^I6!;=<*PY/- K<^CLE M(9X^8PE1L;K0E-BC!Q!G&@ 
@*_R27(N&;2F#D#E0Q;>'O&Q8P*GV&]H:.2W.C]&-)*( 
@?(G OXO.S)N6H&QVO?^FDVO7'JPIY)()C"H$R- 7O:H 
@5K9X_9Z#H.C)]6T-:\^X?$5BKPP1[BK@N3\[52H" >X 
@BE/PF1)&LTQ@5XRK7%BWO[,4GBXXC*Q1P%>\;Y6R-_P 
@OS&X9 0=^B2-Z]9/\0O5)+>[\[/["%)V1^^7=8RL&ZX 
@83U?3^G%T)__M)]M@JT^UI]L +^QX58B_^&0<>Z/\(< 
@!U$8I\#JKUQDR$)H#"_F#*!A?1WYG8$()Z;K1% /5I4 
@=_'][XA.6W72(R(BVA8G4Y@ZX-X>EK]X+)G%:"J(E78 
@AW\^:;[\8&,I#)4%^W8J^<G@AQ6"!G+@^.?=T>Y2>2P 
@$0QW(I!%4;?4=_"&&X%).\",VPDO<QR69<R)Q#N6$4< 
@"P=) @$SS!D[53URV]#KQH!>F$VK-7N5_R90ZA*37K@ 
@V<],G]!"4N)CXU?>>=?/1$)6.@E&8GL, QL.3PRL3DH 
@Q*/T?07>E;JHF"T#G6[>!N]GB(5I+RED1 D(<9R'43$ 
@<6I62KQ41_10;ANKF#" S[-'27C54S*#J)H PT3]*H  
@_>(GRP8%S&0U'&P5'8?/X5#E)LS?\K(6F4$.8QP5#IX 
@$?'(YG &FASF+:^3".X<T$=9HOU(:KVG< XZ"+X;-VX 
@Y7LWQ!]<J.H^YSW0+]=OUXSI_*@>0$NB'V0XC+5)U\$ 
@\^):")105FZT4!;P>],!'--6O@^GS4MS: 3%D(.;O7X 
@-VG"+0R_:VD?S<8+9(H=\)E_7DT]B];_-C2Q\K=9:AD 
@)\7+%Y%'__GKZKO?WP6DQKSUZQ4CS.FY7D%7[XH4/T4 
@5I$5/_C(L#:["TN\?^P%@Q57>67C %?&_MX(C]]QT)( 
@2/8P^?LU%>1J\@Z')"/F/L0L&:?"%8@#@=06>KV])<X 
@/&AW@3G#7BOKMXHM9[4@.4B,^DXSJ3#II7:7RPG_L9L 
@-:7WRBRA?=A&_PIU43T,*9C+N6/(Q@XEC+T0HC37 \< 
@V"-#$R/%6$_F^7M[ _>O3#FNV*-'(,UQ$1^8X[^[A#$ 
@/XT:"'\,]!=1NPPWIPVH._4:&RX(>0L<O\US(,E=2KX 
@4"=@"X;UA*\2P8Q7 :""B6N99.W):Q!WNOY]Q#I57)0 
@=E40FI],-D"EMWD%+^)HOA3_0?;W* N (ETV\;U/K#0 
@#=K)8Q,-#[RO0 WUM@)#U1&9;U:6BSO.1]YBAO!=%XL 
@U2_654"Z,GR&*.OCF_3E]-Q<+EBB(G1H]N'G3.[8 TP 
@SO+6&P>7.<02#Q(WL\I&P9#TQV=:R936B>E:>KGD  8 
@ZOLRRC4%'TTFJ(T[9)3?VUS#F.<3\2I]B/U@&. X>UP 
@V;,'PN]0F9.1@8]#6H!?-NW$OKH[Q59"G,^-8$N5O?X 
@:QFCR F%P7]61R&S!YN!$&@<S%NAYS%H=P@%4LX*()$ 
@RVV>(81XM[<4",=Q36&95$LF'D AP"SYY.'.#H3L*5< 
@N(]F+PJU@+&..:F#)(14RO<JW8\DOV550>JS/H6QR>L 
@!NBR.D1C41>G5?J)TNIQ]&GI8@)^BL=>I=EQ1QJ'.W@ 
@7,<DABB"!JVQX8BQBLB3;1A="C#AD-]%AY#S$XWU+!T 
@%,%1TY+,NS@U_2CY4]2#0@QRZY%O^N/JCWI%7M;ZIP  
@(@+758]X53@Z[J24Y#>A^.FNPXB5UG>/^<+@L ]0YTP 
@P<!(A^;BGI0N0/.SJ3<OY3#[N:C$T\ "SHVQAD+M$:T 
@B_);\NX#)HO1\B0,O+1Y/%LT-?]9R>T3NH4K$GMDTTX 
@T99BN$*1LCGZ_M0#>ANJC'N.4.:Z8R;+A$IP(P?(Z3, 
@$+FYQ%_"SUX3685B;N#A>JWDN]++]+]4%(%/>A3>BJH 
@,&]?.LJEY9FZ^W.;>6XZ?CKTRQG0-MN@S;[1KOC59YD 
@:6,-@,]RXYE\&.4F(WN$_1CV2,BX8^Q_)OSETB_-U8\ 
@N4 -L^WD9-N3.WY<^"@=W TJ%\17PG.$,3P8K&1M('8 
@4!]Z'?D?:O75^4D<GO*;F@[^[2^ZO%2OE\1HR (1858 
@MO/K()ZMCG6?@#9#AW3*!#+/9>O6L*EFE X;6RQ[M)@ 
@*4_A,3-T68)XFFX9+W);8&DOK!F[X7;N?:#FGGJ.L3  
@%YCV0^D\S +Z>VJ;LA'FEV[1$U;.VT"[.\^3_1#F+/  
@!\X:"<@?C[:-)Q*^2(/YS7_U!R@=$#@L4X>TK#5Q;?T 
@[>'# D,U$J&X8^2:VI"<$28K.K9J?M:NM,"<H*5(I < 
@^&)9G35:I<)R.$M"RQW4!7,3T0):+7FZ/U+A+B*1B,8 
@O,YT^M0/S@9X@;<OUX([<M3;MX./8_K05XU,VTP,SK$ 
@@R:*(/N!$$8P]'?[/GAO##<O>0R?6U"B:+RHQ>WU$E8 
@6;V18'J8J*-P*3S0>-L!-JIQC8^\*YV= ZEU9)WX+)0 
@FVH?B8NUAB#1.^F=#\]E]V3"A<!Y6@W7F",RJ<*5Z$\ 
@Z33!=!$^2ZWB ^C()&4@]MBU%(G[/P?_M:V:2=I\BT@ 
@EZ3V%7UAQ'P;JQ\,HE[O:*+Y/FO]?EB.*HPG8QJ.G!P 
@AWA74%I6F65G61.%;:-$= F7DX!D8+#W&*_@1P/)#?, 
@"4P:)SGJND;=(*J.+8]D*:<=<\:O4]&J;.ZZ#T =8E< 
@%0,1X;-_BV:".X:#@FZ.4;P]H,PK +ZM55FK M M[30 
@,PL=;PX>&HCEAT@@>-H+7]M$3&P9OWD9GZW8E7%6+S, 
@>)R7VH]BJ)122.. 7D1Q",E]%V(NS\ZE4H2%_!OF<D0 
@<S1\W;#M"W]8;/0#&6U7]QZM,[N01P/Q WV@+IZ;-00 
@CC%I@K)Q4;74P;F20+<"\ !E*JRE*@25#2:1(T@M]=4 
@AY<:'(X4+2E&FNGYD,^.YI>BFF0+#=:#&RD[A:0]?OX 
@>1]&0'=A92VED72 @W@ 1.K<M5=2AB[(G6MQ%N?17RP 
@Q^,\>MC++#*7MIBM:IV*O_>A-*T=E4KC(F=NYWUBDQ  
@;3S/^OPQINY:MK+XXB_$* :-T$(]MTB8C H'9/PG&0X 
@\O(?%BM>*T@+R7TGIO%BABA%!G8DF/2GE6*AKD_@N/( 
@!,UEX)S,84J<6EP18S(4W8Y-^<+<N;;G5[GME&,U[F4 
@(#[P.=W+0II!I4F;5*<W2)55U<!-*]%B;D]:A>9I;GX 
@>_%$1;$3ZK*DKB;60;7Q5?-KE)%"2LW"]6H.J"K.*E0 
@P[JE?@ #ALX"(L]+YVWC8F=[D;^+8PI$"/-1NP=9X^  
@Y8&).O>[E/A^T\?)_@,O:=]!GFW*7 )2QIM!PF,(?E4 
@OQ1AW^3>H*9LRK<\G0C=Z8.SEX1BV0WFC!V%<-N/A#\ 
@M/:&CMCN@<9W2PN^3W++.RH)6=XR'[HWO"._&[U!WTD 
@B#ILGGWHD-ZFERW0:FG5/;G4V[UE>;KC8/]1LNB()(4 
@_!.@8*/S3%&'X&G[H>F>R>\U(F$D^T[T!W:7UIQ!;D@ 
@]G=Q&+Y!O7^,VL-#XDYAZ@$HM]!_J)DJMHNQ@)R!V:0 
@C7?U[+W(<V<OCR#);;> YP\R@/8QNVA&@8>>FN9Y78@ 
@KERO+^85N0R.XIXAK91!2?\K<**68SS/QRR9O%SS+P0 
@)KK$BHPT_E#+JU4447UKU!E?XQ^K#JWW2CDQW! _A6X 
@0L;4N4I.Q&0_@0373_W7@)@R<V:V.2 BQKX".F4;P3P 
@"P!WL%TD]M^/YCS4"^?-1\XAM7X(W%@V<D3($6,@XBX 
@,W\Q!L*]7\6X-RI\H6@#SR39S)*&^P>\"Y]+U.@K$!D 
@L3F&A/,R>F7L>30[:K* +Y^!O@6&.WX6T.ZL+28G=10 
@W,,#)EZW^E/<;7=Q'.0B":/*3[.7;,:_DNA\K2T$;R8 
@6[(\8DGB>8J?D.B"-D:;[8)3VAL'!RU0RI%RU6,<#S0 
@ILR+Z;C(D_:T>'#ENV>*,[M,F;0AVK@DW3%[%+2A'$< 
@+N+A2_ C!1_P-YF[+-40B] Y1>H$*T]W:[#7JV X]V, 
@;CH_?UJ;L!@8"L"CRG*(+'!67XFU.:AXJPVOHL@[I,0 
@0&7Q'@Q/L33*_7Z+(I>IOYI@*VJ,=$ IN?$M]]JH<+D 
@6K%8$-A4"I>:OV_:2;O*E ]I[0W(#"+O?1U\!:!\3E8 
@4=<!&DYCK^PR"OK]:=2DG"<26L?O['F'Y.EU> !A-_X 
@&'FQ*[^LA447KK["ZI;>)P>"U7I0QGAP7]?)FW J>U4 
@+YTV+$=I3/R MA$^RSQ*0(F!_F=S&</Z >F%8DC+&B@ 
@\ #F4'K*Z*4'G1[K]?=5Q_,1,6Z [8W'5%9=%)>5D\( 
@!*2+J-1"@2L"]]*]13>CN4+E8AV%K.H$):4'BTEI;ZT 
@BBP7HP9(JF'G 0ESA7J?-R^8+)S2?R&-#E(CW2BB=V0 
@ 8W L<6K$,.)@2)U]*>D 29ZTC=%R[L/A,UT<:X5'"L 
@9$"\MRN-B9@V-'2^L\I['0;=KD?]4S_6!NZ:X9(6T*\ 
@:0FZ3$;CG-NVH5[U]&Z 3,=A?1\FE5NY0PJKHC]'L1P 
@B-E6LQ2?*J/T\29XC D5S5UW!P*(-J[78Y8J"A/D#T4 
@]]\2;Q/B'H?XKK?,511=M')<%<5KV..B(1MDI28Y6[P 
@,_"M1"&R^O[JZ6^ 7$?%[<7QORCGF27"@Y*:SX,O6%$ 
@=L5T6375+.#'_6.?O<K0M"*C495<3-%:5V$[!A%\&VP 
@-[N59D1"!^XTB?AW-RN%,C>/T/_"7JT<T3)&M",$\ZH 
@PKE*K?]TBSX/>><U_>;7/+C#J&[)F'@0FD@D3AKCFF@ 
@S39DT>&^"0*_&[S#\=:* MU,U8V?N*@8$E/!3J8Q>L< 
@DT&[-O[9/;.V_>W^9HRPUOW3:JQYI,%ASF'V/ $KI!0 
@)9S:H2!_R">3#HI'7^?5P$X>;PGH O'ZNXU")$#VYA8 
@]MAW$I=D:]/&)9EPYA^]7=7!#H)F&RXO"Z?PG#\8'ZP 
@][N)*N%GXXE3G==L7'[^Z2-O<$8N720R1#<YMMCOST0 
@CG2K]BE_?N[=-;!\V9XA4M0I6[\(I.R9E@X);_@+@B< 
@9TR<!+-26$]=;=<'S)=^2@1\.D:16Q!*22)\,4V$&5\ 
@,1BBD0+TW*2P9,XR?3@C?*VJ8[S*FJ12E"[TG+SD%J$ 
@@\E9Y6W)KM)G]7!"GV+]VYX^[YALPG;)5C6DG8Z.@OP 
@Q?08^1U%9C,N3$O:INW23U79J4$R3&<]?W_FMP[Q[&, 
@O]1=9H"/]W@Y&\"P;B(T/(/.T?_Q0*-1ZL'A=D>)^\D 
@SI#1(DB-&DOX04.3TGW-,X%O3 "A:;P,)3?SVY8 \1, 
@JD&90EM8.FPMX(34L8E96_N1Q0K'TRW21:+F26 7#&( 
@!38D;X6*Y]FB!Q+;1_$#BQ,2MB]/+'2GD"^2MVK-Q.@ 
@"1R/(!A8O:8A^K3C6*[#%%1\V*A1EQ-\U]S/-51NGKL 
@IIL/&Y$^,/S@+:)"59[#WM1'>">:+\^P2*UWO;_V31X 
@[.F'4KPA1V^N>OF?5^V.).:5*D-(ALI50(Y_Q\K!D;  
@@@7H^@P,]C#8.,S!Y[-;D ]5;1RREH_8?:,HZQ14(U( 
@$['B&X=IEYF W8HS5UQ!T>N4U#SGC!XP!!Z5#3)$B-X 
@,$]21*L$!67.GRK!7;C^)D60UHY %+.#'="($.IZ9(T 
@ET/;4@%Y^%K46^.F<^,ZS 5C6,03L)NBU6 9.M/BD?D 
@MNV^+)W-6A('UROL4T!4'JET7H^NB(-#!WK!R6MX)[( 
@+EG^@&CRK5)Y=H-GI 5[25&!?="3T;-SDN<@F^*Z9,( 
@WAD3U1LO4D+4^X<SX@[HGU*,O.7Z0'7C_\:61("_FE8 
@ (5]Q#L)=_U$:<?9\CCJ==,)$A8QSBS)TE&]^%J=*F0 
@A$T?!(@%V8-B?[G]9Z5&-4HQ75&_\V14I#6(;3E=!R( 
@Q7LLZU&2)W+^/G].OUU!<Q14>!,[EB8-B,A#QHBW"ED 
@'J?9#SW6>A+R'=L\>A!J30Y73/) +R%K*A8'8)SP=V\ 
@E0N]_P'>K;?AC_/.,@B](09^]K9:M.IADF*X;@R\F2T 
@F2SV!?!9K>O0VLD\FHRQ0#^91(L[QG940@M]SG!1;W, 
@CS -2+LU95B3QX,GX:LV&*STWQD=P7'HO+]+(M4^'DT 
@^7F;4;=7V<Y>T4+P>(/1M1[)J:HC87VF.D 4 CQ00,X 
@6'&M'"QXY84\X*HP?VR,>DL^*Y[HS1VN[KDQ+<BHS&D 
@N@@?^,/$#X..XE-H7_;#4VQUX-)B'+[U@[^HVE<Y0'0 
@M>:^0>R"'-V+DKDR@&8#N QC_P(_ZNO,5SR,(<Q&YO  
@8':-#L*/!(APTW<8*!#"*$)Q#K.2\-O\J%8=BGH&O-$ 
@"L%VD!;%\(="?U5OP$"6WR;'Z_TU$>\CT;F/YEE]X.8 
@V<+Y^(%*!C%U"I1*XGZUX55WLM4EX1O[;&3#_507/P4 
@$ "H;R""F>_L Q]II+H6_7N.:BE:Z* K8OH=7J-?F^D 
@PW%_Q,SH*-:SN>1N-(71'EJDX@AC?F?6N>2[R_2B^Y$ 
@;9?1N*LT4\+3G"2"O_\X]' H@WI/X-AW&+HI!?+ FZD 
@BZ2]A>OR*^]L1WL$V)=I?1QY/9!JW?][=V230*]0CQP 
@D!4OQ(XEDP&@DS"JH)?A=BGFJ&'E>8P:(@F;LBA'_4T 
@G1GM9@;3[><3;6AO] )%W(2,C=27"BU?<.;F"-[FG:, 
@ZY0DXD)@5O$XK*HX[.'6XP+])#*- 5FP_[;[';?E_%\ 
@VMA'6%YB]0#UVA<YL]B>#$C/1>S[GKN4M^@<!%Q)!Z8 
@'X1T_4+TWSQ1C9AO8% IQP%'O"R*G5^M0E/+DJZ6XMD 
@(%RS-N.\'884(@LA< Q\TEGB(G@M8[D"'!)!@+3H:J, 
@TF.O-<Y=\$U(5]+3HIKX9K]B*L',0% L.S+BPOJ&=+T 
@F@&^QZ*BEWIC5N1&W5M >?'0BU*U_I^KRO^)7:'VLL$ 
@[>G7V:;H.0_"C4\+ V)??M\5L'>2[M[F,H_-V5<.;AP 
@D6NX?;'#^(C :)&E+H[>4AS*RW4-=6:W 8 :WML0M:P 
@+;AK#J!HMZ2P>MDMI>TO-J[@:/YO"TX$\0E871=0^\$ 
@: 0AU2?+><84O&*J,0&\",9NEF%^,<./6>Y5Z#)UMZ8 
@N#X=^5V+&WI*.HXK_8]*2[<*=[3YL 4!WSRGE!78H-P 
@ WI]\!B2KL>YT*()0FENM\44M8*:O+/05/Q$LL-KM]D 
@?#Z\IZ04G]Z>U?_R2=E'F=6MHME+)&')MK261#I7H\\ 
@.V:%ST;7 K"1P+N=?0F8[\<"4<M7MEG;2/$;H9N=ZUX 
@R)]*\(HT&D_FT;T\UV)TMCY(B2 @ET=.DP'6NB]QF"L 
@!5VSA&\M-2*#W!@]X='YN*JDW"&M4JLK_ )S=6(@(^L 
@*Z5>+Q[:2$"!9C)GR^HZE%O,QBE]P*^AUT3>'#<6SK@ 
@P6X\G?&>=I)J(V?/CZ3D3X;&E<9(Y#P-=1;(QR!S8A0 
@*H S%:-@6R!M'2GF4U3D;CWIG2SQ5C#_,Q-H28NCO)8 
@FVV/T$P/D@H<T5GF"^J+4TIR;>6%SLG;T9@^V!-<"/H 
@-YI8R./\AS.ID_NL%.+?#[\/A3AQ%I*_Q[B,!"]+< P 
@EQ;OSX%&.OB!AC&_;QH/:GLU] Q.F$TA[3^:+.V\):4 
@+5%P?5-CW]Y+_H.-CT+L#$]D:@&9M>F_,L@)AM!ZL2@ 
@W,D!+\'0BX^KR=0,<C^CL3Q7W\O.24!ZT]Z2?VVR6O  
@\"--Q6'Z:B1-2H(*OQ 9VCV#X?LEE)_P%&W:/_5RL'8 
@%>V%%7!/AYXF41J&F&5:,M6$^W@NG42ZJ%%52GIJ93< 
@27!O@RW02Z_.="U.9;OC=H=S-<&%9V_N+ U:A=9V2K( 
@X8O:!<])CJ?>C*;&[?A;FJIG>?3#?R)SO&QCXKK][8D 
@65X;1L,.RVD%_+UA?Z_GY 405^-[O/G#&#C ?$/^:;X 
@RI-E+E$;CE3VL4=JBK%+/HMX!-_1=4+PA &S*>VC*Z8 
@* 4I]G1WD;Y4WY$X-ECJ-D]"W8$FVW.X!&"3LLQ:$ T 
@@9>\3+G@:,FCO9&EE6 6-W@N=+U"G@00;=UT 9+8QK( 
@;AE'%M!47V.Z<Z,H5BT>N'T2L\8\7Q;4<^WV8@G'>+0 
@XR#0TE5\J<Z:^==_6]P"V<1C\%D^?]#_M\?<#3S/NX@ 
@"7=5+<@FUCZL;1@0# 9A=&>*[)/#87.<D#>8-B90*>X 
@CJ3\%ON)5:<SPX)K7JP:0.+V_U 6-I<?SGN[UP4&-"\ 
@P-5R?P-LS+Y.J'P73H9'!@4F,6)OQ<G?J/=) :GU#*4 
@A47'S?;KT8J&#/A2:RB^F9L#=&GI;>,RU4HMP/8FW2H 
@4*AXOZ]U-[[-H-*HH\8V 7(<>1V)%GVQ,-ES<GDK)U< 
@6,7;+!L8<8$,!@$?DJO[&LB-.E?=I SV1X@P4NVL$\0 
@\B(<<10FV%6B+Q*2<T];;QU8Y5M72BZY#G1]3@>]((8 
@.1G-B5G^GD6RYSRGU=K\6AY2=QH></>;VTD)^&(D6\X 
@5# PQ_,('Z):/3;9&Y<(FOA:DA!L[U? #)@5++#8?BT 
@Y[(XNE?VUO^]IR1[.?EI[<@\8DOUA\*%C,Z+XM<3ZSX 
@/WUCWQ:UM+NQ7<8C'ABIG+O&F\F?,)V@1'/ZWJ]P2F\ 
@;A+9K*;GA["R/8A,G@^=VAMAV=.D[KO-9LQ(@9NX'H$ 
@0PG96IKGZ<Q*N$KE19 81O:CD$QP#N6\@);%[%_"W>D 
@<&BFJYZ4XCDL%PZ6(^%FG(T9+&<+9N&Q4XC1,_[</ 0 
@ZUI$;VM:\OH@^VP=&RA^T!?"U0BN5ITU%I_R&XB!H<0 
@ZWJ7/T^.3U>LIUE^:B5A1QG:<].',<4! K7GZGY[5QT 
@6$:RRU\.@N!R3FL6C1F6$1.L33\: @$WZ2YU:->W(40 
@*%P"[S%* ),V*(PS M&SB=>U)NUF[?)I85,&TW&;%LD 
@E;/-:_H9&^ZNWDGEF^\C')*O#\Y#/3G1<+(E+>]Z,74 
@))0C?-XC%J^A:-7H&5I)&U4[F5'WDB0+K*KC06#/X*H 
0>NBZ+1MQ3GV]9AU59.!"E   
0)[J=,^3<W\XW5^A$=ZAN20  
`pragma protect end_protected
