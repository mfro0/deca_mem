// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
oWlClaj7YX95YSzCKFKCqiSz7oNHwe3rkNBpMjabumCiQk7BR023LzQzjOtcRLz2IdvEXRTXP4p0
xLZssOH6dLVBCh5nn6o1FadhucyIrm9HbAz2ItBUKXOzBGOFyIiRB4e99+OCXIOMKcgBhc3okCuU
0hJCldh5McqshkFJr5lQRDqePkN2cTvsFEerqniZMRLkwDFHmln3tn2CL5o5GqGfJqfWUdl800xW
QqIWzKBMdi6vrmuCufBTWYY7zNXMx2M9yVPgjXGoUjUm2Re7iLRdLUjJ/ewMQhBnT4hqmT7drWri
dQ7duw0owjY86sY+auvEyAIPXsCATM/h9vH+2g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13456)
n9hN5duyD5EfdhZSpxIZ5uZwhNtarJCw0rd1Ium+maW3i8RpFmB3uBx134bJSgNsBVWiUgGnQg9k
eMrK5b1J/3mh7T3xZ/XokUkfek+w4XmLPLxahYtsyl9rzwD8VbbvKw8PkbYC9DAOdTzQmTTG3l3z
JacBm7G7SRrgj1wrrqGIS5o0Bkje0oAD69u5jqytjrRy6HDnnHtP7Ilmcs6XiFdLA5B4e3/i1AfT
v7J/ZChTdSfW9WWwn8F2u1ej/F5wnlW+WjvZAI0Q7Zrv9gW38gWmbOq/RnTabWmucdlL2BrHn5TN
+g6g5/47oTyhSCXHG1XsWlm3sNoEx0hvwOGW+CWudOpv7DAftEZN14JZRn9Iao6m/uFoUPMtTz8L
KcD7sx08jZd/5NRMrwGXvS//eSoW7nxFoAP0YZROYnYwl3D2c5XOI2caOKYRXcTdGvWBX1BoZHIo
JgIquKXWhsidsd28JAqw4XsIwyYYK+7dwfkEn+5jSIZw8UcEjAo7N5KlOsJb4mbzynPlRjb3o1KY
l97iJZ6ZCBx06JOlyK0k/c/tI7DytFNj5rHBIpYN3LGRAZtsDzsRrfhnZZWIeobrcWw0YqXKAhuu
bzceJalmvCMrq8o11bHEgv6lO8uEXwFJobV7QJbqrZBo0RD/7vZY/ugCQCfieegkTcKEucLaUDSu
gpVnfgHf2h/WHc7XEs+Jnwar5vCXEgzTv3sw2qfnt8AUbPxu/V7RuVcgr5dRYaT+KzzrOHe7p7Qa
6D5F/cOIRE2Uk8VpizIHVhNBKfxu+r7gFtrCT8e8vOyWAgEPVv+ufIctjF9Iuk99W9nOJo1QTH2o
x3u1pQ8k3pwZDZHWUbsRvtgVEnyfVfMnLqK8VwxnJgWAm+uz1tyxGlKypxXRHbCqlZYOwQx1pEqq
/rQGim6e/dhxkbW0k8Uqqly8mmZzTZz4pAvWWxwZi3NXn1WtMUGOyqRCG/us4H/0XPhtV3XrfCC0
0pAYBmq++W1zkLmzwUhx8/ksnBhT5B+mx8ZsK/V2cI6SyGpjUV7a1npPB5hQzndFoPRyxC7N93OF
0g9YfygWkoqBpZGteJUguy1sKJ3/vXI+6bAMCqGaux6vgH2TBS4uUhWnu72oTnl/LoR9dAquGZIn
43wpZdprVFbGJAQN/FFrDSeIElbXqW29Wdd468/jmN8xd0hStKt/fVLR3LnwZG1cu5DrFTEjJO3D
tHaY7v5YkS0aSz2YwKn6MbNKRAFlVyNbdnW41u5qBqaCclRK/RyxuXnPzQoVcQSs3Qn7yTzyl1lW
gnC49T+KaYTebxEW4Yc4VZdLuIIk416boO2IQCY3xj4conQvWT+IayAfEdj34qDroO/elV64YoHu
BQ9SORGqtJ9a1DqXgPaHYyS+CEzj4ShCO0N4dAUKtse/xts87Uc/LyE8FcE1gs0GNiRR/FlqB/Dn
32Ej1zJjA3H96NQL48XN9QKrP6tmhlXYPQzYo1+sAE8L9BQISQ4YCgdyYYuCMExfhUmJCuYl9ejM
zT9bKP8l5wxLc9e52xNE2bZzgrv5wDas/J4CaHs/MdTDgdwEZErcTr/TzFJfIjQ5g45LADp/iS8N
6dopTVb6NfuR6BYDGMiWSNQpEesyXNa3wZJH/N/n08WUHY8HxsMwfPyo9w8wSCNsf53VYNGPTXFz
Vgb3aF1aEQumZ3vX1DN+pYVaTqHUrnrxAYR89DIdy77rA0/C4BkXxyBkqTOZan6sp6vpB7bCLCFh
A4beNibIE3SfdlV43ErOUL+DH1MxooMBCkrlY+H7qunV9KJwxseQwfIc5Bv7sJAzFqWU+hIMuqav
29qd/G6bt2e4WOm9A6CommNZszzMn8WPeK6loCvZTedALicOWuINhWFxq9BBijTfKV0K0VNnt6fx
xsbmlqTsoDUV/9AY9qOiM1mRVaYpc7VH/wplHx3eg4iWiMW3Heh9byX+HHQz57LvvK2LmegbN6oe
AOQTN0UVwWtkxzM2yR4yaGEtbv8nZZ1nAM9xCFkPeGbx7Tku7EP6Kl5yhmQP94YT41suTyTi6xvA
PwP6sg0HOXSBPgDbg74wwSp717L9s9fC1UKC0o2epiO1aVA58jkHa1NRqPOP9gwNg2IJmjseuMc1
/RC0q89ju1o2kTyDk6Q31/Qov43Uf6VAi6wo5iv8QKDQG8FL/MYO+Q9Nt7JhjOkkD8iFwuqDnbfG
fGGUBdngDNJbu+aYnKNsnEY6uL/ctYuIZon8ko5oMeJwBSaRI4IBsBkQ1U+r1AYEwMppqKAfQILa
NeUk93877lgjSsYESskJVUbEGzlyxoM4NM7Bg5QsGwOuTxyLhgPds2B0y0c95ZF0zAVKcg5qrLmS
mcs93+62JJwb4Z3fTtRsQVlkaKH43Rz2OaKich6ufMmFWpty2aGv+M+obHgPNkICt4BASOGgWDtu
Bz/gcRQ7or4IrtlPYgJOEoFZ6Ci7apfIeJqvebjgGKeOQFJsvx3yCsmDrX3uAmTgHoN3gdLz3Zzn
KaKAm1Fxua0CJkXDma2xBk7W1HYxR3Obm1IkaRgKpO1eEJ5tNTtHpcy3gpIUztDet21lbqPMvQCL
9YJlYcjAN07J8vCbb3dXhTvw0CqzpXHl4C9C4gXcUcxNtbAoSGf55712ymJdH1DuhZHB2fswnBlh
3EdmP4/0cL8n6lWw7PbrooBB8yMt4w9YffItS8AnLkwMON1CA+E1wWIjqNCm51rxsnP43rHcf6Pj
UmGKLKrRSoLMzt6eeQ6azV3a/TUzojm2OwztIKfhfwz1GEnR8HgqRmoD98mguuUTg1k6jTMi5nip
VUZpmQRHHU1sGuOn6o7EoCpZlTCebXc1g/DPCcdtk2+xpifjvj/iCzktoFcdm7UJqO485kb8XwFs
IyXSRMDsa3PfC1gZ4rzTY2duPLufjmwZvFIR0oG5TzlExz1e/TPxsJ1ahkXFqseiZCW9waBir6v0
E07AW7Uc/saDfFAx9GCtmBgxt9Vi9xe905lIfzOPUsdGHpjmVfxESgda9ZYyIhlkMaWIswISAB56
81X2tx6G5Y6CVD7iSum/nqWdZzPUduotorYR9kXThZVnI8y7gToqKtbyd1YXCxs11oK8qftlpA4c
+IqaAhauqPFkBpauqAFSBBlI1qc2IKeYPVwNZ9mILOH8OWrnorP8PjbOLhFHbAZFnTHGvZECPB2g
YSM1+2vIe6svlgxBm3qyd5CTB3hsjj9ojD3rQC6stynRqmxsL8434sJpmJf1rRBpHGEb7LqlyL1h
cGgtIPJZ4qCISCEsLJpFUyGZI9uVwgGATLDSgWKsFSqvArvF9IB1jAU8HZwbZqLV7qCZVV5Oy8uz
rrJ9UhTekROMmMW5Hvh1QaDhvSY7CmseqVygHxspTShbHYeIyyUzFCP7NOIVWotT1U3wHr4I6wF/
b+V5u/JmFEBRIWjUzsTG8nGCKTp+DwOs7YjP8Qfp8SpMDjbGgvSp0xpMDxYOkk1a2CTLSnKRauAb
g/ANoVmIlzqRlr3oPB7BCDSTp9UbyXO6ZyZZquJdY5XTH5Lv072eHVea81KPoNmATwcwv/sdfZhP
m+fVsPSRRv+IpSFA08sCxHDybDv2Ynx3AHI/fPu5Sco4qyNbEsKtOZJPDcEiOjYOtL0azIhysDM2
ZCwEApvcLSseKDN7S6k//G7uXryJW9601py0VjXMPCK7E8UByipvFTPfdolMY6kDzjNX4y20gbnI
LwXFrOrTFnaB/fF/HV1iOkFl8RNY1rxBV2IRGSy/H7dPiBJCrPbienY2UKnrav0B8k2nzwZoO21o
zP+jRZrEarIjpZuh6fSbVBKo8vY6pxfFSok0tSv8nHK/W9EZhKaMocdKSdlnVEoM72qAoRGN3W1J
j1Tome4fvz2r2jo3W30IhS//ynQtyjPzpQoKRzOBK224KkQIGLmztZuNeYXxeCrAcdH5fBcOwpbq
v4/QefbKHj/yu8d8eb6SWDm6qRI1h8GtEoX7mJq3DdhmW5KgXKwS4x2a6hv+0FOnej6ergRlWUWh
PR6v0ot+xIiDq98mOLFZqZSF3Uj3oMV7Hb4SbsayHTBKLk8psESFiQ9VObwBk/3CSi8+Za0yCWA1
Wl2lZhNMH+PCFDWcHG8pTkvn27jjzI2ZKCyAWOjSxCEWeH2UD9N8Eu5x3/4AlSacGmPlqMYlh4zM
/rKNDHXZOcTuWAQTpLKEyb04iN43kUkgePohXsnvQghuy/GZzi95tVEVhTaPjlwsx0Nga+/8ztfi
y4+rli7IFwmYgB8S2ziZSMZaE91Bz5WCr29pzkD/hLIwQxZbSdjmh342epQxZAYw/DQ0Xi1+l33N
0fkOkQsZCSaubtyMliA44WpX0eJDX1kGJcDwlrBrKs2Zd5dhUH/yGVi/fD+pcImP/w7cq6qpMsBw
nTXBnOHMhsZ5owoaeeEi2WPzD0ZvLVwIUhp+VTuozKFnjh7doh/40fO5Gmb5NlFRjBagG5INQXXK
ALkMmTLV8OdwfjQqD19jz8tpBp043jOYAultD8Y+dfOXq7PN70WY8fg96IsQOv79TcMEK8T2Wlvb
KeqmVJnn8lfXSdRFU31NzM4zp+QY8i9mF2uFQBszC9EU/ub6RfNc1mf+7TIu1yIFWY8jx36DevW6
GLxjCijgu8cEH0argFXlwrYfA/I3QgjOf4S138HfCKgSmen4x3oTDEaG1fNTNeVlhoveVncimDQY
JTtndP/MWUBDhfNmG1Fmr+3oD1mqePwchX65JUCwRUsow+k4BwWdu0Oy81VrHDc43bYufUnwPrWA
p7lQalRvZyfLqSRSmzFIlX6Z5LnYnVLPir159fKvFgD/fNUbg/l9g7/gIZMSDkmXmnH+Pi2lRviG
/NiD0oDcZ2oj8GhNaVwOCPbtWXq7RJL+XiKvJpvUNV19dQpCBIQU9SyIIcq57Gjt7mIjJs9dSla1
YbnvUIm0/xoPGgJQfOQgIE3DurM2anTamzbDW9whM6Jesr/jUPF1hRnoPJPlsDC0sDU9tlT0CJ94
x4frbbTUfaTrgT8Z+tpScHmgzILt4kOlps+twq2ioLgKnaWto6eglTqPP/kqeT5qHLV0/fAAvOnO
3IyU+UlvLJU1P2mYB8fRE9dO7zpjhbufv051yxUudg7iatRuPcvPeIss6+nG1mBRvVp7HSbag1e8
UMqO2rJ8gbhJD+tBh3/IOkZyDZXbC5/sjHd5R4uJ1G7JIMwodbDtFPKVkqFwRQJqzvLdvmkPeXD8
O5yn35PjtMUds+W5I79e32PQOHtTakBsIMILjwsEGloc1QJVBAck7F0R8qmlWJQ/C3yL2ylMFnMy
jqYpdZwa3NyAMvVg2iuApChxffwAJvcTALcC074OvoRJ/mgaHylZjaJDaDlNLejyCyBos5DdeeZZ
iNBgkc+yEeC3R+tLXAgOjpBryVIvN6jc7ROGuCuSjNEBsY+TK/vwTfs8tovV1SSLoeHT7u6rCYBF
Ursj2XDd7et7P8YsBIMhuTc7RxSs176nZPY5XZHSqmmyH/yKDzAgfS/jUjPp3wewZfZDFXnpd366
XpRXMjiHn+gk1X7VcbIXJ4UpO7s7+v76DK4HvwdfQPl6dF9zUIls0faJwI5KwH/3DDu3YCZAAOln
MHb0i0dK/WYAQTY7HrjHoHure7UMa7OIoQAqgdMRFIcE7odmcFg6y88lvX5e466WeHfN8T2rFIAh
lzrFx9zfN7nKFxYX7znCdzRtID3duryCFKua6EVSni2/3lSsaav7LbAeZNKzII7yy6UQ7z2zsNR2
/Tly7SDZXn2X4r/yvrICm+yxcYnWqhovVbM++7XzpN9mpG/a0eMDSdVGbpX2ejydT9iX+eeNzLQ1
zIiOAa68xJzsLG39NtbrawIE2eIFjTL6Ts9qJuC+FL4yLWeAzkIlyVqdkE5LnQkY9sSVRoBjWRUy
6GyWP8dwI+rjmfLWTywurrpb4fKEGxzFCVrRJw6nX1m8SS4EvZWU89gynuVXrEE8GTllhxWWIAHx
7wxvnyopCMHPABpcJ3pp9ry1q8QvhbXu0TpCzYgHej8YlbM+n3qcRCI074KNkEdbfmeJLhsGpGdg
fF+EDGLmkp2EYsm3LmnZvvlmgN6q2+0XUVizEKjWhQMPWB5f7IHfJExS/xvplEbAibjSC+Sa++V8
WXQPyrNgGX1uadQpFp5Y/+BqgIFScABTcw6wyibRD/KahywtknxchKRl8O2xDVMLeYwnqd009aaq
H1YcK0Ww6k85CWRoEFOYig3eGenTt9EAVrACi7WS8ZoD1eyHhK3swM2aM/r1L6s49fxc1fSHoenk
vy1XVqbhAz7S83zK8U8by9Jy/cqCn2V6ypdCkbJ9TXxAyK0GVxXk5/GUXubkUWC3Er8iYsZkv0vX
b2I7R91uEqiowJKgUKshD8nheYm4MPPIY5WuW7GYinuY/aR4cpqDk9aUyBA+HtePt/TTMMtGldwj
HbTRCywIhuGjqKOshFIfZeQDboxd1IHyo0z1AlTNFS7a2g9IU3g3xGBXKYdFRvsCxxdHkqHvoNPw
QXj9cRr1qcZL4HfuzyNmPqINjBjgaAfHKPUH+ijy8wooeclJEFY9e/GD5gYmpI73tqW1ne7RwnWM
z50zPVdrCgXBnGEan8d1OY2pxpVtWmu1WLIrcWxd3Ie74pUpdsDC309RpheQFesH3FUGQvMviVae
7aI1v5g4BVZCcJL4k5gGIxvRaKQNlmh8easrAk3cLX60f9KcjU3Scv8G0GN+kwFJjOi3RVu6PAc0
Z2sVU3+j9IlbjUOdI09z+6E2qXWKsjxIHs///kJDGtxa4xxdLSJFJEh/bI3MwyuQq/0NPZPCZ+VG
6yn+C3cJ2wyWde2oivAZ8dkg+vUWjJvnKVE11fbezueVMx+Iw73nG58e2qZlR5006gAwajN8jOyB
R+nj9neGoioLUYQ/MiHzABXHRNNwbM83KUB4PcQDHSll9XeksyP/oQUs3w0kYWVqcddkx8b9stvD
S4rdeJJUrRFXO7VgdtizjmXja0bDAvGbOQI9CbCpHoOTDU9vYzCRnHjj4I5edH1OV3AC/Cdxkh1Z
bPcckX7tAxZdCrlngO66T+AEA/khD4euNlN5EmR5oFtH7+074S9kYw6oiBdHdnJLdfMWDZHrGkXG
b9+A76ZX9qKYIyjTmxMK2ySVoAxT34fUHE0EM9uR60ABZCKW9JOW/3CBk9GdBLcGpPQO23JA+AUB
A48rgU+AYbPHs3YzEA/3R+F6GV0lOGUTPl1viMVCpdIl1yZM4Fyif1YdrZeoDkVqqp35nvnikcP1
DBhsjFb60+MjKKd3FsjhmqR2XPJIjWd16hyxwxe91yqWa3DaOQrAqAinFoR7CdaKE/SdsB3moD+Y
7tg0XXKysvkoFvjpIgHmySbVvDOpQgOZicOjX/dwhdYQuvFuGY/8bwG3tTXntwSD55FZRBB5N9GV
/1Orvj8WaaK7pE86b8srUSkyEaAD2JscK08Fdfy7k+th3f8rP5Z/a9wAsM5cRuVnip8Frkq6lW9l
WNFfkozEf7uCMoC8j9QA2XECdtEISloozf1wXEqT2EPyJeNAFolCLqPoMsTJfR7FLI5sqcEpWVcs
bDewDwVxMuWhnsQyWnEUjgHS8FINfISSnZs2/hbapLZaNDRKSLbXKqdipdEq744yBS4j8p09Xpz+
wZNn3JjJ71vhZkNCRcNWMAFdymu1hLfjpbwgrNceOWgtLPKTamMmbO9Do5jMPdF6ddASV3XSXetv
vHBeOaWHFr05VLEH+nG1t7yA3jvp39FMg63r2csHsSCP5bYmoCNI8Jv+ZNMe2T+D7H8k5LwT+7W1
ktnRr7j9omlFjzr0pL9GPBfADOAWpQUilaKBwh+mRVVyU0EYPxx/KqRlkTWruZnCXJBYbf66fsMF
8ckV5adVL8Nc0L4XAlkLYI6cuY7tLFbWm+7QdM9Ohd75cibV4OyXe0AefqxsuivMjvqFrFWIw3SS
L++T9qi75YgBl0Jqg74bek4xI4FbAUBg6YnLV1cMJHbHIrC1nQZ/Ah4Q0/WqEcJiOrZiLzmMMs0K
NVd6o9B/bWMnfJusheNlx9brUlElJ7EAx4ytP5BfFLzGa8UyboIqHl45RRwUhlljHByn6HBklfaG
G7h1RvXQfG/va4QBDihIWpjXiXEm9Yl837H0cB8rETPp6wjSz+OBLImg8PZiiQ4az14cGK1+tWN+
g2XdmtfFrw0CxIXLWm818YxTOQNyVQAPq4rSLygeCvLKbxhQSGY0UL/sWhznVVEgC+YBRBzSUCqz
JkoX/mRkqgKlRCiRFJKbl0XIYvXdU/W5ikS/wdWSEjs/FLX6CbB0sAwuBtSBZZ9a4T0aH3IkbIlo
aoFeJlraKGkW6Rl+lT6Mq9qBXPqo/GINjsTzbm1qFRXbqCQyMCgC5dZyWM3/ESi/KErLhKUt1aKb
nSestw1Eiva+HI8khlsnMxVms+T78onm+YoQ4wuZdbxV/W7x462cQ50S2zwI7ufZ4voRwn+NthZ7
WV0Rxqmocc/TSwLDVj+tB/Sx6V8iBO35KDHUgjqo4uksnDzdbZqtMJEhcgzy8RYNohNR2C7EL2ro
+T+lVEOrN8K836LrOmCiXFrvXc/wJR1Cg05AXR9JnHWVWDd6h9K+dT4hOwClOgCIV+t4QGTiDDcP
4q6uT8bwvHl8I42ALdvgkm1N0vOHCuZwzYmIk0AocbUl/EA1tiI3n89oMGZvIqWzYjhG46P9jAXJ
I3Fd9ISu432efO6DeexL6PTfdTlwaHm5NooQiKtXRxvIJsVW/VBKT0FWMy7nbUE7pPbOTjzAxemv
EUjFf2hPvISYbIAhylTiuj7bloNTfndv4jh9asFx7DJH/+Q8SnrxS2Umhz+DSli0/wRjaT9Tagr2
3ZUoD5JRBCL8ZmAVnzNJCiiBc1X5++DoZLB2vvrklUiQB2r6xB0ukAHC9heyMqHbppM2RS/Ztbb4
O+ASF5uRTWCPMIELHcPEnLv3nR8mZyvfqint1d+pHzrTd2zb8yf75D5cLOo/1eYjXGnlp9t1YdB/
pN6FqONG8GD2I//oSiuKKX9ixqifhibD4gkA+rUYhLhL3uGKDpVVTpZoWeHMB7vE8uK3VvXSoxaW
mB2zdgVh5E5Jid1SQg8uHnUJNWNYGfskKy9TueNetLIQ4Vvlc5ORoOVAkrfbuLeC7jRo04esPW3I
u4+X7O4B0xDFJIPZRvEy8VqRI6Z8FEVKWfIVOH7YvGUsc9GZSXwMM8silhqtch6dmGJu/HuaRsHn
0kad13U/PiHW4BnB0TwGE5ddoyZon/ISNX2ehzvBrigUyDBjHjbGQq3JUBLff12JmFDI6UKf+oAV
XVPUpfxhubFA+LrM2c/SEgVswEyRqZW953W98h/+REEDjKc/1tpBg5BG4WD7mNVt7IN7u/RJV+65
HCW/YHQakwxx8eyBe6Z5of8ELEOpPJTZwwVhutmRASQ7lBMsObId1zHxPWpB3TzgeXhfysgK9L1F
bl1GzJXmZ9xYZiH7hwjflDit3715VIV80j2q/qVRGBQQotjydvpwqRqtSI+Y36cfZsDPoPAeU6DB
MG5Ue8n6++2g/G6OgqCQU1bDRB8RcJp31vbI5CprV0n3/mairZHjQcJX5Uqcs7xfUYbbItmA6xxa
AECu3JulNCnmBNo0Auc042BlhrfwEmXIy27OTXSjcZRXchIMLCOhjOXPunoGkM7iO2yxmh6Vo6Ez
KzTpEbPuq+g03AASLS4Fgw785mwatp15eRmvv2t7rg0vDPYFk48nfHXADL6qQFgHgeoVMJ3l2Vq+
nQJlkU+7ce7EO+s+1hug1sjrjB3sC1G9eeKaQ5A/9kwiokKCy96Jwqce1YaMDfIjBruO80T8MTZ9
sk7iYN9DfWcQryQQ7gexgWvxDFLtP8e24kf6y7X1ary0fMUAVzBiRVWXydED8Im3sSkxpclZOg+A
vQRdixvSIFG8BuHEXFM68z2TJ+YXb6LK+FUTbYZ6aGPeUltNoUYwq0AtAIcY7MgtOUSH4xU1IDiE
YJONxmT7XFyMIvG7s7OJtV99LeMFbyIZF6jSatKF8JkSVUh0WYaxi565+W596xGHjYN0VoDMq+hT
U8tcNrdz9zy5RjTwgKCJNf7+djbtdR3NBYnpnKBIt/5ElGfrk/aJsNAGDO6HbBuu8XKEUfBqkB65
+fVfmwhu8rqlYY3BGnTS3ubzxe0iLmeBObPhQoySI+AL57DGGZ5zzIC4vdCt6u6n0Us8jgJktbGA
XBgLZl8oROQJu2st2QfACBw5+te4krhi+NMVnpP/VBmXSQ0OoGVYf/ljbbSUPX4XR7oNecqxaOTf
jVKT1wvUGmQFHPlP4ExVNdGyycoo6O277HeuOKBfnK2CLhKzMoQ7LbPYuP5G0HJ8W0X93b4pTBJI
n3QegBOhTBgQCMSZQYR7NJfTG0Tz0Y1ASdDnppYo8N5KE5kDPBd3boBPVFtfq7WROlXqg50WbTB5
gOthVeR+5APQRpyCIs2kU3ZDZ1yoAi+Ble5Kl+hHCzFbh1wQ94TReDxosgbZwBF3T+EQp/gWCQSV
hZIk7f6KSQIk68bK6tGQC9jjqjQif8Zai0D6LfgiiZ8U+qREE2/P2jc+Pf8hmZbyZfh6fsiDst2U
HVIm8h9RxLEbCmCAWF5ElWoZYKE46qRjDoRxNvTIhKm9q1cEfKx6sKQkWl3dJ1YLsyEGMfVcOJ9r
L7MzgXmsYsbGOKbVvLtOGAGdYvyofY+vHywlMsWnO7aVgqlDNbi+r+oMexBo8sJUU2KnN/+ta39q
5u4NOmBXmhYW3vHcQ/rapcsgJ+50zDd14E6Xsvk+m2Ee6h7dlXIXRuImUz2DwLaZ1wmpPl5XArwb
4sAscexwAunw2aRDi/RgwVTHkE3ZrSbdJjQz5+lUfkC9ZTh2j0kqpFpUj+UxqycMKTuPQh9VmiEj
+3qV1YxlI+MlmGbIUAuOUm0P11G9m7lQjavnIC8OiiDnpZ/xSuRjJj95H9gipqxPz+UMKVRx1Is3
OcpSwTNrigYtF21esNWBgZcR+NKjX5FvQXTkj00dS/M1R/1n58b5s/WdDHb1oni9lW8NT/oECYsV
yZjftvJr6BtlCdIsn39IcS8NM0oS0oGnkcWT+WbUxzkM9O5Dc+q10QSuMvH6HmviGTE5PDK1S83i
Tr+cPyCyJIN/XzBq98LdPf5OL8H6UTMnnaUi5VWvPDrtxUpX2xpzS3tZQQ4pTYaq0Z4l6Pc3ZDl1
IsRHZlmg7XgM3ldrXrlsQIH7O/CMt0m3B7QvTF7k45lTC3EHHVw2QQqtMutZMKQr5oz/QMDahB4X
KcewLb1Qxj3z0N3/Iqqxy0DpUfqbKs61RYApY+yYnITZ1LhwDBHz/Xs8dnoYKvQEG0H+V7S8nI7a
vKiOzNqJM7R/EcJJjys7BqJ6nHUda/YszeMgIE9s8TX9661h5DikIxF/RkQ23vXKKXYU8t5Y6ObZ
kv/9TBIRDcGJM36uy9iv+Bi2TVAoDudP/FNzdIgnZSBObsplZUhKAlRcBQX4Coaa7hdEw7ot4TPb
25sy8k+XGDiWQZoFlP56HVG/7KGR2WL5TIcpVMhrFZlySwLqEFNy9sjLCoMUBQOFJ3h8RxDy3eAu
mUmfc43xd3SoMydc4OJ/7tKPR/nEJtrjzwoFM4JiUOucXyY0c2o4qYMoMkFqiI2cq8o8mjD9AH2e
A11xtjIc5SZeGKFEQAi6ZdFMaivVLVcwGC3BiFQmynxVMQ/D7B6r4Lv0215pnSQ53V6tgK4PX+wi
UtVPRRCnLA3nh2wuHsGu5CNxWxIW3gB7GC37fPhYQEI34pqAGrYGhnmgWCtHMdInLd+GHoJqVExg
jD5fGiVWBUJe6JsFKvw8o4xI0qsdSHRyezSxJhlDElIH4ElmBpfEJ3fnOX274hjIuZ9nnohahfah
fLkA9nTJuSiU9clB9B0KvfEYVHTINBdEyPJnBc7FCz0YQFEVftZmm183twAKmgiJQaVEOFWx9d5S
7bxCTX5d+yMg2M2qZ+UiHRQqw62x3LciHZLVhGFoRIBNzi9gwloNqvcvbjghU83A5FEnqybDbUAB
t5JZLn1fm+uv7QsANEtw2jia6jHKoDFCtOKxW4PVGEfYewryeqWmdxusGOO2T2f02zef8jJQ65di
OI38dXdz60bGPk1YXviWLHmFemvTrFjniSdre9O7EjLRZ0P1Khx+ptv3B9t0Ed54D0g0ueaTyYNw
Gz84qrzEe9u4Jh3kUS4zm7+HyCaN0AOZVL7HoVIR7fL6Ck3hvlNp87mpCBWgzbpjFyTAoN4CffRk
118y+wfrCJ8ip+00lf+4Pq56KlzHAZ3N/cNZPWNAI/X6iKM0zSk+F3m2nhk5i4SW4+dMVSLPf1Ye
utnjnFeiPFuWFP/QQorW2x8xKt6FQj+NwAxLzmHTx2A69WjsHlWqN0nUoFZLmJcxBFrIR7UgZPhr
U19dFIjRjXzcv1x2S0gRKhSi+MYKhmLvGrv+jhKWe9rpsRITIdbLSPIF8tXiM+nJK1HmiGhQsERA
S3+2VUqV+j4/TwHAo+NSo3AowIYCRJYWgYBbFK65AmqIY9BkLm6Gp5kOfu+QAsDLzONVXdtmz6AZ
JBaod/lRYQMLTmjaCM/grpwqY/ilGSNpx71yR8eCzjIJLQIEuvDf4U5XQn5jz+/j11d0JJ9VK5M9
zwl2s8QKEFnPZxFB6YMAdW5kw/LBxLHFbf97IwGCliuC1ee/nqg2VwQ9gISl2dvTsRGS+8rAYHyG
jlwsp64v9SdQilSICvw+tdscsbRw34u7RtL2HOlWXYxsZnQ9jnhGDnSNd8ZdwpPICl5ccQZgV+Lb
hsCAoDZTVQNx30RnE1nPWTjFRQfp0SeDGJHRJTD980Tt1GDRYAqaErOpwT1GvPlr6dn0HRYCstIZ
aPtvp1yK4BoHEiznXStpgWYJ1MNkcAn1+ZxMTpWsa7otoxLuXvm7U/llAboD+nnbo8fIJPEnU+/9
gXFGgktJRCc7Fem4IRxEY/LU4JHc+ORN/NyCchHyW1EkVxkI2jk7dP8mq7g9yRZKlpymqWtDGKkZ
JsXyCRA7nZYMte/hHPWYXtYWuanPV69ep5PdiMzwfYT9fIsmRWUjT51ekOVafinhJ2CZ//xfEzR3
uBDCiRetDWoeEOpj0MyDINpJEJEF/tP6o6r9/uPLsDQl+qxDunWfrYdRafGe2bACzBifxIl9P9wi
0ZUJBvAZeNRFAdTnnOKlkG2U7/wpdWAzusNxcFq+DBUx3RhvuBg9yVoy5Q53m9rm77ak9IYXQhDc
MSMq0sb6VXzQFWSALNKCiGtE5fhbE/Gl7zMrNpqBrdCq4dEYHCqbQTfczyuTFSpkQ7DXbf1i9v7P
Uemw4vypBJTq5RxecxjsOMi912kgn81wM290s31oqpQ7yycgFAQ/MNOI6UhUYyKSVfe7MLvXkIo0
fNQYq9BulCoDtl0Gl1s9tspNq1K7rirh3TFMedEY+7BTotSu8wEbFFHR6BNg17cBccWR4/Me86J+
ZwY5m2O1kXz+vyMFd/V//PLh9Z+jZf/bxnTSPHGg14g8eekvKUQ5xxnfhGNat0NzcCE/4BoRcIU1
ntzgs7KeEtEpwDe6AH7IcXsCOFxjjEsVNk5dfWtlYOn8KtgCSiSbuDWWL3x108xToJTGZZtYTtuT
RdqhlY7CTlPPZQm0YHEdMKNex6UJEXR8eMy7cWFLnxtXKYUNfI2ZalPM6kGCOaXBkCrFGKxghzpg
fJ5RZvXnLLU2Nv989fO9CYlBL2myW2re1Kb4W27RBtzHNInAxLp5aScXz6gp+GxoJl15RO+tvbHT
UqKYMAuhDpA5zrSgifCU2Uy90rhtdCnJ3QTWUuzoyqmnOfpWFI2vrQBdSSTsiwKdz+2T01h8J+/y
dkZUkQ3dYR4EtkHV+BBurGwSEnZpDFc4ucvOYpYLylB0ylgDlCEhdzS9eAEGIL47utlp+5tBpSE+
wWFFh0kQzPSz8rX1TYv387UEj3+W0GO6LUdxBK7/GM3szRfNn6XI/l9Y0lzIefFfMSq1trC7Cc6o
0O+4xGbCUgVUZRBJ81RxlPh7paL9MXjT6kFpJv309xGx4qRhJwmRfo2uAXqdJEjMUSFiNHJItzSu
jcRsSvgVHXCUUptRayBJImm2JoQO+01YarzG6AxJwko4LdJDfTa7M4hrZqYzI7M3ZveeFUOcMzEI
h++HNl/hm9sK+jYnrcEcxAp3lh9PXGHbXEwVl7sMKUPRrmrqribsMd00unJwLJXdstwd9buTevMo
46mK3sWEP4Q5z09dLHQYtfngZAComVJ3kxhSP8Zaw+y4sz48kMb+gd1AdwVuTVn2tJU2yMYv+yEj
fCYfvIa8o2KPRqxkn4LZcTO+tBEqEI44tcY29vCqjW2mr+SDfZqNeeqlmBNkPBG8Cw25v4Etzt+h
0ncHJ2OlLEnptm+gTulwCex/F5qHl/bQ8C6FsjQZMd7clik7+eAuG5ZtGKAEhjNejGyP+CirCl1E
mkMtqO5ggVxKQqEJf6IcpZrZ5N8CDLDW4HCi9iLP1wta6kGgJsJfkGFdxYGkbaxKf5s7/HGglIu4
K1VUv7LlIpSPYwI698peZly87cKRgGuznikLQceZ1PbeEDvbeRflioWAWJAlRjmuiUz2Vc8vS5a1
AtQ9s9DI5nsrzfMRQgRlnOfaqoR9fgyrx0BGKtOxOEWIQX4+yGoB8O+h6dlg8bJMk2cSHy6lsZMr
xaDU2CZUueJNrKJF7UAhjTXyaDCTzKVLg2J3fsxjUNp1XbFtHizQ9WlGwFfFzYJj3Qisg65LgAZT
YgCq/DHnmg9Gm4pkL18PU6PqW2Pn+iTMrHR4lBgZje/5DTd16zugwxOk3+dKK0FDryJv4TmHkX+3
kcTVZiCotlSiSTwY9oV2/S+ThoQDINF0Qe+TLlOVkhmLCj4YAHmfqVIQcZV34evjkYPN9Fzg1AwM
8IyoXDzSF4tU5W3BxOfnQRtpBlffKKs83J+uXHzURDan8RxZeJ5qDX8hkIFcZKjYO+a4LQtMUffD
hOCzpk8Gv7mtpDJfYFlBbOviYXWJ9070DsBYW4sDOz5gmvDvELbdtAWKFC1qmdPXkjgSd5tOB7nk
0BXUsElHSjX2k0VpDmYxmUQLwWOmpFAOTkAYsmV2uXKLZrPZGuPnzBhqf3SRXiMxg7SDGbVCprCL
lHpjCDmT6wLhjXbdtq7NAv+butxeoqjUh0mLHRyQRTUTBfph7q0MgzfDFIdBmX5E4TgGgOOvDpgx
yr6hx5MqqqiRM7QDKcMj8WzBfoRyjmSJoSFANDtsSOwr2R0Or8Q+ReEF+TWZfaQsXRBqn+DZKKjb
pNClzM0r4Uro36qgK1e3dk+m+JQBUl/F3S0MmY46NyV2hEPssL9R3rM+3hcNwENSpUfJ3Ok/DM6w
abvGs7yi+nAJdQ6jzTGM18m37h2Ra38LWRLcQtTsN5342ieSOgTDjvovv/jC0c3EV3EC87Z+2/+f
5PlzulP7SAmPOJ/cSMVAJ5ERseXCecXucWi4KsjYR5L/rEKsc4hnh43iHjhOpHAO1PNW9pBpBSbe
vZh5Vs35CbRxAtKvG+lNaTGm1DrULAR3yuDZ+M+a4uJfWi+fVbEhbjcaEtbz9oYHAPcugYGsxTjO
VuokWrdFWh96mcW/tocXe5s6e4483ipPC8YP/iIZWkulR0fRCAYuKRI6Ct55VResd17Fj6/+Ihlc
pcdZU4B4lWZH68YFtO4pF6HyfcH1RRyB5eCq/Cnd/b+oJDvHekdk1cnpIrDYDBmDJhfdZ2xv6HPl
fNWA3NSjIQOGemMGFbU+XIPc47va2bUkRA+hlIxZUiEtV4+4dJ8Ys6/uQsM0wQBGogM3U14Xzs/T
r7/W0iIi+3WsrGOdi9+X4AcJVxC9uy1p6OPGPgwye0fg8hWFoKvxjOr5ea7xt49xcijdxNBlJSRj
5Gr1lYOqpctzR1Ierb7UIxfigV6+YGAkPCtIz0be765c0lPWVMSb7N4F2jOwwvVkWHz2qL2PdDjR
CyU/abFDImbFCfse0fs9EJupAcaLXdUGn7hHqtSAmh77+GgoT/BzVv2xYQZnZT2zl3cAs2lsTMG0
3yj+w2zlX2xhW3S/+Ucen6EgxDVqy8gY/gZfaKAJrGBFPfGqoBGbFFEFww+dJZxveiVWlFYMrcfO
XEMxe/zPBzGEkP0bOkzh6zRWdOEPNggFMs4CBPx/LGpdoHOBC4BcvtpJYypigM6qFa4qQMw+w4s0
Gs7rrMhFbCyoQPl4vPDaP26yxMk+nzpSIyesCoPum6wvhkqBTBE8fRKSM2VsqxtxeOVe3kz+9KT0
5bisD82o8dB9JgpL3MlW7kqrhX9y82uuH2rP6pAAM6DbcRH/GAqGK9X5no/FOUGCCqcXRKzpW4Cm
maNMxRT4TOz7pCZKhmPr9fxrRH88uRoPCBF/4kc2FfO4h1obk3ZpM7KrRC1BEPDBimjs41vsZqeH
Xfo7Y3U6Xg9+/SaeYU956pQCPSw1DtPY8j+HZzb4VP7K1FsPtLPym5Vb2TQUBhxHFQQveIJjs7Ny
TStRgOKB52u58v3aPYA9EXR+hv7oJtGLM8iIWGAhfLnMeQcj6zzD+Iki4LUfhlO2QAukeycCDFud
/HLKz7O3Ozg1Ly6or4Qno+Pp4qDMxEp8Y/lShEVP/pznV4H8qmOB0TyY7Nk3BgxugJCHQTcW6jDf
PT25U7yPfCwMD+DPxvcBv0It6NzfkfBsXxC0I0XvjoyBvsHxu+JUoE6wXGu/dhJekLXkr4iw2t6I
zyu3qByEmbhEMIANB+jyhQ/SkZMcqO4760jlZwwiAbbqzdVqdEBfz4VRYj9bf9mTAmiycC9sL9Gw
/fCbA3AxFPoCy6JATWYoc/QuNTTXbJMDkeAWtSeV5YsuQQxeQwaSYsnhfgssa1XG2/4tg4zoBoWl
XEL/mgOMH92Q+YT+7vu41cmGzC9iLn5b6u/R2ED53j0g0qJoOADhi5aH8sI9LGxxVmOOTJ19KvRe
0IluFZ0LKmV5QbaTLxELrXJ0oxuuYbFG6isS4EHTEem8kPp9vKbUdlUMsBW9PGW1XXksLkjZhfip
QIvT8yPWdw3SGPjxq2IwHKjOBuMamZBqQlb2D8uUD7sP9jd9iPOfg3nwQAQG6ZKSWWzNqmvx+1tB
YeCy7/IsxnHhbkPwn887gRRkcoI6esN6l3Hdrq5Iq9t7febmBHTWLuBfeBSMbiGhvfcdBDChzcX3
mkA2D+vcDv5CKt58Pa+DDaUyAv1TIJqks50CDWkA+jrACxWmzi8I7qM1+ir3k+MeycuACBjTA3/I
+7w88GU0WQLgIsZbJl6MmfOio63+4HwNNOT1BeU/+aYEiA+qc3qPglaMk64JXPpRzY0MUdynE1om
GOXEbrgHhdw68hFhLgCpVYPM5lqviH5nN6USvJN+BMmnm4znm8M3pMmppXm5YsLcXmULSwfKGYtE
jJTojezEBbMGBl0xUAlhdxwkJHT6biQL6XOU33lUwXc2gVvVNgmmGOojMfrypXyyfcK00+zABM1V
ghaTIhUmZGeGWS22UuaosRtPqSyVhcvhBQyv7OZz1oU8/445R9GrozUEH5sT1dtcOQ0mgmgIVTAE
MALxvWIdAIKCan3WRAhDXFVNewliK2TQ5ZWcPK5nnrQJahUWmsXhlvepTHlwdlo4naska/MBPZa3
L4RRz1123SXQycf2raVAwoTQ6uYvWvu4qMOtjQ2Q8A5S5t73NVXzqhWWMgthmQEcpExRPvHelQVy
ENE5uJgHveK7OIugjvjc7ANDl+V5KtkQmdMfe9UDBANpIHnWpdCf1in0kxwtB6aks71ZUyAJCYnL
Yp3y9iJkmYT4+eoLtESOqcFwr6Q6MGsQBQx4/9TUicjeLtNDpEVdN464ZwsB8ODNq0ZoOoJ4fTW6
+C1o2A==
`pragma protect end_protected
