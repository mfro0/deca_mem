// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:05 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NaqYpHfP24uhjs/7EW3o9GJKwkLV6tWvaye8iCSGKmfpTZ0IkGFtJ0CRqc0Ge3ts
I8ovGwWKQD74M0l2brrSJ6515Tsqag4knP81dsdQ3hRXX/RhXzVE7ofRvzqZkG1X
cwrPJ5wXlDlSbMSTVdGzo27zAdgaoE9HYSYjqeh91Fs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11184)
WIWDbq/1lOFnnc19LTEy7IGCfY/3eSw8Kl8Pe03awDGhHzab5oa1vxK3TUp3dKG8
HDyp/zM6uacZMGOf6IhRASNVIcZl/pNDZhXqjtg+6UQSu/HvtxC+i6T1GUImdMtt
2pkzw/oIPUdESW/FfYVQx1cnYEa1EppYyzHxXBPhd0xFpKNSiWAoQCTgA6dvQgaK
IliMD78LejOvqBPzyr2UhEAc5qY1/hvdK9PQAtrvEiSEWTiO0XJBO/a2yvEDFWxT
NRCJq7+4I94D4SbtAoavCgmTIQ4QYQ3jEsiEmuISMKLvYGwihVHY3jB0GfuGZELj
aDgaNmiMlgUy7ZdOMLd8EcfdBNAnKiJ0GmP+fWjsMKwNmjDJ6kdIBqRPrXJctvZV
lpQoIPG09+fHUIxHarE9i5gWAQjflsoWv575VmDqDBpdS3q7QVGU4il7eqYkZt+8
oHU2Tb4D8Rz6cS7FkJ+HfQh65dG3OrvtpKe1ENH6ODkLrR4DG3785XFKrVQ28dxl
vp0H/Jh7Q0UMt075HNdZkPiQBZ3K1eDjQkL6DAtw2AQmjEhJDejMHR7YtM4PWSg8
ppWza79ejDkPsiyan//qlHZXuHnx6mskhyBzpx88GcM03ofN4JymOhzrcR+ooPVe
ffBX1NLEV+xOmtOT483Ox8ETWc4bBe68z7aqwLunaZiX6475EWxyQ2UErg1ZipwS
GgVfPxZ2FQHvBGY+yaASYW+G5AqCmf1pOBB75jqDgJ64lcXQhDa0yg/EDryiP15/
Siujw6LeKw76HX2EQfZZpxUl95NqZ6kt0cJub9jn942XuBi3iYBxFp+L4vc1RBk4
j3O+nfjpkFfTHX0/5tnnIA6UpEeRj73Qh7QxwGBGsIuoQF/0bp5fygj7H8lJrOFK
FF/2EYUsaEDdfuTOcfRU3mj8pNpeZeCI91zSK6Q393hIUae9mtzPgXy2C3Slj1q/
GIWVPQ951EQbhtHwh7xvzjy64t5JS86DR2ISDIqWxEELDCab1k8joYosjfbxTC5k
QP+HUgyjLpzIDO8aNOYuOkDAtTtJRiI7EjGnPcTuqoT6a56vhQyD8KUDXrJmQfsU
tCgZlIjBqA+qX7qLEuvDwE9uSn5z7aghke0+5HfzcPixHfYF/vEHL1Aade3jT2wJ
wlOk3N/N9OLp+ne2RIW2saOjtJsyp9Wl/qbWmKHn9l/yH48jhvR3xtPB5uL7RFrY
HCNChEst6bsSU8f6TXmkdWVKGb5FcJn6nJ805zLInQtPmYQOXmfbensxjAMwk7xb
7e5BazVyrPOfp9zReiYIQ+v2ETEgcFiQLEL1WrDntOu2YBhFEKtE2K3vxSjZssn1
+L7ADGFxx0QoRbATPIoBud9Tv6NGo0uvm1O4FOFJo9nJEshLnFKVmMOpuzO1Dr/7
ZasYbb7gYVD2ben3lF/BWW/EMPa8OCD1kAMgEl7eIqUZA9RLALaGhg+kEEUCtx6z
oh43gmmh3n3DAMHxZp5wiS0v3QtOUqlvc5xfu1RSLozPCk7OeGjonMzmyjh2WO9s
NnxKskKSC/TWtkCJWkm91LMEaeix7zIrKbourf1qLTcBo9JO1AUfHoeFKQf9Vkv2
1plu6JL9Sih3Ae1Ia0QCtmXBPdsMQqV+VaDEZIJXoLtClDxfAzkxMS98tcOa7m9q
K+z2/YswT4ZSLToDtXmzKd24nwtj4VmMtLR2vT6ZxLYP9gC97ENjfJl3+quOKv//
qsjKfLvplP3OcuU22uN7aNlad5i9wTfkcKfPjCa3758qEtyT3zqDCvDyn5xa3Zx7
eO6fOPJcZPNOsY3C0VPZnOkG+stDW62u/eWKY3RBpW6fIX4YLZpzh4MgspPKXpq+
mZAA8bsHdYfLgWQW56rh+/XJfbx2RDbe23nFb3GFVWQBv309Uopt6RbboV6NCVhj
zelUO01vZ0r/aC8y4k3tBl/RevRihePWObNgOoZRYChOVaGftHfKgEZkJuQkdk1a
tdgV+U9qt4yDsETrrNkmUwDBGHMg8qE0JNnHVbdgIIhWYBvk4yCyd7D2QazuMfv9
u0HuvNHkgiU/V527toI7cPOhnSm18epPtKPvsDmRQh7x58wGA3yOyo4boHptjqZ5
4tFhFm3vQfRAjY2lhU0xoR06XDy6p5YsoZo4Ep1iErPrM1EpNAF78I/XN13lOp6W
IFaMNGViNUX5HMaPjEXmHuCp5PmiAs25q3ex33q0A+88ZSS1PMHSfFK48X7IOnmz
6JwxVbuPUszUyRQ620gWiKY3st6UExwaHTQn/+iOdRATufzjuT9p7JcoKAgho4y/
8Z39pC/8qBb9fyAKQ22JRFEiUx4dI0UUqzPGEFw4Wj8agXz/8i8YO6Vos//x8omx
W+Ic/yHf4TqMi8Sv1pxp7HAAhCgeMaLylW85UizWVSIMH3m3IjDwyj7BVUAldBls
U9Uha/3H7P+v5FlNRLoid+H2+/tLvB1of9Q+WpWZfFuGS19Z0pycQiZ8MPf0rn07
/F/T08ezsFrni2p52icITk2Aa0cpgY86Shj3SuSzXUlxFJ/kGC/rCLKTmNu6XW65
apY5+OTW0GoWhcyNfsyeAGS5a9G3YZOaahSVHAahuCuM6deNW3xd6bL9Wr119H4i
6Grh6q2k8qZeMxG5ZB66Aa6/5eB7XxX5R/GDRm5bk7EPODvO7ouy0GQfdIAZ1sBO
UyzmX/ZfQ9G3Oe3kgTvWykMQxLBaIDuP9llVOh4gEWlSwjAVJ7KvxxVO+JQIfIN3
t7q0hLS6TSkziN76G9hB/V3ov+XEfeVwuluojg8cRjbBW0Mfcsoi78hRKqFlLWj3
k1kK2RgIYAQ9sfLJu7/4uG8wwM5SVx6CSuaBbQN90K8o/Dv5IVwPf0qxZtEAclB+
CYTf0W5dQEGTlPbBSAoVx2oovairUjbWttx0gDtRiZymMHyXqilaoSXTmp8H3pF/
tu5ej7ZX0J8PTNqxA1da6TVqKuUe1HbdikEg2nsmMTTnJeyM4NEVaeUDtNl3hwMC
wmGOr2FpIBbarQ/SZINShMFGRnQt3B0Up7yHK8Bgb5PjDv4Dad+TrdRVwBJBfItM
xxfeNq6HMHcWLXJ997LyKktPQq+GIS+ZbPrCt4NI/Wd2U+F7h3RP+tE4TK4dLaHS
Zkm46J/mzMoqy1R3fOSTsRtT3TUQW3MVqEmMc/c2S/9fn+ZYO1HNBEC3VPRMcA+l
9XfR4YSnTIYwhNnBbTK30fAFICeY+3Rrl1atBsGxaDPXq/0XLYAJ4xs+QJnnYROw
xhOHFtRDma+6G2mc7H5+vBOuSxwzhhjVy0QRpyU1i+hapyhcXnh1XtNeXtpHEnwN
wEC/svTqGwtHoNgTTwzjb04zads9gTr8sKJ3/SnpMOlMx7V0AMSv9Jxb/aYebh+C
xbFc7ajcBBxSAOAow5pJdIuyBo1A5U+31crKKwgvZ8To4eJ/Hc/5HBWnQMF5sGAW
ERdyAGGPfieAq/Iy+LJP6DmCd0DQqoqH6Yy7zeud62AyKJPxxAus6NbSL7UI/g6V
hSr87IkMb8OReeKTZ0Vrp7Xlz69ssGpO94ADgGkWJc8nexKXxVTdUx63AIflIlPJ
vBbO4Mn3leU8yl3IoghkShoSd6ci2c7ece4eqZ3enYTfhzrQH27rRQoDFowy3Tnp
JBOnEgHHDC7wucO/IbpIEMdbwHNS/KNqeq1PMNQQ3reVUgNXmRJqPKm2UjtGFCe7
VOFmJfRfVb4nZJO3e0tsdNsmhssYtW6WSHFyNM67ttgpOOJf4zSJkr1WCleoMgNd
5SkfQk7Y1wzrqeTm8WcIAl5UJR9PX46S9VJLMGn6C/p327/ilkwJSL2BrRQWL5nM
wXbNfwoGMMkAIJeP4ajwaBQw+GsvDk0F2wiwc6kZltzBzk3EBASSalX5OeU/VKZa
QC+fgZfeVhCCG9biFgdtQPdSchH96qJoidEeGhTn9Ux4Ef3ayV6tRUopeP3JIo5a
i4YBK4uV+Qg2MCbq7x7xeax7Fpc51VoBFQGbvzEvwWqQvTdGCWCHwfiLzOKCrxe7
Fw3VNPSmtxHnvILeQj2bQT0GPZSYD2AVV37BMi3vT0t7rHckdgz2Xhz3csokU6YG
1m/1qvfWawcRlO6t3gwONodg0d5M0w7aeB5mL0eKc50aa1U5IYBDVh2feB1GxAyd
G+upCljzimSuxZK43z0QK8qWTj+o+ODEuKIefOYjhin195xDN5qDHJqczSN4KY87
Iu0lSPLnml6x8bvW/yOhc3S94H+KBoPzN5bNMY9WzB1UND1o0Xz26mgQiEL3RgPC
NdruoJ6ALOyYymMpb8u9DQh4e9Z0y6D/gAXPfm7h2PRhCtmpmg0HZfM0FMwmMs8g
kv/yBK48o4EE6eCtaY+CLd3FldQfIlPdEQhqIOAnQMNbHeM/WKrQm8B7mpNqtuS+
7t/3+/n74TCp5QzNBKkED7KEWP9X97rbkQ1WZ6W6p+GYVDGiifA1imtrP+mpz+kg
UhRY6zLgsx+ABQ7vYxjs+lSIuZ7dExqewY0QXejanam4pWyeTVXQaBDPGYO9EZDM
802syYu36Nx9AeE8nIegEso3CC4NEHtZAam0Lmak8sWz8QWb8eIeuia7krnobjAU
cBIdVGPmUqR0tpWdironDexuENkPZIRU3ENaWB9KcNmA5OSDZSjKUS/R1mZ/UsQZ
vylmkPuDrRfBBIEjV7sSBnDFBB9GvKXn9OImoODbI9n5Ys1YAAXVDPfVtlkpmAIj
hu0SlnkUjUW4Db029ZEW/eTbZloB4/RfSdeT0O99t20z0+n3SwzmVfGetyowLSb6
eJQHJfvOKFSGO5m45Qa8WbVYxUDwoTwrgEw3UsDhPINyRVHIOONIx2Mc55RhxOyw
NIED3NWiVjcF3Q9ZTeFsL3SU3Fx2MqOgYogWYbPyJlsUvtvlciD6M9HgbbW+59GT
BLMaB8ZXyGp4aT3Vn1Fkr4dmfXNDnuZGo3dYBf2VBc5FAi/HkbJ77sHhAEv4R+GG
CHnyTBbnpP+J6VXL759tHcKlGFReqGSG+63WzXzpNUeO8US7tk4k+phIe42J2V1u
QaIpwPIjBO5GWQsN9kdacjsxd5v1A5/sTnYjpRRXNCxu+6Cq3so6+1/FW6ej8S6W
o3KC2pQq2CSwpGh8TUVsnrgxXDHHwAyQKMTUuFJflov/mQvuS9jZ2aXkXJ2hB+qY
jE+eyn+vAoArPfwKdRZxdHeIsiRI/Ot6qEdOaP14i/Miebkh4Qq2Y7LBqWKi66AH
H3i1B/gQyihMdWSR4YYMfaqEc/gpger1RPfhupDPmKsD/sKJ2wj65eXJ5Zr3+kjA
3yeAzvaMXu4sYGJgxIf4meh4o0bIeUgk0Yp6FZYIS4toRalVxCRrm0LGIeQTUvcs
ekjRSGPFMTR035FY9sV+TJkh2VKCaBPhM90NJia7DJbFh2v5rvDQN55t6DsWNd0U
ThpjlejV3PUHAquOk9pVe+0c6TcZ0L0du8IRQz8LbpXnSB1DDS/PK8QisKE3KVR8
0DpwFD+xSyKwZLXE6HnOhuwD6LgkCf2XxHgY8A4g29Db3Ui5L6j1jxLkbNgkmDMI
E3FDd9tovZ2AOsfUfWAbKR9UF1vj9yN5aJ7waR48zpsktK2E3DUvrCqRT71NbhXl
+vrvBt631cDyXohGUNbWmXM0HLoEYmB0NwTp106XyjA/C3Hj8D5c8khzA6c4VEOI
JilgnSeCqyJn6E8qQrgE31aA6p893vAoDKtH2dmzQ9mUTYFpfd7aGUUDigczr7J5
1p41IRUSZtJtpuesOC3Ll+9EBqGLRZPN4nnytsXP0ntG1AKYJAY0Tom+I1K5CMmn
PlcQd2l4rKdi9rg8pNBZGchvNH2IX15zL7N+2LDe+J8hcixY3gzEgNt7UFS8O348
hCmcbQpAlo92U3BXH6yR6zjfrnIrLVFm0DxMcRx2EPdU5hwYclF3eM4RLcF4ADTD
efmlRmVg6/cOfVczxqszX9Pvs10n56yXJAZdCXEjTuCaQ+CqY72AUpzhgVs1JuFR
Oe+EX9Ox1BBA09nQpaNI5F2MCE+b36S/zAmOt/2zqNJixtYsd05Fae6uKX0L2H7e
rgZaBfzfQ8GlH6tSrebLsLF9o4nYkjML5jT5eVAODq6AosLjsyPxUMW/ACjnOrKH
8bhXm8DuRDwqH0pCmX82WppokSxfrTSPSgQNYyr+C7Jpjigop+k8kzwDTmnS2Sz2
m+97lQVP8prrva9I2tPnRxHPSoyU7r9hQEY33/8aLreDskNPrHYkbacxFdgdhKS6
bnPTM/UIMxo8a+NQ88kOTW8bBDcQnxV3OdWBoleEEJQ30lWa5Fu5GpLTJtk/uNFa
R07QaDgngRK2uFmE+xrCfWxN1F+EIXatIfYSzIknm1sIqvFn9nwaoygHD7p4NhLJ
AaiRutuTkcktMdd6iBZcGq2VkOcuaIl8MeQbfQxbsOm+cMXjP4uVSf0TiyB+otPs
J8g3qoaYHj0i4K0HFuPDgJiL02CFfPr4OID2b9FKHkNtSc/UwnZkMbjiz0b8UXju
b3p/NDP7k63AnQWEUmcTLNSFj8q2zEXizEGNuoD1uuEWopM3v2WJVj1xjz11HVh5
pbUP9dSyuUUzENHtxMzWGnA9Hc0n59fm3ZLeILW+PxTl9MXSY3NH5Fty7g2bR/Eu
JVvLa1zZYbaEC2CrCAktbAmXtH3b/Z33+KNdUjPNj8xyn/dR+UsvVKm63d29aErk
m80bUibhY6cVewv8xCvMPEQGBPDF8Goe0hNgbdemgOYk0pDqjcKx4cVooDICwmRx
tDbcnEgHq2IbI2r7S5xUphORAVvlZEdSlyojrDZmGaGKWDexpduoxTwppszFz0A7
j/9+j5l5CpOtNElqJrZ3HTwqKgxErRqTbUgQLduEuo9Iu1hrqBJQOENzBLEs2YeF
r2hQZ3j3EvHnTQ8rQMhcSLZiLfPXBTbXluJTJUypQERjkHepww6V/I0HgPaJYXxB
pWk8h9u3VJj1yyuQDu+OGjOT4G43lH0p/HUwwfpZaKhN3lN7OnJIOO+UX6KwxZMz
Pd1fIChytKJUFES6IQ9DzBtasgKoAiCsmBCzzTBpCNASzxihPyWKybb5LduIrTg9
U8sNs9FgZn10ETRanamPIbWqmY/gwK/kQnWLfBrAAOvf5AE46if23znee7An/NDH
h2+H5N7KiPkm1a/YRGgaAN2VARC89SqaEjQfWz4jhw3jdwFYdDevstmtVvUJ+f7O
iiEl9CBuzN4u+4/FlNagG25bg76mpSXyir//TafmC+fR7KPMhMEXifDrbL6jbKCp
+jF3T8v4PRmRvbDyUSHLSlD6zJ9mAIsMlxcSRPzsEQw1ZacZZqTMaJDhUcUgaPVg
71Z5U0FWU4Lj9m+FmKEzkrVZW6YY1yEVJZo1xVnZdrPjZLkMkOltlcNb7XKXANF4
EAUeoHJk94655dz2RW0yY6inkffmeno3jg1WZHzwM+rn7WLGzJcdTpXCmfnz6CUg
D4m5EIVUU7r9o6zVWELpceOS0dqgBTjVIhsNAywAZMaw2mK10Y/d1G/DROuEWbf3
rMEAce+Amnbb/NEhQY1h+InR/5czyMtzqW0ETOnVpVCRbWhzvy19QKRDlWdYF1fH
ezq8zqNahFHxY+ovgiZ70TA9zSQwJoI2pfUouLTmeeG1V0FtYTtg605TFMjj6kPG
IpdLClkOxVOh7lroi9MNXTUtwyoFJGv5tF1IW/e+ZugfN+11tCWFNPUq0jyVPEya
663+iHP++Tgb73IMA/mV1pWpyASDsEMJczJnQdRZFsq1F3F/Vl4qlWknYK+aMALn
HSmy9pmxGrMaqhAgTHa3PehlHUXZ/outc01w6HmPgrDx5vxQSQKyVDiAkdmrezMC
VCBpIHbSSo6BeOpOq39tpIzGvxlFjOnDWDnfWhetcKasehdbTDbt32SrfuFUM9rq
Ww85mrWGeH/9nOO7BY+gWdXSBhCrjjC9zcbIdFLDcQ+2kwo4HsNheznhAV2HVEZ2
7wNzuurCUeguYBiqHvcHJE7pc3Hq3QFQaV0Chs8ChYGJLxMMuvE0LvaKd+km0nzd
qaCu7ZIqeCeBtzXPP17QWYGE+wNNULa+O914opa5ahbEr/RcQXSFLO61EArA/Q4B
JhxLM34vc9hFbFpfyaooFiEiKX/ErrycmdmJmiMvAt6+lySFXnw8nllUHqe3pooq
oVm63rn6kvvoDkEOhXQFjIbanshuf1CEBQCjPDe2xz9bsb46YgZQgLNt4V0saMl1
KLhAG7Cjbasd1BfAi5M6kCnOMtlB6ixG89N8j6+PfWDTfenVRGPpukHmgNVsXIob
0jz4P0oulnaNBrFq/kwvcjCA86KKWpYOphER9v6jsZOSD5OWfGpKLb45zHAH5MTH
WJW8kvhpbYerkG/5Y06us0mR/x9p9Ia4WUSIjpwn5nnB3JVeaFMj4CiL5bIOoMmO
mTDoh5KqoUaVPL26IKJjgnryop0nRQ36qlT3fmP+fNPebnbf61qFSQp1kEsYWjAx
cx181VVjPsP2ZF5y5D+MRJItRAvijodSml12EW1X1f75Nzcpl37Fx4mP4tCERabL
ZIJSNIqqeV5uX9bZkk4jLx4If3ARw1fLB1vowuWdkDCagjR/1lhcySBp64I4wFBR
Eq+DB3jnyzCY8F6GvzBXouu1KQMaoHjxjPMrIJZOURvF8pw3ogQ8Q5aA2Y+zkuQ7
LQCARLU3LWcSLi6SNsipm3V8BTjYVLV2xjC0doYuys90Lws24ZxDSCTwysWcbHPv
c/Q8YngErZxfonux9FuxFxaDc7gROL9T1f2pdt//H26CAHwcrWnAybC7I/sIjJwA
yYG0oMljMkXIDD+RPmOsolUo+6Ws2qrHGPlnrrUr/WPGnWCdI1I3vVPtKb+3+VOQ
xpGO/Cp9ciYzYc5n/0zWAd/8JLW8TxRnDN8qdeV6/+FLVJusStqdQqpH0XM3Y+hx
sfC+pMJezNMVYc+kZBy/cb2+1BpP6K4kRG323nXnnzvNsNB2EJxbhlJJ+cbJXK+m
VVYQ0RxVINp9fTPpfXezOv8Idsyump0hXsy0Q6GX+Mc0vMvcYV+fLxoH0rTVVAia
Wqrqpjwofo82u0SRAhYk/6ajxqdnbuo6eR5bnFa5Iy9lEW1ao/Si3JF+KES5kHDF
SDu3NnUolRKmsHx68ypJ3eifogItUx6QaSUQXVY9irZiCWThPBQIjy3AvY4mf0tC
KBNFZGIUOQHMHwK9xHGbP5lX3k9Dvan2EM5nSG6WVTcycdALXMOz1nGmFsl91/Q5
xWNvyZj4+uM3pPuqqBYwg1/vpgeslTb7b2ClP0XpThdYk9C/dANRmkZWSYB6lP/c
1eK6Br0izXfTXn2841LdAlde4N3BjnfLxp6LZ3SYsgxp6hT5lQblbGc33JHOkswp
4keGZoc0xWVTPPHXBlGaoApAIiMlMsmgsesuegMeYUG8Xzsg/mgTYJg/i6OuwadR
0fNrBWgzNB+eIaGH73nEfdhT8rnnKU7gmtGcm2pqHg8+pENZsANkkHqlribnfLW8
q5zUrqwnR8/NnrkAnEWgkHah2mfEGsJLs0WnYACbkX9yFnGBi3QEMz3aAFHfSlC/
2ALxDeJFiPR02YoazOAS81bX7TtDLL3nN88reuCsjmQ5uZSsnmFI8wuqXlurZnlN
wbVO+raIeAvHPVFo4v4tvPwMxwJpruMpJF+M5ej6jG1QcHF6mybzicD0DfVur3eT
S4O6EQiJezll5NRx5k06Yegjfd8++qUr4VUVyuWI+RjhByfyASF6xqKuh3EqZoVb
usT/XpwFuge7qS34e5a4hEPP4OS04Ea30naL8NbiK3rY0qXxippC3EukGitJjWnV
eLOX3Zqm0HA7Ux4i5L4ZOmOuyEXBZD7FERlgyECf97JgnhU1ANBkCFZh2/5eslLX
qC3FhBRQsHLIElVwS3k6727sWRewCjvyY2b2yhucykSbXFn4aas4QY6jfzBwXewd
YMDpZeYRgiGhrCesptodZq0fV7CUumdXs1/LL5Q7ngEyZmMGeCMlstg5+3Ke4dw5
31zyMFG6VJckGlwNQcyvbX7+KOEJl9vhNbKgEnveXDkRGOgRe56mfyFfdW5ZJpaZ
Awt/2p+NpsSveTkILQyxsAu4L0FZABszVlHbyJB2Mq+6KWSnW0VRJ2fMvm/ht72Y
Kv3oxSWlwd4rS98elUWnXd+LG4iIyqbrDZnYmhZxKjvH7fg9egbceyOTuf4f95Vs
0qQGz4BxJPLQKH7LXw0Cmra5w/emfhvx8ID50H6RtHdjG5ymaycSBJHWmpkZHDTT
gkdkU45LT4BmsD/kBDdDx6vrLeZAnoX3facd32LPL37nBiRHEyr2zmQK2viJaVQR
1scxPiGSTeWqiiA2qHt8UA8nd6xsbZrHB+PX1TPP9OkAmezrDSbjdSLlBv4ZnQg+
0oc7EqsA1eeBaQbEb30sgdq1FQp/jPBSR2HJ4Le6anLeyiNrJs9OSz2THg0X0tcG
TNsX45mZfOOHOUvDYJmCle9In+6KccIo1QJbd05Dyl58skmz9cnrl+lBKEDW2zHJ
bhkuNAbwDhILCMNYz48RIgBu9RBGFCDwQN1/SGtGFrPHA1ODduAIeNXl65Na78Ar
8afxac395AZasGcwrq0jbq+AyL3PtTNZ0CY6fg7807kjjuCd4aNXn3UPer72Lpaa
ZqVyg3a+hepby17nu/YGByDRHDGY6AOMMNvLsPUxlXRO0ltkQ0Je9bQ/hvA8aHhL
w8sIR7c3xWHb5aarFyCvAtjM86f6fFls+PeKvwdlN7LwGd172mDDi02LuH0V2qem
pTn74iaBAjJrzFVCmaRwNzdok4xuLao1zyXs7GbUlv1xYSGpGXBTuAW0wSzRsqKl
T8GHGB7Xcv2tzaqz/42beLC57X0UxBVfes00QR/q4ZgisyNjf6EC7+Aaxlt4o1Rc
v1fd0KHcEonYdNRDQuX7jrZGBGkxEgnpQFPp2uVUJUIwku6VMNBA56d1yvw30FAt
zrIqKv0wlq9dNiQfTZQCJxSE/R034D8g/soRkbGOk53OVPQQ3+eMWWjCqXU4XAsj
410Qnbh8onsW+Tg8etZtFV77NYIURPMgyHVZBehSyeSxfAOV2LReuEsRBj2oWCq9
f1RYkpW7SJYFcvWJ0ybB5K6zbxmakSa495k8Ge9sOT7Xyzl/HvLK/ZE7xY4QwvsK
ahxI1jDrAdORySJ7nWJUqvpuw68YutudMFtJWE5c/8Lzs1acZMORqa9I9SVbfcYd
AYlBD2MbERmie9RagkPZKzx70bJt78s1I6BwqyVxK0WKqBF/kuKf2PtRSJED0Pmq
UtZ6HD/9GK8FShIT26D/OuqsGEtuxLfbTJ7Ua6mq6HndLFS4Fa29FDKdnvSpoHyu
Bff+AMGvUWmTUxTgLfzVkkeO0KEU+y06Ue9NYqy+TzonrFV2LUGErKcRbQOPQVU2
gVgDO1q3kgcFRASK10Ll2bh8nuSiwlAXTzXkb1OuFtEAnECXoLQ1BVyEKuBNuOz5
raH0NdJfPY8KIT3kU5qWXY8Wf56fkzXus3envWh3wZGybE2lt1fAkR1sl+TM/PMp
+dV8Giq6nzteOVYELzSchMaI4m3X5D+FIKHAyu3fzlTJFr9KJe/E/rPoh0ZUD0/R
l+72GiVWmW6q191C474w2yWXhmEnfvKsbV7vfhKqhLTBJ7wuObdpByiW6orfxJU4
Vnc5dUw91lPT3RYmNzhD2Nm9IlWksYFdlYqYoAUyQ/3FpoNd3XpuL/2S4eMHeZem
3yqTFLFg3zD9IUty5XW0I1aZxpuo/0KFtUkQfVt3qmNGZPT4p+LgOE6HUiGVbFKR
fft9t+U9MNXxY6wk/9/LtR6RXCtvbWoFiudl5QTIvhfBCYbGBOBkXUZwkPj4AiH1
j9lbX3j+NGKaeJ8c+/gYyH/PaqIR/Z+wX5s27eBqjh0Ftz1i1/9KmdhOmg4yqt8G
9CdVUgEn9cRmZhcP8bWuMN/6N18PqgwZ9B7vxBnuw3prttXf/+L/nRGxwkJqfK4e
WZsZGBLOmYC/vC71aE+0ccLQbOOtlvfmgajcJALE2mYbhP9g2ASqu8MgcjRAcfD/
c6GiiTrdsDNJ/RmipEFiSRLQqhPzVsTnmSWUF6faN7mULQDOhfx7L2GVpWCU39kp
nI6AD8R+rilsZnSB6/mta1dbts4MUnkZpa2Ju2ofv4ID7My7fxbB04XGLmapOGx8
E+M6NMp1Xrj1EbQWc9O43bkj6pc2ExXQ4CufRY0pYIhGd8s1Dq0Yuek1RtWJj3SV
7zvNQRk4sgjOY8gPldOg9FAY9gxzBBRo9ET7yQ4q476wU9jHg4mBKXBUZyeeYf9h
KKnLZBNnaB3W5wgx6ZuwzrU9IPsL+qTK/QHeODh2l3oxiWrbEJhqHxPAglLtFOWO
4MMiU2x0rgLkpbzWmiALdfVENx4eyTce8zgMIa1gTjVTsmL4H9FIwz/WIxMjJtSE
qmFi4qJ3WMR+WZEpDRIXZYFB5svJbYwiIA1IX8I5xrq3Cwr00+8MxApsSEaeUtjU
I7SeDnIsZJILf0AMNi7EVqNA/2JYME148cYFKzJTiL8Yux35QCwDUHBCeMmDnLKu
xT930QFyRskHasYUbQIHBV/50w0u3xWiHozDEx39NvkaTLbpYINUXuOEytUDub5s
LKbh6rZJxW+ejwChPPAScOWnwHzqP0gvYEKGGZzd/l+GAElfHf6Xo08hw76e/bY1
SHDwNaDXLf7h4VpKvmEq4i8GXPCc5PY7L43CyuDTXjUo2F2CWytaTZzQAaWdqOrW
/L6YI2/oLblF4x00UFGDfPaphuWLZYyL6OZqRkQsUvXf5+Ci05pykRcKj2VhFqQd
KEP2gUiNKdAZlWRgWeBnIdvWB4K5vhedJVEa654lpOoZWxwq2MvQzqX21Iv3fjYn
ZKVdvXqUlX/FHd+l3hPVKdjQS2HXFKobqOo9bwuR2Cdf+gREWSRn+fHKQPo1FTaG
yiIxllv4BBMzW6BK/OcbiwFJWN7QDlw9qzqkA2HHGwkAhfZMs7HW+Ey7b2QA9eJZ
aIWMcRNfOe7k1fAZJWfmL8EGZSF+csWFbcO/QX6QGg16+o25hIsv/D+0LaPRQ9qE
NF0NNWfhQnclYIJswv/bpTsnGNoNfXp0d0nYNkJf5xMEgy7jx31dOhM8mcvRtu/S
4/0aCZKQ32g1faFVCcOYjzw03RTwLiOcOZ9KMYd1NfBa1m+QaSxaOeRm7YQm4Scc
D6gZY9j/zbFt8scEmUJNQ3DMTGtFeyN84o91EcOpsfiB081aRSR8dvrIQgIKQgKV
ZrAIfEtAuo7km4OdQXP3i6OsuMhXeyPvAesA2SlO90MYzALC7uJaYbqMySLmep2J
yWUSk815gZ3GGe/Am334Olv5dLvLC2pje5t4XC2oOnjh02vDmxkuYnOVvfYOMCab
yNA0lYxSB2ntL9yn9+Je/jGcGlhI4t3blvo9K3fbfXPOHS3K3wz3cGYpOmyRjZbc
DeZvSXWIOPZ/wuULpmTrMGyvS2GNMUz2lsSqsWvkoMYBUzJhpoTPb+ZXQStWftWQ
fcFYPk/4Din17kkYFgpVsYugot4tT9P1Wt8OIUX3lA/LBT0l+7HjvGkXsluGjLMq
Kojnw9D85Wym5SRRYrFiB1ELUKFA6ZW9kRERS/Z5TY/XLJ9CHE4jKXgjVuZ2NWvg
hckT0RmyUAwA3+82I4ApQHGSLLoWr61Sy4nkNhtjBnTBv7xSYkvHcWJNW994f/Yd
2Lx5u1yq5qS2uxlvg9fg+0NcJUNYumXXbHpaKeRcH6/LWKMR31mG309PHikZXTYk
zkPsPqdCNGHeryIbFzvq1tZF91tY2ogtRtL8BltTGBkW33faG1FNyUrUXu/S+E/G
ZiXcA4Ua/8bZhMN6XEXxivZKGStR33wbMOgFH13DBiqyyN6Crs58oZ4s22le7/Hv
u7DnowZ6angINhJ/1h88xN5kIFTh4oAbmMaFh6aOkt6nTk+UDeUBy5UZ5hgQkdVc
pnuE8yca5NxJUhyqSYAqYxlo3ci8al72+8g2l0MLccahszr5SHYLADupJcEFfXTi
nza8G2+1Tl/o9E0Pmxj9lVva4cpfLid0GM5Kg3IptfHyPsJ7teD0vVpsaVX83n38
1TNJkbewEm2vHVmy9Ruo5oc+xaucxzo9xOOGFSYjpyigMmLmQHAvuDaLySfvrJC2
XswpAmRnmFyRApNgVKsc/VoWH1KJ1JhygMfy+Vo0nZYzKVYflkjx/5K/rvP7N5YF
OQz2hjVv0T3ksqr+qaaHAqwXsmHmT5Og3cLwh9geXd35mmGTJrMDfhMs3KFIxdvt
5lzv7KBVclBy0dRlRLDgEpEieW/K5ntwyB5VgC5vio7Xsce+85Nz4wf/ANzdGD0h
Ya7xHs7dKfMUL98jECVCwxldz2OMtma7MGvp1p+587WqPFsmaLMvKC+syPw8fqyv
dHiuvOWMwAbgMSnT/16O8zPO5PAQWDxKCwyVH76EZ32Ivz5sWHRUEhUi2k9lZ49y
krvrxtUSgze8msKJgbJiu+bvnddsXyGwsMSGrbykuUoSvCfa7lxRDEROn/MpaZ8R
Gm9J7XbEFbs1MI2s5saj8pO9KK8V7dCCPt6aJfJ+joXYekxWpUmYR3xkzY0W2AZG
urVet+eIC+iJbOGQfolRHl1hUoBUYPAFxIcoTflF8uY4W43yC6mHsZNi4GVuMJsA
FAE8TCCQvZiyhhbX0/W+TkfNAKUW47bqmM/psRmAJaK2XntWoLKUnKVqGYWoW9fE
NFaAOOS8vyrJfGb5RYnheS96+ZKMPtLeIN6wPInJhH+/s9DZg4ptVaT+R3djK93e
7LSNhWL4ijUWFfAhpDubpOvUBeeBHEq5OTU/qbDrucDr9z8FzPtILwbwZprNk0sR
`pragma protect end_protected
