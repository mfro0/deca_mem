// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:34:59 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Vcn2pGit0fXn5k1sDpPUesYzTF5k2j9cNQXg5ktg1neeG2Yk/Kqn752grCDKMrcj
1a6x99v20c4zq7pDi1JpCThgreeQqIbxyh1IsfX1PglbVmckstaQDjTg5A5abB2I
DTBV8tKL3+MqCJkceKCR6VTRPKMRuGjWz/xm7CCrFVQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31440)
LOZWiYzM2YBkATlSv9LnVYgItgGu4E6MoObVCUN8b6n7ri1cR+tzXwg6hOb+HLRh
HM9Ry65w0LPsCuQPyqpaFLHsLfFnwFyyHXn+s5Bpr3n8F63RTZFpztEpqXKH3m1U
jsSwfvuDhoLSJRIYrSy5zEvjHE7eln7De4cd+eHm9rsbWxzP5rjDsFt8ZZZ2M2cf
YwOV93+XEYu5t5DGW2GkPQO43r7oOzF0bMAfJgRdT6TQRJ39uGcgJ8gIDwPpkAAo
hgCiPy751Az1fAKRqle5HgR67gq0WKcFzd47vxKS2ML9j89rYx3xVYy8wFpkf1XJ
PfI4AcQ/Xuy7cagDQe3Z1tFTmn1ol7jX6w6M63SfkXnVjJLI2fU2kR9pZYW+B4or
p7hpqpclUivCnntuoyvGdV2xjKR9ZLNc8jlkKId8NsF8wJxwRYPs7GNs5VMJiUII
+3ZIGAHT0NBls1FYQ7mEbAGcTxhdnpYRkwU1yvwWrP3qc5azUu3Z2TCo5K9GGZdW
lpaj3A8ga+VV9o/fisI0ini52dkSSuHTwkgbnM2YHzAPg4mpdZoTpOKslsmksnbH
HCfhNnxZYaWOzUzf58cK/h+QV85opY9V45+FdlWvsj77lXbA5ji/DC0of5JmYP+K
0GUzNR/Heb47cO9uvchf0aeSTsE+7hNii8uoeAZsQcNkQKyF1wz14sqQxv2ndyco
feRfax8b1lDXIxg/aiLNlQ7RSmgJAZgG8gDGGdOaX1BrmqBxIHDId+kHVVm2XHZh
BPNHjoOe+jFqtmDBI+oKsi2yj3iqFIFF4MuTDA48GZ5L5c5QljiRZe29GLQdIpZY
1VTtdCVoU/WL0M/pMpnI5bWRwVNlhe8XGUxK36Gd6qGkTmCuc1w/W5SJcGv+zj5j
zlD9mKuSM7ga2lHTT5krJAnCAkClkyE87FBXnpRYgXpztjGTLXX1Q2koUpIPIVnx
pvIZDJ2i4Pxhg2dIGuzqintSaxvDm3P8IZSRBrRN8LJRI7gdTwnNbmtJIulEnVpR
XLGAXbv66FmTE2dBfJMvYewISEipwaykbJ3DPS32Yp1a1CueDlVQdVx6Ziubd4RJ
TjTKOGc4JSF0p5CueloFfEAOCaK6SiDfVM0gkGJeDeFLnpMY1QQCioXe0DdN91on
FuctcBpR5aWUacf4fTNA8F2i2h7vZbROcLjSVNs673srJsjMJc+b8EUqXfAGT3q1
5lR/hLbv7aDPXo5f4QK+ssx6w8izGuxTD4X/NYenwkhbuOKFGh3WcDF8SGdNFVZv
c/Xa81JE+hRFG3l6cEFKgEy/9bp2OwqPl6Bq4bDVwNHGt/2zBvI5l5mz24NN6hkA
0PL4wNz1j+ufzrG+2FQ2/fGiVJ69bOOqEp+YvExYkKh1psbT9kvF4u+6N0FD6otP
RMQ1UhfFy/KnU1ly6ZbQQeslGqwBWbLljrX5y8QGNlCIdMe4wy6N7MNQwVs6xN7c
44QalBvKkj3Kzyx27tkFdkRhmvrnszRJ0VK3vfD9WEpu0bNUJaJJM4L0NqHGe6aR
4z5vLMO6oK8XGkO0+D6nM4Chvy6I1LZM4zn0kt1w04/t9RXnx0zU9rfhefiblbTx
BXHFuzpmGGOVhktvP2TFZMamGs4vE3gn1E/fxNncMUYFNUb7ViF7qmE0PGEIPYmq
/TbCbpo3w5Pe/+FRzWHTc74I/nEt4VCvE+aDEPtEqA0PhmPuTE5w7In/pP0+l22h
/igkGWGvXrBw0ayb272bsOlZHnGT+0EVchlVaOhI2MNlXNCL/99hNbzLK+K80KsT
9E9EFjXb3kjZwZF0pWZ3WRk2bK6hifki6XyvyCfKoy0KI6rleWKgyJUvB0TKk77S
xGfGQKsYa6+y4EMCv2/rpx9AJT1tRISObv1LDuU0tV3TsYKoRthnD9vy4dEfknZh
CwKAfxiP2qboIrgVyyQZUT+RTGZtjFSRYDNfCBFNm6Hd/AFVhhZboRiHdG/uckVy
I835MXSioI8RsuKEIrUKehffpDDPLoRjgVKi3AjifvsFFlTa6oCYomssZC6cKwHU
evRX3iRXfEsOs+7uYeJiVMQR7gLIaXKwnjFnLn8SyhnyePMxCeK1+sZZoeAxYggA
lHdmyhWwHk5KE28Cij5qBPmirL9ED62aN6pf7j82ilVGSh7R91msg4kzH5ILMGgI
F3a9jq4NPlVXMIS76PcREuxk2eoYgRKKWZz3NSklbHtgQC8Z9gaRmyMAZpNiivnE
BXwiYajLYZIdxapWPCk4voCJYkrxJx0crZ0D0InBBLKLW4BGQDL4YmFdf1WgSwVO
ELQYjjLtxZBG1ZOokpZiu5MQHboz32ArBOlLhwP7Y7QxJeSxg15x+FWN5EtmJsfT
btfWRY9FcExf8TR/BIPs24NBqlTPpH4UdSB/JCbkftwDdINCO+fSHL4bb4MJoMEn
2wTQAg9273oThoiCm3U4O80eR/EA7XBBGO/ZSotcwO8cqQW6bXB4gFUOZYe4EE00
Atn5ARBFZKBUuekAnzEWu1JcbuCeETjEB/tl2c1Y/kaM34bwNZ8HBmv1I4dl1yQ1
lLWkxISIfYYdCOrhIHbhhTublhuSLeO0RKeVuCkakfpw//1XBYouhSjfEI1BH74B
w0hIGToLbfYrR9xb6Z0BhXdrNk+/HRrVlvTYj8yoffSbpoR/15pnEh6G1jyvcB2F
wLT6RzjEik/aHdKBzTLmxKYNMUGtBce0mo1vtFvIIqA3wGsjxAPhZXKlnqmOdmg4
YiWixjiPc7esXPEBZdqCuEggZrvjxcqOVY0U4HoFEvEoErTmRNmowIGr/ZSmy9K+
hCpeImOvKVKmPuG3778BK/xyJ/CMXDJKrrcLqLIbJF7gkAJL4/sBxTctfyxGd0gv
ioDeJgldrmSfOe7b1vrtEB7i7vHjBbCePtGSxjZTADq7AMKmN1X1jIU/mH4aKUC+
1wAgcIDE3rJCwfzvyS+ROpJ19GkRJW5X8oiHvNCSteUigBPdElW2PNll6M+ZI6Q2
eB20RNKQqvIIVzythuYyWvE5OG4LiBDwjCTf/gUUANYWgpXyc1VNuT8DV/nsN6Ch
/mIj+FRQRUgJj0Gz0OA4Gfx/VE+g1lFqMWQ75ECukoIb3lnas8+kJGECB1K6fgla
yVDD4rkqKnFzbEI6zq+ITS1NGBYZs0UvwKIs1baz5cUPP0wpnxXXRjcPwZVspxeG
+nwvIoV89wxCzHTKXfpCd1AdQYZq/Abch9fckBJoQPGMLVj9pfKZyacMd5dzM31b
HOe15zVEvcYDdbG+THb2J5Sm6OJj6tpMozBv+c62kXTI3CShA3SiZQDzC3y5zPp6
yAADTZ8LRV4BkHuY5JtQYIXjKD5RYi01qtuOCyp7UDt2Y1tviytgGojuiL/eOV4H
OVjMNynofRn/AMg1dGtU9N3h9WZaYv3ePkzp/kPAK0lhze780DvsTS791q1MJwcr
/lqCQgw2s20JAVPoxEbebs7dwUyrjSNj7bTBukq5Nc8Y4Z1srgFhTyzVXz+k93TF
oO4c91TKz4gPxROxmSx6QLxaKg0CMqfBxeHwpTB/OxR5dVSQgOc0tdgnl/dQs415
TlNz6Yg134FO/7U58vW4uOm7ZHyEaRjw/CXPGA4n60btymiL6InRwNLvcKGdrNqS
G/k0z84GDsuNlFpNWq/KfTz73m55InNkrHyoulzPLSRrLUHyljz2xX4GXMVvPIBk
xoY9hNuHIiJfPb2XEhFjnmIoG0hg+D5M+wZ8AxxGjIJpSf4P5zV3CsxLXzOCFo6J
O2wsoEN+JAIabi3p2XvlWsMmyqWRcgYxrIC/JmrmnobumVhV5pIQ7rHP/wCN2/CJ
boHIcTsc2/Oise9hdOSrhI9K14ubatBZTR+SejbjBDuUH0771yFtq1czE+k7KNe3
FUlFs8xe0VUHdQ8QyG/YjmBAuFKDGp6N4pXSr3p2jdwQJ7NOySlF1mkyVOmrWCE5
Fw7M+CEGbNE4i+KaIz9eLYRxJvdgjCiFcE+5oJZtVGL1uxcZFEBEBLbMVRx95d/H
6Qy8XeIO4ZoVtCaT2Iy/6P67trPrzfJNjUBenQzG2zVg6KemWOWI2do5lWZZbBcb
QwhhzP0pDx/efcm4mxH5K7MMRVDsV+RaWMg1hQ2RFOA3JDHNeeBXL9F+1bVHjhxo
LJW9P6S/RE8vrdptICvDOiUcFf4HV1zH/MEtLdvurICnQNDiuuHjPb4ZVSCXzstk
9fYrByZf7MpRVEYnLiDAGe/LZsh7Q1cIn9U5uChExJQjo0rmSWWxPTReXbRDJpH6
6GGljecRHw36PVlK7fYi/Ei+hM+un7iJQYtU3zrT1IHRxtL2cCsEhIv8FstxbJu9
1uM8WKlu7P6tMtvt9sbm6NSFx0xsP1ONXMtuWCWPssnWkmy7IN1ZepX9JYlHyzmN
AUyswjE5G4zGgF196J8pfKcH3TiMKK8YKyyY0TU/+VU3QASchh9zk5PWdy0MBo91
MeNMdmCTPHD3QqAZzFVj2gSkdlZd6b+2esPoOe9Err6YBhFHCGDNq8A9idczLkBq
UwPE5/y2/R5pPI95scKL0wCXEji4HDkqOeEBAUDpq+FTG7aB9QtdtK84pQkgUNCQ
bz1wa93aUUB1t9UOERTkWuwRTH2mOan9E2RpZAAZmPW7IQsVXvRxwE2Y99rx9Tne
8o6+2RdDMsB5ToeyVYj2CnNULGEGKVcVmcDuZZACQzYGRfa//xy9FKRVeGnfoX66
+4A5nHs8tVMoXu2jmpVX3yfNJ/bPj/dzew6Jb3n1GoRFmt93rvLxS2fRv5dQslso
w3sLM09ETt47xlSvIS1F96A++m16ZGSAjJDe+Yo2O869WVXVSozAB/afs29lWVuL
aIPVjjXXqXFxcuFCHOort73AXj361u0jMW86vJ2TBGjXROmWCrm9c4Y2dfNcgG4M
ylOHVLnXoomEyaub1sRN8SW8eCCIAcPxMuLlnE4qtZhPWP9n8ShTKpIvwC23fQ0U
vxoaJfCWoK6QPvB9pSjblX0E+aYIVhA09vR7qCcyi44A8SP5RySG85E6WCsxeKat
N9552dtm+rsh9JGnVhsdBCPDJvuxEA39of+8DxgrEHYg6DHyQHc3Jff33vR+hJ71
oMW1T9WvgHcPr9F6lv/i4hFxEFhPPxnLPDtg/E+ujxqlPufhvzVzCtk1nrZU4W8a
haQF/FoS8BaHitE34Kz6yj3NH/4IbaajekDMXG/iLz129NGtIbWrTcTLEia1/HNZ
sspc62YOkoEa6IS7GxoeBemgdFaQvh2Tk9VHatAaIAEflN+Mntl27o9zHB1a8sku
vysJTvKqkamlTVO1/hclRJ5RrWt6gpGf86vdfj8O2iANPBjapYqzqEAMa9NIzmhJ
MN1ehrQ3qyoP0ko9K9oADNfg0doDgZgq2g4yZTd6ErYr2b+IkN69JyKNmZu5yvQL
87PTHcSrJOa/7EUF4vz22esjjPbqrPSrv+SXYTUBsKzzBnTVF+q+qpkueYA6iXsv
HB2tg7d0vdM9Fgy+C5L5iqhSh/fXxxX4tVTVSkZwwTPzqUVEzQh99yAVkBzOlWB3
1WduLj+ixo2QzVZcXFJOAwsukHvZgk0kZGGT448ZfyoEA3kZyOkLE7hPP/6WgKiC
AuNzdx2gYVgY3EVt0uVlLIWYvkj4Am3v9qAU+QA29cgvs3yCh1SRC3FTUh6/Ctj9
384X7054K0TSCcILApKTaLkomvGOkRdhNYZrw1etWZgMq03gp2xPMpFFmovE8dBw
I6PsDAHOjezI74Z24I7z03zLt8TRVLFzDmNRiPSXjGug5zumRVouOsq/VtRkgDuZ
6bbv9/C8YRrBaSWU2hBJh1mczOF6G2KLqGANXQEEOKYExKyvDpSTVBMtS1eyyggd
toe50+6tJ0lZoFG3pWsin6S/03vCt0U2o+WuLGkzBDVuZldJwQ3yt+Dnvjw1vi45
lcNNs8+8hiH4IDkSXdfBV0Z5URVGkHj+Kg3SUGoXdqOtsv1R3OrykKpLXXL2cGzg
BFzy5DsiRI0cAmEKOdkjoV5p3oIgil467gQaJRJHhwp2gn7dYwj8+jlO+lnMHx9j
HdQVX2tZtkb2FkXlc8yD4hIdL8KibTffwAq5lJtBZvtCsgOMTyp8MCuMA3Q4p2og
b2J6NJ1y3vffyR3ytQes8Zawph10zswrxsabZFXYtoUTndptUJL7BotlwEOZfZw+
u4WFB8vjYKClITR8GzlRLwjuJfwjdrRdPrcfUEwWriCh8P2JXPTK2xYNgQgrtJcL
Zm91/lpRfn+be2yCfgAHZMQ9qGvI39ORfPBj58RFgl/+jSfnYxi2TaV4CdrkQAqw
3wmqWIKD3CP2AAUMU16pnP8hUriGvxDrprU7vX/Q3wMAOwEtq/NQ/30VxHV/Wws0
ndK7lWv8O5knP+Kud4VOckPWjGg3CqanFUi0mEWvEwM3PuS45+GLKCqwDbaYdtC9
efj/kJ9C6AkEvSo4YV/m9BcRymwKyeLCT3c0CLn2rObD7KUydQ2qfnNph8Lp13cl
T4DqggNCLvtrqFqVbZRHuhZH7muYHaFloAJGc/UJNiKDweMIeswe4lM3AYZQGVws
iTgKKNWT+K+S++VUDh3uoHKGtTAEEEBGh4koVfkaOGbilrvD5SNDToFsDKHyuni2
16hRgzr6ZizI6+EF4NxuPdPhzuseCcFy2bnUzAILcYaEdXqbsHi0YLEl5cjy8D6F
FvaDpMUli6htK63HrGvS5YJLFRZKg7LxtU+DpLqpKE/Jc7KuEMpOfeNzUOLSfjth
1lGntCvC/vspw72DUYH1TYYHzX/o54Z3x4t3HoUiOGWqNKYuEIOaQ5zwT06KREfM
ZY7j7R5fKCO1PBCHPCqzOKxfXUjKgLSAQtmWp/4DMVJ+nvFrXqWO30WzbTujI6vX
EDW/GkCydv55VYggDrz3X8kW/eBop51WLwfRdFZ72tvWfNgiVOzx1CZ7JRKBu081
mpYSX1DZZt6iwb+UyW/csNQMXQi5S9/yTxg6WlLaYvsWBLbWrauh3nIobKJSPQXP
HlUp48B49v4AZRJXXBNcCjiU6xWweERX+elUm4/93hZc//UdzZnHOUDn6vaVJptM
bRgX/EyUe12BISPjvUFKIJR/J8Pu26bRL5Web3yfN4sVAv3Fvstgt2ep0eilQuNg
C03gYP5M+E5WktELDtzYoTi7IYXKeGsr3ODQ78HNa1UlTYvUEfnGlX4IjcdY5bbo
U8608CZPlbdE9CmYS+xU7wQlqlPrIn+wbakC66lzEbnthwpPdPqc/0QUnk9HzH2p
ufERmdrcnxQfHLYrMZhhsfJTlDb4SOsMrWcDouCDlvOw4YBpSgFCP+57llOo80kr
u+JgXWV+FxEFopAHEtNpCQaHLlpCB5l1/mtEm8xpPsPUL56n6xm0Mxbs1jMmba1k
3Qy5f4px4d+V9yCPlClSBfmeUxJQfOzO6OaIBZDuDxWWJ+XDZw9MHvf8fPC3isMS
podzSvpD6q9gPUr/yfL/n0AcxH/OmS0ejGtC7+TOo29nREnEc+rvsEyMymEsPkKE
a9eC2rWUmHc86/ml7rItRGVESkYWHYJ+fnDBicun5cWJITf9eaP8jLDqLKayZWpH
gHLeOLXksbds8oGWY28zJl29uqJvL+UAkTFUJTqSdCfCaYoKOZAS0tCH1/PJktRl
kGkCLlUcQUgC03GuOmwHDSs/rpQ8Ae4QUdu2feX6CfeQLdVSgpMBGADmlEdnVAFk
2wyQvJ4sX5AumsuYHKV4SqdPcmaEiKWA8ZVa4Hy5F5VTvSbYp5Et4TZOL+bFK1qh
fKl+ruCwFHe/asCRyWFWgEKnY4yUjKC+ZoVppViyRaEazPV70ZQWC1aZxo8fY9AP
I4seoYSbGt2EAW0gAnpQsyjUSMF9C4n0TGYUxVWIWhMIrqptWAYkdLkjdv2xK2QT
g+wqrEthgAWsb1+1K6KgVL8hS0vwIAtvx8XmqXE11tNP9ydfXAuO/fMwaRX7UEDs
xqxhsDl4e/3iejqJLNc9SqaXnD4TXfJVcXYDKtcwRIOMOh+3VJHfR3pRfEKSQ4vr
fM35V6yvuxAF1nR7B3uCiszxZYqJOIBzw/Vw9n1pWBnehCYaHTgaN8GyfqvtmKog
kbmZ7CZWlkUKOfZ+yrbX81MqtTVEgpoCu3b8Oqf//cVdPPeC4KbN1u1JzF8HhOHs
5oiZ8H188arvjyh9ngY/Uj5Ldx6wMZP9bQCJSps8wwwdplOqEfir6aVtzkVcnKYz
jFFb1wEUVE7KxmMohbIXjguh03oXi/9SlO4WLxOBmogn7xbvJ/r+Xog4oqzVL2V4
+xplwjbetTSU7J6FflKy7HJeTRnH/IoAAe3ysvyv5R22/WoF6YNoKsknM9iHplg3
wUkksHx5+pP/NDINJJcCUcHBOGv66XOZKXytj0XccdAsd8/SLTmsVooXXM55eygV
gtvULaPQlk0TquS4Z8gDIsvBLbRd8YX/L+NlPtjO33ZWMiIm7+fYQJsgzGHvKSac
WddYbCvCIWrn4EPV2A0uUAeWHAXeJgLNPi3GR56D8JSVQn3BjyDvsvMqv2Y3QJti
SjFThuX14f9jYdvalhtSp4xmqAh+Y1H/m4XD2StYn8Yvgg95Pxg2BmOIuQbPS/lN
PYx/srvUo1BrWXjLrWiJYLztu0TvA5zzGpdxH7GdIu4GZsN15kHwH/1a4NISDptj
XNnfjTRVHyGrZJAgWlBNQjvFvH4NLgBW1dVlIHm3q9hzk5ogy6/kP/a9K4Z84/DG
kp0V32bxM8R21y+wTC+FMd6J1sHSRgS5AzWgLZy/DFiOUOyXkccovw5iV8MS3owO
Z0hLixI4evwxBrXhU2/asbgTIzpzvR3wK4/pcPUpNeigI+B81vDAQiSqQK/9cFm4
F7DTfT9R9HIV4Ukjc4B9VnSqucX6lZ/GZVbGPd0Bm7qzDC5Wpx02IAatVCFrjs0f
XS6ZGi1sfoZMbANeaGbTToK3/vMw7muUXlCKI0GmIFDEO/z2l5gZ+xGyq/yhtYpe
a0ebpYOUoyJZ1Day8pHAT31SAu/x2j0k71rBzrhVAzdtk8m+Z0O8KKUijGhfXRUj
JIt6bKtRXINYrZH4fm2d9liTTCPUvvb1//49ln3sIgHUWGFp20Whu8Y8nemfOl2x
q99YC5ZhK5kCu0Z32EQJnUU4sT6X+6iaCNeCAigxHhHY4DO3wZ/nsG39tuxXcyOY
FRyTnO/jwhJAljZsWDKgAmEzhRndpl9zL5Duk46VOV4SRSLQerHnM/7tf5hcXa44
j8X38InoXeKhvr8s7AeLi+pApid1XeN2ueJ2lZWJ2lPH3Ong12+SgbkXxFeY5bzc
mEwBaqvZu2zRAlEO/KHchzNbokKG2xoD1H1m5xtndX7VRCyw5mELGeyycUDNrInW
6HH1ilzMYUKNyYgBJqWv4VYYVCn48znqhPlwprXbf0HeIZtn5MaOhdrDZ3nWvxcG
YIYFmQ5IgjE4XXMO8mf8MujCnC6OjKQDeKhmRQWY2uXSeNP4LnWqIJg8QjfN/BYY
g2nsjHL5HeRVMhRuuUL5GjUExDdwwEAVaAwha24qyPlmHWV2O4IRMxKbMJb9q/jS
+JzXivH0PjvrNlyA1kwaE5uYiTRCHULnpg3I/BeKMByGsv8eIQnDYl8fXHNuKDwx
OMTxDELSHpAMzdEUKYHenVKPFA833ibR54E+jCi97hkikPjGQvJMz1ivEuHxiO5B
XG6TZAvnqrZftH+C5CXE3NO9DpXQk8Ij+jQdHiYtjbjpHIelrrUqs1tbmBBFz5oW
aGsAgQdpOJ3F9Uh3LGM5rgTHeSA2Lxo33CIw/K+Vj4l/1PJDvvTOmnv40TZQqE7o
sJvS0buTtwXLGHRPQo4Lxe0u0jza9yCE717CUMH4n/l4IlGmlj6kAjSSjT230rCu
QbrzgxrLl7pStSxW5s3itl1yVePGTJrk+zuWbZnn47kpxb0L9DsD9fP0oFj9A9d6
y70sLiaXubjQN3nZHu6bzDhnHdj5gwThJgEvxpBiPkj0wy+UyrfB/Rs95c1GJKic
hEOVMBPxaZCOzqYYmJkBBNv2ngAD4A3yr2OqLDbTXlKcVf0IMgQz7LAN10hpDcwB
ho6aUhM5BfcAp/fK6TQu2OI3O48LoY3NfpiWbLxZMYIwVAB97CMfyk29HuCvVfph
rbmDNzYBi9aOYu0S6Y+439U0ixIjr9nMQN1w5uSdj7qGwCvlSL5uYzstIkNOwWaK
Vk3PNEl4gmTDC6wQKzlNB8gI7aEkEUeaZ3MBTbwLei/TnWaW4PY5LvIe1zRSBrnH
91DrpkzAecDOcLGNGIp3M432OvsfVoj7YzyOZ80rEOwZl2+G7NrKflASgHzVOPqt
n+WC4VEjXC3DxzJHP+F9CyOStjMjy464pMyZeeOH55jRqQSJX+SEgY1NysvTXx+n
vNX8oQl6c4fQWR8uRaFUpuGHsc2e4zFEUlp+s3gsTI3J5PuqU/bJ7oCI0OZF8BcP
S1oP/SrfS3Nk1rFL9/RvdZK3ccH95iVip2CXtAKG8wGFNwOwPHYSppM13p9Sfvn9
ZTU7/T9l9wYelCKzTvxB7KyOoEkrIWY1dX/K5UfqB4Y35JxUWLrEG1Dkq+NVntGN
wygJxQA6ahfJU+gblrOOTTboiObHguuo4kAog1iaanuL+z+A9+NYTkQysLTjOV0Q
IOPrY7G4jqWcGTuIgn2dwSTjB1EKj/ofwFblFOpHbR2tmTGxVEgxksgkK0gx8UlP
LotoS6Xp+23VEKj9R5Lla9ZoW5MotZUmsGKnBd0++LE1XlXTMum3izSYdYi5cgvE
mCFdnffEGF0jjVe7ki5LSIVmVGKvJC3Dr8wIcVW1lOp3wDTVibPgECId4oq8M/jJ
dKyp69wuXdpqTcAj7MvOnMTcPZB75apK2slSd/YdTEKZFPEgksbUIwwBvZjcf3SQ
Yw4ckxD6n1Mo1uMtgWbyhcZET1BCxfSyUmJx6mW2M38v5lL2/sPeqmJXW1WcxSLv
CSLD1Ab1rQBxDOcJais4Jdygq2Cbrw9VN5+PI7nlODCIzilBZ8+qjio/AGgqHi30
yrnWi+/q48qYN2aMCpgY1EEns2MDCUyt5Fd9WFrDRLWM6es6dskxxgBvGnBY2wkh
QlvqJjiCrkHEBraRkDsw+Z7+rU+Fck3rOMbgPbt8tRdPmbWlW7j+0jZAmt9esaBg
MDuhxlIjBYXK7C5AZKR1BxDWP0G13wTNpRA6TurpQGyuKxR1q8R1ueG/S0aOt4pX
BKYOYSZ+C1/P91xY8wtrHkYs+zhy6iTrzR8RulSPlMmhBy9CZrYqkyCSSDnHNvtV
djSjfAlRqE3naYidlwx1M7d6VsZIU1osVd+CF2T4SfqmSXcb4ELgPY7F/Bw3K8m2
ksAlD0PCQ+6TxLV1Smb1Gd8lB1QKMA9NQ1KOaaNNbwUKzfDeystDeR52QtUkHthp
qK2gPsNaTEB+vS3D27Qwwn7d+lJk2nGRPrw/o31/GQaSgSXxpXFIT2i5auvBAZVo
eqKCgqP4RBNNPrRQFV0aAYWKj4E4Eg5HRq7ZexjsS/gv+pNE+RETe+BneirZPYWR
TJmLFqnJ4WBRk8hVXvFOq0J6bVRQ+AFrTt4rTIxbqJVke/+HRErKdwl6b8jdgudo
0QYxWT9TxoxbXXu9K3BCBwbKWRewu8qLJ+cJMLX+qqJXuFMrupKAM9oG4hzwvvoQ
D8Db1NdikWzY6MBwACODhSfq7eEwwLIkd2IGHfBF5Bjfxq4iu4jgRVnfxEo/B9IP
X6KTd/NkrsFba7ewgc9EslU11YnJma7JErVnASBarAdpnEx/LTBaB/I0MlC30HqW
o2GJokfHOsUPKeT3h5c+66WT6fT5krs89Zp2nlo8k/HjNTRzOR53CfpysbMl17lY
LEzu43kVpLfI1Za+bpdJDB2xrxd4SsPyqy6b5re5YwizU5bmLeR5wA8XYKm3k2Nu
RSe+oc+GIRiJJqANdMXcFTSHviz/3g5AH4+yntaVvphO3C+wryKmaFOGEnMWgnjQ
FhKkhDvocR9ka/0310LqTb4zE0kBd7VL+bCDP6/7/bJTRBRMNZU8FVjYhtH/L/Yg
24S6/Gk3K0Vlu+XpVrkXpCw+Gj0XtQfTyLBqkeQJA9ssAV69lDXjzVUKSEH4ByNE
fD75WikaIieLNcvaWAMV7f0kFFtRRJOEkftdtDV4M89H3fRxozP//iSrPc9Z2BF2
v2wmEK/Ogs8MlZXHK7yx+1fNVAAYEkxBw1+uV7ZSqlOMGfh9WpjklgcnvFxwRJe+
Uo2nPgITmDergJ9qYCSI7H03xglyifCC3wVo/PEz0j9Q84kPIQdKKSF4c+/ugbJF
9Fux7ypbkwXYhKM9DuF3iX+p3cHDIu9JoLVzjfY9FmAUkzocC5pka1xQiMs4ztFc
VfdnAABcgWwHCl+iJYxgTa9LHVzZQ6Q4b1ZGYMqcYrK55T59xOCd8Os7zkcnkt0I
fJyKi1ajKerHnjN6L9YzS7wPZUeGpBHqm4oHskUhbDM0HBnxjlqfyA3WfNGWx6Z/
YiST/risfWrPw8Y/H8Y5XmdxET/MCGYnPt834Y8toWjAvdpobNix65vwE3ObgUn/
VjjIGmYKJHAy1hCIyQcjmeT0abm5z36aU2pPcxtbIk3pMtcKac5Gabxh9oK+4A7e
MjAanXtDgtpBSWyUqx3hwH+WIlWpGUNYxUYpJ1X3NQndqX7aVpszbTE4Edh8z8bV
fy5xYEBsU01CzqerZPB0RHBJ/dYysod6HmIF41QSPYXN9hHFmLjsXXNG62pzqmq3
OIDG8cuoopAQR27J2tD9ccHL/yR+z0mQ5tvTmQ0B43iFzHCTobGhs4bD67PEK+kN
ymr09g+D/14dkT7jyOVPQlf103ximR2OSDEWISmIUvOthYc9GflD7J7WG5OwM8Bd
qrylSr1h1X70qhBqr894yvV4xINJ4n2aiRdSoKOPtR5TM+BZ4my1njvHt7vAzOrm
wcCU4O0Rvh3LXh5dzitJdSOP30VqkWfdUKANo4fbcpgdEV8OdVNApwvpVNX1jSuW
gMVGIeuA3j4t3ULaMOQSnx9CtNGA0K50Jpwb+rIiT6fmsHOUR/APBXctQ3/eCyxo
66P2lctSDyfBglpVbgNMrq95irF/iPlE4GbM9AL4vNCQ/a34uT+0yChYGgyoyEBj
Ah22wzKtB9H3qoCSkVbNvL832W1Dl7SFmbDPJlNnQyUkhzjQKlh14+yi8NXZbG/7
PQYuXMj+4x8Su03NKroXcfQ0Zx+ujevryDOBfKd+tFks1RhefKRWHqYuqyZ3PI93
uOSP5F4vFEoJd0d5i4t3ASRkagzMWAQlvrPC+rAc4L1zZzm+tuJZgw6c6tuPkMa2
YaQqXFZQJUAjzz/9eyt/fiAC/Lc0Uh/DTh5rmU1aFrZDLJ6ZzQB4VUGz9tkPZ43j
wltFjnMW8Y9n+tg2Ak0FUQF5Cd/45eezKEPyucR5IF8VvIC9Lo/fsfOBX093Bu4/
dhoxWceuwk8bV/9HmpIFHJbuhNtZ46I3Zn4KnZfqEljjFn9P785ktryU63+JAOcW
Ilv8brKjE0DX94kKLL9mv6odUwbd6NO4Zu+HJDRD8/hQ0nrRIUensU95LgR0Gu9k
OM6DZ/QbSAfYeiDmhJyHb0mT8YyMjQ4c5G9tm/vIiqXFM/+T5rkklTCy/4gNWXvu
YU7klvLlp5at90FFPTp67WwFrd/cx9lJofw85LOgF+EciDOcpFd9pkd6X/9Mm//j
/BfdomQJJp4u/Ay7A+vIH4rcZwWk/VFA6niE8Yy4cbCeUcITv1FvFrOi+C8nwzA+
GNerSfCKv3cuUpixbSQ+k71JCLNiUvkp6n0UEdjBgdGWBU1tMyP62fli1DZ3CQ2q
4XVXX4O6D70pfh5WS4m2IVJUDsTFrAoY3dGNr4N19fu66Q6PQSvgq+TFO5wWLg0H
97dO5MJTYBIe+gxfifpekidOR4QPCZULMAoFF39v1aiuLm5IGaNFn4GtvT1do8xl
r3OmV6wmSCWnxnIks7+fp27sOoCDqzKyLQRjH072OWgVvVnPYNaiCs0jmGG8L3to
IserMAabqX4f1UXYddKmX9y812Hvkf13Sc8iPrrFQ7hd1CdYiRCI68MaSQRpFOsM
igLcNl55k79LWSiuvicux5zng9k/Uwkv0t6iirZM7MExk8ru4v1A6dW6w/twY5+O
Z7rR9IO9kho1J6ysD/1IB5cB6iqLJ3b/V35QmW+R4Iyjb/b5S10A9PNAEtm8ijJV
HfsFAU9hkyDfx41rhECylAKJm8cAopdDtMHKUDHtpyjKTgkuROR7QEkKXD5XTa8T
GBkJcaXv7zEJlAD63RZM7uQNKCWVs/Euk4SefijZyWxydJX8rZnSUPrBMdvV3zR0
UcQbNgWO8/8eWCPHhkXsvIMi9ELMgFbuqUT5inatmeAmnUX1pqqrW7fbjdU4KH4L
bHtS9f6h/dnyS99lP27Q0Zh32AFgl6XfL0l/zAMgiY9wofUB/e0yLw1A1Y7rKMxx
oxK9rk4o5wgEzSZWoWeKVtXATXFXPqDzLnr68ABwFEPYy97xXF2WmaiOAhMB2bZp
Kd+/8pSBcSvaQ8VsAeroAXDpLcY3O/s0YLfE/awpMm1HGOqxKqatAm+avvth7aYt
3j6I6H1JiSybgOBX0B1RYBw/3nweon8At3guhw1k8p0qEB9+xjJb7Y6vKUvCl+3g
ZsaOiefEs+eQdADG44IMvOB3TLig0y4byLvTHM8ipkeM59bQdwO4wfsqQxmgJHMD
nC6+VG36XFPmYsvu+TCGsuGPDdbULOo3FV3yBcIXccVnLDyctYlOvuwo/tGFf9Tm
hll251e+iBwe+E2DkKw781SbH9g40cM8Giv+Vp5uZKCu/mwvtHdd3BlS/9G9X2mi
8e5RXVzZtHEtgXyt8AYckqp2zlS8kjVq5ny8e/6PAJvYeilBYFGZ94OrPXigzCD1
A51mz/UiUU1Fqw9AsyaHLmLCA6wFFiII6qd4sE8YvwpPCQRwtuy7FwjFu4Boib/c
AeDqpF+m1NXlKxCX+ase7NwYROE+9n9psV70vfNThwVZ+0eyvsMHUdydVWQvkffQ
yLzdx9SzWIp2IUMj7F/IcXvOZgnpjLWNVUuC9AyFbBpfo1dFYmgEba2/jmNSlnpE
icnp+G8ia6r25bFSwGxJlNyVT3XxP2roIyTzBRdnB/OuDARJh6D8os3lXqepEESp
gXKTyHZN0uQ6YvsXY9HeNAk37Ag9KCtN7wTcjPf48KUWVM6TSHaTH7kMoeq1ApQa
PfuTJPOdPGzNHzW1+RV7tww+pjpXM/M9Fi7/96XDFT/Xt2s0mo38cwWqJZgS6Ovb
pi4VA1h/vPfTxDFdJzfkSKabGqBYnvjXctFVYxmjLHqchoXZlkdCZAGK70BNc1kF
1YSdl7MJteAwmqQgmq6Q8IG5DOqEqpLnAOXqEOwV/eJ5STm8GSmheuUak5WRj1Af
dLQvtb0jZ6mGiFFIBkWLpOVwVW//sfPVQD9oIIlRp4C0lyXbPxpbwnXMONq8z+2O
C871mgLMwXJA9XWfZavBmsC71qpMNB4KlQJ7aaiVEThEThc2IY1GocS6ztFjYJQt
oN7lgUC7BWSiNGqk3866K80TIzZhDxOVeHquVF4g9Tcb1oST7/i5LpH9eeJbFGir
h1dAl4zwncTvNVWinWxRDgl4PwG65KU1b6DxCtL7P2+bcn1vcGIi50VQqeoxTbXf
murR9jgWCqYg2aCQND3iYGls+pU/eWS7mkJZ1ffBBbcERuZ7dCx6mGMDnA8fMyLc
MPb5bvxBSyCyueXof5n8pAiQNP/M1KEfBH1x3FBfxAovQ2I/9pEQGHZleP/1SYhV
9ZAIl6qAkaUNAM/PpdHbFX98mHQx+MpOAojKfTGBYSn0BdH+sTW5iKeCkk1v/XLa
02p8x+JI2ehdk8KJzugu32qaEQofF40yFsgfrkD986igDzTU4bf+t1m6YNPoJ0Iu
tQFIuTqKXN9JQ7Dt42HAAEpI/KXtYREuI6s+XEp2Slwumhoecb7pq/TirSAUMrYe
G/J+k6R7wPNH5cOT90ImFdmYT1ivd7BQ1csdICGutjrD6qvnzwn434RyfB/W+VYV
NdK/pmBta4GO456M0EmRHXCl0qtffSqUPCVhRYuhU+83ayHu/Yh/3kKtIlP3SfDX
pGvkurYbn7091unakrwzLdGjK8skGCOicxaEH4xpBpNJMFQGEKbT28qgVbB2uLjN
DLJVGIIFGu0BU6vQovpuA7+GGIRKW+0TIeFQ+Dav69K1sfp+9KvgQSdkaqo2sDjY
5wV4H+qQkY8sYn0ONgp+k6+1nsbypM3DulXwWTkXHzfK6IXRSTDEePwavzT4SXKE
jwGc+kdUB6Bl9QgwmDEVgWWUxr4xbtuWp1iOceChEziA1Bn6o2mGNkpUK+f32T+5
SKD67TXqLJTpTw3sRWbMxoqO+lCK3TdMWlX4YqiO7vIUbls+iKBxjwz5J8dNMu+a
QT63IZQWR7sy2GS0dodCZUgagjnF4jiI7e3pcpXuMFQtJv+n/tTV1TWbRegisYJN
57C4Z0AxFkzE5HqwqwSSnF0ZSTbqKNkxSlHkXv0XEccDOGB+wcVXsOX+UY/2lSVz
hF5APa8eKDMUexlLP+WhMYmGWwnbUTx5w3OVMmqmwpbztZayUGEF+B98tkhjuEhu
qq5/A8SDl+v/nDsaBfsFmQBrvGuB/l+hrgxSA4H9Z9YwzELDXXRaNw/SJ85j1WF9
DPwOKgWk4vwKREXl1dUNl7mqb9EwaTtAdWGfqVUpFIqYVcRAuSFZtR4BYMMTHB/B
i6q8EL3DW3CVCCnkN48oWLnzAOktvKwrJdkgZPkqDvv+EkZ3lyNzQEeniwIf6k8/
nl7cg7uCwJa0Y09UF1hu5X8Dnr2z0qt1eDfkuEmw+j/+LBzr0fMAoCnzHKRmDVki
aZYHtmKvfvGKOPShSpxv56ve2nSV3O+QhEqEnlBJOqNbLSWYugs1da3ttfUxQRRn
uQKgxmljGvqaJdR/tfsNipAr0QNyB0E31Ic1yyXIXTrH9pNLO7Gx5N7gqHsPZRvM
TeXy31ZfRkBTHIdQmIyyvrDrIqQ5oSd9we+BdQy2splMR+hWdLuAI5X+tCc+N8if
hjbYBKstToJGt823WOuj2R+TojXuCCe/EscZvjBRCj3SV8JOOlz0tCV8qGv5Z646
eMvUPur6yNNIOXQvQBI/E09mqMlMM4uYoXdsJ1fLbjDe9eKp56c74tJ8L7OcxHE/
HF2UTQthvgsOZEAAeUSFCAwgI6vTOMKlxklN4rdgJb7A4ukwKU1fg/THfD0IAbea
a0VBLwKWLsh/k2ZvPyerZ8S/+C7hAxIIBhhroMr/mC+toqGB5Q/Uur5kCOgU7cyA
v7vR8HmpMplOWU563s1sz/aCc4LWommmf25VOqJsPKHGQ0V6+VGUA7W4/bdB9Jus
fA6cnxnVWuMxCOlaeriDRZEok1RfBuAg2EGaDkMx2kpV4AWP8TL6osZ44Ry1XJtS
2FaSe7Q55u4XpIHAo2PM2VRhdalSW7NN7SfAP/T00t+epcIxXvxMGMXFNGIczfen
rcY/UkQIv+bpHz0lYGIKF/2vaD9X5gwfPji1YjkiNIGtBwYRnAm7Hil8JQF/QuUd
qpPB36Ivwygb1w4/IjkA42WfALJKab3gIsJSOyEfu94MeNYjLP2+lzv6LLuKp44c
ejtABywAZPcuCr4Tn2oe7yez7y+epIS3oCg0vQU1y4YKCOdxBSccnyUxqmvGR3CB
JGG3aV4J9CD4ckyZfu0UyMldnI3lVmW1nx6+xVApXS0PklgmS1tcT2eYo10ULx4F
3hhPsYvvEDzRDF/OIVXF0B/C5ZV+/GBnlF8FOBSMEISJCJYPx4jkyk/gDNXPl9Yw
uEGl4LSF2sn/QXJiH3n53x/xdAZ7gCQE/J0IAnyWtABk8UQxSy91tFDIID03AgYf
dIZJtYO85kdc+2M1AxB8T5sWThRYhKaFn/SyvXeIl349/2cSjKguokL2caLLoD2R
1JBIa3LEQsP4WzAs/h15MvQ1cSxh0djfVBAJBmlfpzByEhZLqS84SYvUjjvQWgKR
hipPWevVKM6CRzON/kOSf/5nYVPeJUDHKeurGkLUUYfSmKVy1cNAzUlwLVGD5z64
TPeEtEi1qlB9h/FP9/EtQ7+x/XZSHo3YVHa3nn3l9Vz85n/sJ6suhJRoF1gD+Mf5
o/GBvtsIlNaKwku94XSNyJH7YbLgJSQA2kwnIJgGmZI6Ah7PcIaA6mvk9JcAynR0
Y58WxfoFScatHvUPTwseEkArwqTORSxWgYgDJQu5nbCmJ7tah3ian5ZT5kyrq8mF
DvoX46PncG7QfYyvrk/3ONr9GyR3tTYuNUBjxGeI0VHhSLl2Hq0pjvMtrawtBt5j
QAkx/6/+LduBbuB4CGMhxBTiAkRWeoQam1p8KUHQwTWqTfgG9L5KC2AUQOZ00JQE
+yoy+eEsryYY8J43fzP5gHmdkD454eyTGLGi30cZIlrfg9579ckFCNkP8eEMVcSu
WUCGtXvs/4dLvsP9IXbOfCc2TJLgC4m2XKRJ5KBYLIuD+uf3GMVfs+NgEhJS9bpH
r/lb6uYjgvULxF/weCEWdftx4Qr+owoaiXA3SY6sn+FZiiEpjdYeRhX5NHYs5HvW
zLGF9CMTYrfFdUU7s81gTufafuqsJ8uJUNpB0d/wYS4YI188LVZ78yfhwJz7Jgdh
ewjDTEaji6D/l8EWxMr3EjqObK8EJvll5NngrTP5tXg0b4VCtL3dU1A/FZJGz8pi
BiKoXCDaa9YibBET8mswOGwTta3YCnvioYjcDazE0VFnouYPHwwmr6AOt2P91YEk
9W6JduHTNjyzgkD5XQ/eQNmue700yNvhQBk4QkwQN1QPtqGXx87Fe9iBcg7ow5wu
5NcEB/uaky5JbYUbRKDfphqPSgCZu4f476YirfL6ecIMLL5eLByUoZGsYa5Hv+Yx
MkMcuP4lATIEvA+ko/dVK4tu2+BTF5eTmbgDKPRfvOhbHE77RWUeh66fZ4+/vDLQ
96Xg5BoriEiyARt2Eo13DHkN+ooD22M82KVKKIx0v9Ugobk91Va272U23x82meAr
zXuAuMvdDLSCCi5CJXW5hAlTIoc4rJvCjreyl1MrEgiFeAFgM0iDDgVX0rNKyp2U
tStCW93dBRhjH5cGaG8Xmueeo/Umx9UF+m3rBuCbq35fQMfJlUgQFVdvoCyNlGft
2akaMrlWeps+8atTOyJtjpQaCq0xkJ4j5gYQktEUzQQr4iyt2rYLwVg8dxxIEoPZ
3+TEehcg+wslR0ZuzPSEQqqURXL39TKDDbinRRKWQIooQ600WTPqy/NvElV4psem
QG2tsxPe/e51OuWzTOawyRPhvvzpe1VcUaVeK3DICEmxmgLymyP10WBtzMfZ5jF1
b3KnDLb79XktM934K3f2rT5hbikeWaOKEPL4UYHDF2XK3sHEyfVEOTnRTYdnfPi8
OMjf7moDz9P5rAzjd6thhiJTW/feC77VYcYotaeaiLcrn+px+CT+t5WGJUD6rsHV
FvDcpnJU6KfCyJ0KhB2UShbbx72ug7GNEGwCobHYXp3FFXPINa4EPv5LJD1oQ+vM
7RH5DP7qJ2emZt5P2mfg0qV51kZrbWB0n4utjvMuY+/YUAmIsHvrogZ8ChFZCeAr
s6WAONd0c+PNtyGL1Oz+V6pLpV+QuOFbbfh1LC3jxWEHcgIP16nwE62YDVTTnu+I
oaVxnLRliUMFtD23/m2QUcVhfNX77vzJOdBm6p0+DU97hrgC9qgLuqLzk1HZZb18
hDkIOyAW8tki7f3NVQsA0LhDsh48djZUF6PTVHVywUdvDhqKou34UNS87dfvviXj
kODNfpazQ6zBiOXrVgJm2v7kb1RY5HUDC98uoTuliBE+23EfvSy9eqWmQ781xP0o
mhdGFFsi7cXkrkaH4XG+AUGtW8i0w5SgtOjnnHAsrY4VXrH6gJbbBt/KmDZfPOSG
BufjSquBqMa85D1M0+J280BW2242ewpFMuRy8Vs6kYGpndiERJJYmCpZpw09gJgq
sFTjmggiMiNSJiL9UyHyFeGmG4494vebemIQY8LFB4AstKzjNdrNRjW+gashAEZm
6Q0VbhutqIgXYatnuNRK1KiZATaHntuFJdiyyr+Myeqd1j8177OG0FcfvUrDXWl2
UMU0adgbdaP9jaWsy2Kq7yofkB/DrSl+kO2hBY/cuzSLOaLazBnOfUiaWLMUERdJ
rh+ZtJoF7hk1CLKnXiKXUGhfjyJ/jqiKaEc1y48T86nDWaMj3iMfLqsgbbvbVwn0
6Q2XSo5WV392Zokiccgmy0DQm0ef/RPjsj+aIURFeo7wonN2f9t1XOJNBWCtcAVB
cyhmvHon+di7Dgsq66d/dulkWZ34tYuoTsDlBttjCXeL2Tt9PmtWZh7EPptmaI6Z
6I3tPt+bZ9lZXhYSAwkRzs3y+7+7xJ44auAWg0MwRKasOTXGo+WsRetK+4lrBLJr
ojN/NGWsHpxfhNAUFm2pkXR1lLT30cc7rgbUEamBKLY1ljiM3aXJB3l6u/OrKZNe
caDMliC5tGdX1b/29cW5eGucb5NXWFq/kTIbfYKFAg7Qa0EQ5CExoamZAjAbQURo
DJAn9o3UV1utBtb2VtfUAsu8umuk+UibCyY43p2rvkoR9u+w1ZR4remHMotqZYKe
MCRBs/lXrQgl3myEdYYFpuJBJjxY7DgYCyBbnabpFC0Rqqfv4mZWcq91gNutSDvQ
PjAKG1nda+QYzgxqNA5u7XSH0eXrw0L/O989of5Tuw/MMGjAZYbQwGvipMely9Ko
MmkfHWuOKxnOF7hcXk3o0nEaHvyNB8XNUDExG3+4f7BeO2wk3f4XHkF7wQz6RK32
kOzw9x+DVfyBiN7WugWE05IoHsfFnOIu21UlsKpG8Qhqlhdj1TlA6DyEeu2Tg01y
IowbMMAX+992W5mpyQs9pvSReyxWU3zIEm47VKbXffnbSEmin0WJaZ/wiyLLQrZw
T9vE+LQXthQf2kQlVZhkM981oph6wkKB50ApVB0agUxQ9T+EgR/1TDM57MfbvD6V
DQL5YhMb+zvwjPXCt+bCstciDObe/KeUgqNXQLiAd7nr+qH0U6amiYn9pELNmarK
w7k+svo172QhbeSaP2YfRzSjKeQcsMcQ0mYd5XKAJAUMagLa+XVJB3Hb9DsmOzWy
XeVmUAQ4wchxf+sEgBRMrQJVroezccf3wuXG+tJUrpKULklkT1A9wcU0gzZUatBW
+opm7cNtBzxdGwY8QcgYjjnLd+w0wbnCaqVPIf6/tYzA9W84Fiog8dQRcrB2GOXg
Ii8gbM1a9Ex65udUS3LW14crQcatB1n4LOc4PMjCgn2JKlLkHrsTYcgvZLav/zLt
xhL/kin8KA/TvS8w4qDcRe9NMG8KAd7oeO+emyRi/LK5p2YIIJDRDR2phGAwmXT0
kamQ3+saW4CGTRz0ViHl6i9T5ZFXWdTcC/O/IqSEtTkQ9xXjCeHITTs5QT+QJT++
KcZlH7RI60uSuywkwRPoypItYjGMdJmcejLuBAnIEcpoYyTw813laRIvuZM0YEnY
1FxNigKHFfDrzTv2WzzJackOBZmcFPw8tDK4+M8NuHcGNjp3bNDGrgLJiTKq/Z9c
QH4jP80JW6eSJ2LRWolimQ6xtauHq2VPvsKcQJ532Si6IlBXUrvb7m5uKXv5lI0a
T5WkK1sFHvdLb9LnJir7b0bumEnyYIvS69+QHLoVbfwJh/op6VC7B29/4zYgxT3g
B2gs6sN6O+5kbxu1nDQ+bqaeJZtG0QLQC0E9L+1pV8R9fvtAX3a5YVjrYahsSHYr
aTA37Ci7Pz0u604QH2UzBUomcaVSJLCdHdaG2QarBMKze+aDCxc+i1x2I/G1FdTY
piMsAsWuox+9qmpv6sZi5PUSC2JPJe2AlO1ueb7FE6TOUrahpepwp97S/4PFFDe4
ujqZBOk6eU8A8Cj7NhmTs/m5mRe+fTgnNoxZWK0ZKwSh4FEHzKyfxC/8U4T9c2aq
kfMegkWUzskjmGaqmq/xJOX2xlc/bMNdvkWR73Qwx0EK9S0wAT7HKK+hq+PJdBwc
6HwYTbWpvVkD3/mnqFsptr6J8pDahS+tTp5Lgknfrlt852y7kp6mWFkjug0sgZa0
eAbiA3TPuFa8FW52TjU9uSv7FsyLNlSfbY7ah9ejPNSQUzeuSEZpjylNEJkBhbYm
FQ0W1w5B8V2tBDHVuyasSX/lfze0f6Oezi0vS7kPICd14s5e+SPENHFlYbSmBshK
M79W9o3J+tlSf7EJNLNJOtz0Au66IHsHvIsBq+Ai2mI7m0Td51+PmZT3UsHkj+A+
oHnzmPH8jovWcLE8hLH3ZKrp+QtjRp9qA/Xvw4EMNE84O0DUZIsWh4y6sJWN3I2l
e6/NOyz+kCo1O4cMs4AdRm/HQ4O0GSZxyM+qMqWYu9N6SNL3suxFM198lv1ovRYx
uHinRHJAFztGxkG8OVxCuIKVXacMxBBFmP4QVtr0/jAjnJzOSOFLfj4yp70DJqnL
q/cEiSYuApG6v8qUWQstuK85kOYc8/J/pz0Vo0WcoXz8TAM3AJ5oDk47DYQiqtcC
/m5/dTqGVSBD46y/PkYWsXjnjn8KwoTbBRVr9qQaN8sbQy7SU3qqEeVpPB0rKcWb
X9zxskmwRKfz1OIeu4QCg91rAkhu9IFDS9oHMkTEszmp90KjyiJHW4H7Pzx0enOR
zqRNV9p6O8K04Ot2PsuvmaRkMOnZJ3GY38VvblTxqJIkXvgzdhL2rc0vibmz6O7l
iyIvOszoHgYbWCtcTvHjz4CcJ44LO03dIuLcFQTqOtn3nJjDwRO+v5STkfo9b5U8
H5kEZRV0nQsmBjpbDVFkvIxUkirbzjAgAtQEJsnlYBIcF7HDXfQjP2kInp8hJrfX
wXs11um3ArBMEym2RPLQxHYp29hSk88PQPhidaPUNDF6v9kB41VPK/SC0dNLxWPo
H3zER/8TRKDpMtQLbr8qJW1Sye257/SWbHLKTEx+Vr86XNnRBiXcbwGrcGwQir1U
QWecMs0pqGWz2U/LLxgr8dKSCjfcXXR0WwblHSxom4ue3lqrs19iDKMTpm5LUK+Y
AqTgEq+BhDZsqBkJTPSKMMoNeRCekcPWoFZVp4XeuYxsKle7yrjLmBJW1Ti8P7/e
r4PCOGshACs8RbsKd3NEQ3fPk+wrPAq617BqeF3eWH1/5B/m7GfXV7QZqGoYV7H7
HxrsNY6uA9fTXJV4onVv5eX/4k4WJMg/uRw88ZIVN6/AH02656ki0eLlKi9W5bhC
PbDocLgQmAWUj978Lapn+CIeR07t0RmnSDEfzwjtzW+MFuVUgT5R+ATgYqqVPeJG
YSdpcGDgF0mctTnY0iESrFwMEtI0ZjIdXY4Qbt4FFd2/iPIcUpYABNsPVk2kIhwg
E9sNbS2VKLz4zIgFgO39eU6U4c4Ym8VyhuhYMS4W4m6v2v54VBkf5+GSzNAjlVJO
Ql+D/wRGxB+OPCmS//ID9IvJuWP7OnAY87Lkq5XCTbXJtELYniznOEdDiGffLs6e
jcYXL98S/yHne4uSECcd/auXWrg85pltRziW6rs2KHOVp2RcOctW1P0Lsp6FHQW/
TbxV3xUEWq89cAw89wvKxj/CBMPpK71kG4xY5F/faEjmNL/X3N3XzPcu+VjPX0P2
nrTkzxnjWhF/zgkBotuijS3IZtJjbVU3ZMfLSBdLNGhpFVVZZDz8n+mcVqzBkgHN
g+aNstz/CU6J7Xa9AgOQfFlUacCdc99v11gTrQi8YftCt/YlIt25F+TS0oVPEgaS
vtWM5/Rs3dyLvUU9xDqYrrVn0DHwKrO2M1xV6zM9jTsm74tpncyb24CmtBUaB2f8
Tk8xu8BjEkh9p19AFXINDgdtrwbEQ5xi9q2yq+AU9L7nyjJrD0LDCtvawhPu1Yok
tsqrgCDtp9zwx0ZBPw+MWjADcnjda8wff6Y58pYu6qHWOwEA+w6+PUDCrCrdHs3c
hzFq20PMt7+pRMkPdQpOBRQwIMS92bq84H6a+ETG6UveEuoFeBYvlGCo8xCExE6n
X28qkCOZsqc5kb6UTK/c6y7NDogxjKYLU7jGBPtXMOodpdEOw3yeToVonxu7OcW1
Mjh8Q17vu5+1j74pAc3nzK7LFQJf7BForbcJlDYW2MS60QfesMjvkY3lCmn9K3/9
DEFflP8gk8w7CgPE5B1H9sxuVS2LDyvsqthnbfQhQWEJ3f96+XmUUk6tYmueDzVB
i72BdCwXReVF24tsOhUBF6Pzh4K8UrRr9HQYfa3W/VEAQcNHGDjKRVdSORApUgJt
ncuN+q1cpyAgJF/4BkA7AGjzsL8B5QB9cJZrzw9/5DQgvBQ57T31sWjdNhfO0pO3
Er/TPMSEnD8aG7am4z80H4AzaiiVSklr1Wjy6ceg5Jqov2mtoGVb1mpiydI+ZWy+
tScN7/UARuO8WQeYNic49mc4GWosvYLFh4CjPSlIl7bnts8jxVSEAMZb61V5xUIn
0PZ7ANu5qGYwnFpUSFL1jYvlu0Rv4W5G9ss5kvuZJl94NCIlg+3D10ACh5J4wdSK
OyYcY3N2cpVw9H/+jrSivmGWjG5YsTNx94w3FyRGNUbIQ65cZABS0gGILL9gYrr5
n8nzSURjYv9IunR5KzAD4fts5OpuIvviBvs6S+iYrlijtuD9HzCEbuci+uc7EkMI
iC1+sqxCI9WnE5swqs2/dy03XJtOGyV7auASgHNns4cgS7zCxIz6tH5F9fmSNOuI
J2biLm3Q+OWEOJGyYs3o2OvseBpY5J/F9wbiBrHedJvkRPRmEvVu+98shwaj+bnb
jqTnYyLD46ePfouJz/xO/Bsk65fMBtqp1ZzuWH09+21mSSoQXO9uXEExTk7kGd8s
kOqE1XO8TC0qn7D6QcmxyfUNYOhg26YoLhd0RfNFmPPPULt46tQ05PIK1UDlKiSI
GY3yPvdd0h0SUCqegazdGqZv9amHz2LzqVBYYqIkaQyy1uStLQFXD9GruCbRCDn0
hl4vlXVTirPHcA9nFYlsfS6zI7gWMPd/Ee7Wuue/yJ8wFoay1LCqKFDvX+bP2qNN
rWDo9sH7ecggznu6+4aR+cBRfN6Rk4P1VEOwRWsNGvHqBKWQUPT9CRS6xK79dBPZ
xzy5bncvbz/0Q/0g0GDrsu0BbQe0LVnM7hP9naFSGn4qFbD6v6wEL8vqoxifEmIl
eiR1UfDRF9N/GCGCgkn6rMlT4Z+W6dOATP0Nth1EDb0zTjyxeW0xR2+BUHaYB8de
Am9acehFejt3F0YrMxbWvfFCJ/mFDwr8pVRRVDyM92rY15nm8La1iD6s5MtcfWnt
ifYFMm+Rt/SUUl8rz6q6tN5VLPAvC8nN7EfBITw3WxpS4Xsa1s8uXdaGCAf2dsu9
QSMfiRovaCTe5V5Sgii86ulg0ifferQ/kC1UXeXSYHkFMs8PEuEF3pljJ48fa6TP
1HIGEHXX6Hft35YeAUb+TpjQzeh4alrEQnbnAzdiU3v8jdNa21VrEKc7xyE9FvMq
agelyeOy0wuWO+uPfvOyVEf2C6WNwYVSEn9AWUHZrcTXMO0AhgazQTGEByIatxjq
DVZCPlUOKqh/rw5rFY1v6yom85R6PReLePt9B6xtX5e8G/EJIXgrs3002w41kncr
JC0reHMR3/uNOJCl/TDC7Lhv3EO6VU5PfQ9YWcSP00klJMR2I9EeunKWRn8jHs+x
hLPKyWAWEG9WiUPbUVzShTwgtibeTTZdpTgzubcnKqkSetBGQrsm4EA8wTGSfjw7
0t0zgpGVKUAnRhbDpgtJtyWVIKF+D61elH7+rHMvHwDaeKyvHUXvLl0yn6fviGbZ
vOYBWQkD/THffJ9xDYJ1T7ZbC6Yi1TF7+tSAmtCjhGsPLEAhrKnx7bNyR4aQgF1M
KKw+awSWQhH52gUhozxI1Nx9IJDBOPEEMjkWulNN2seDltwTExyfBEhCVovCCddn
TXxqQGKqQjNsOc+8gxnZPzagOn2qUVJ5svMpgvZal54/hXzZFDSNT9U+Tj9NC3TM
k6ORYbScBgTyGUlIZ9IWTH+w32e2xxKUfFWFbj7jVVwS+3yvZO2nJttqFm5ZdnjR
JcEg6bkHIudRJu4emYzFl8gZobVoII7RmzVMpFG0OfaP01J5FOo1nFPEuuWhRkTp
VN33FOLWjbsRU4ceUwKlUzFZqvgaMqKeKANjdv/cDV8zTGF7jZUI1qGhqwghx55P
OtEjeIN9RRPmcmOp1/8vbGtvCpcUUwVYeu8kXdxLQdHoB+Ek7wokme6APz02/8ic
5qKy3uz5/GIo6/VJVwniEQ/AOuUgRjoR7X+4rwlBamDl6D7kj8g99SETs4JhknNf
s4lnH0MmuxFjcPU0xsT70VTxhaQcusWMWJKVKax4srF5OwZWRUfdm3dPla0VfAsG
h8TopV+OIZri9UzZ15qcnoT2TIRmmxYXbHAcgCUonMu8tLa3xeptEK6SiFkbK9BU
6igtQxEL2ruKifxZ/8SJ4aD2g3HVgb+CM5/oaZCz6G9Xi64bIcY4WDlA0Johp/lG
tOLawe7Q/iRnkJOKGYDfvD/3kKI4C/Xm5WMbTYwKDlEJ2GL02a8MBJkO4CC6D9zV
grrU+BRpAGj2vu0JcpjBabraOCX1j9PwiI0FW83OoXNu9pX3H1uvrjBKm67hbZY8
RTGGPR1VXuVhzVj9GhAGB38aclfj5nMm/gSv2+ssEC85/nvf594ghqaA4JgyZF42
FxdJgoQtuh8nRGVdMYEWfFKsKHOCmXbIHqfc9CKwVWAydk/Ld76A+WGnNHBILwlG
L1Epl4GrHDFPy0slTod3H/VMLau2N7MKS391MTE2oO8sujKKY7W50p70mjRztO5X
XzrAyhR02hBQpa6iyGAjwROVFbl9trl0tMEQhLq63Fhj3B3/NJmBfa34hMMDsOzZ
P6g6doygq0VOheCnR9NYupSNASk4XYI/caNjqOgXcr4eLXMB14w7d2FmIgPWQHWl
XL6Bcx4GmR54dkoa67MtzqApzaW8RDlR3lTrGOSUC16liFWaDEisu2GuyBxGhkxa
Zhs8uzFGM2XBqTBWXFZRHPpzA5AmuIGoP3cOW4rTlFan27oWHRRDsPjiBCItC5CE
LQUR8x/i00qXPGpsV+A8he3lJLBxUCVBgUvPWJ3u36/mMqogDQdhz8sRdsm3CgE9
EBzorLq6aIpF5VNkdK/aNCUC6y3I7ImeeJZCdBg/FWydil9C0ww0fjC10ovgbSIL
1w3LVwijamjjBgOwMci64Iov4MUPrHnW0zlai/tuyr9ZIn6jwAkl6wmX6kUATrsa
JogvJ4GT9M/HwigIao/3C86cg7F5YUoaP2PiMcwTvVlwlAT1bNNmXdkoDjkiHUID
dXn2hAHsp2ItnAn7+Lh/BZujNcu1UWpkuUH1Q9A/rnAB8wn9GFLR2876XSJDLc1x
r2+rdiOXUcz3iEqWbtpiemHA4Xtd2/3b+/ZW+rjZh2dFKl44xYkHbp72REwADtpA
kez/9FtviDopEVOA8yecRbktGO9qyfeVK2fiKHFnSsfBin9Q90KuPhSUV66WCKVv
i6Q0YfnuNSKYRxyc3dJIuSFSGZdtmVCb9qU2+VgRdY2wlG8d9hcZ5NvlnQH2iIgy
/fEXhRM2QpyUgG6PwVnniPbhiMwEn9xzEYH5zOMdNI7zy2CLGZU0CTm7EGAhkZB2
9ZXCztY/gYd+Zr5OREZINQyL0neyT+oFwFBaNFifqb9ir3LzvSo4WrhffFHWBmhx
ni27fVx9CrAaR3i4dUKWKUGF2UV7ymV3ZIVvDN/0kaI+WMOIs4WzRohJsNQU9dmj
cL5yju5YAZvOK2zydRu9IwRbgN8733NdRDoatufbHYvV+7T3XtlH8/KmsN+KF5tu
jCPXGWxGkagJYDf8qATIx+lxLe1O36UcXtynnwY/ADevotfRpstpZkaorAiZXfqP
7roO/au7fxt+8UfmIagAue8V2zXYYZfeyBXL2Ulew8dDGS6VJiBHZOO122lb6fYd
XEeCoW5afzO50WQsuOrQLxzBMlV7yu5xHQ8sQPvmHnO/QU6PnaFB9daV98LtAKLr
5WqViTwYwhpQ3vGb+mTEojN7GyR4V3k8KV+CO8wfTpHs7Lem8C8EL3HPNQSU4XTB
RZ/TEkuISoQkJCYd4SCWeSW0nrMgMRN2cUzHb+YwQ0rRTDYveMgxHCZynveRP4PX
8MmVyDTInnnNhizuE4SLXzTp5IRQoIKdcq/gEAAmGPR4U0TWGCgYN1DYQo1UX/G6
TUuNiq5aLTP7E0JNoiRkUFvC2vYX4p7aplu71pgNIxVaZIHud6nzDg9vBIRuHpCN
EkAUizDiPNMN9ZIgupR4nEAAGC9iS+FJSEve1xIIBwVkF+W0XmxDw9AvvfSGlt93
sIcdFizSi2eAakDrPmBRO2e3v4HGLhgn1G4GCIz0ZnfkpA6tzYBvSzdrKENcivCY
Xhg35ajvL6EHb+E9eveP3WNAgZ7bHZXLwItBeWjVShD+i8FYh0TeklcBBckvVjbQ
kQGXxmkmLWfngWcQ0Yp+Ja21+tyllV6yt+UTrhJy8DH2cKYah4xUz1DcfuYf+O+x
w8x2GW6T57VzUaGS/CuUdBGo00Ul76yO9wbjcwzR6i2jXU0c8j8gOM843Q6IBSGJ
jWC7+ZZ92O4uUsHuTEaIZ+TemrlcsbntrUp+7Oby86uHqKeya59Z6nMJrAjA8zpf
kvsCzjNVfgTRW8RIgeyC7s16yNqtFMU53s/EClGupXLIbSR940KxJCTaOKhmPqVc
SNu+UERVewW4aDlxUtVELqPWXau7z5M4C4ICTaJG8KUS89MdCFUgnmXYVBDNfx7G
Y6sUYqV0Iwnl8sKs6U0ITYck/PgSdlJzgKgL/ryj3K8eLLJplm4LuQ1tHpp0fwvC
BtVBXLr9I0WqYiafb6iCWl44kXWGyQloEiKjoOkCY+5qsCoWJ19+75T9Fd8k365J
7Q94/MMyT/NKXXOfAcRZSVQ9YuPbfTNnN53IDfd2tkwipIQpSb9xgD9/D+4ZvZ1i
4G79RApnFhmD//wYzxRh5GVX3O4cP1GgTD5BBXgNgxRbcig1VzZp+iGUaoBf0IAB
RXJF/0TickMTg8O5BWgdzd+QdQuKwO3gEsHJdG9VqmK0indMSBHX3PVTDBZz6kWf
RcT2F9zoBe8ty8CZjqxL1IA4r7GOECDLvpDir2H02QiGE2IdtIDxk9VNvvCu2yUA
6y+2CXk5XceH4Ur/F3F2U9bax1ExV5SexmV7nxtVO/KK6AVzTXUStiCrHEZ4r0Bs
GKj43i7qylb2rXJlPn9aXrPvh9VvjrosvfjuwqIl8G4garZ40mW4+Evce7InIxUo
7lQBu4bBgQAutMlUymX+kE5roRW8kq2SsZirHjAoO4Tt2oFez3nSQfO5PGQS8M0I
OChhkstM+tS3dIIUujNOrpdj99gysPZgA9pPFTLv29h5peyZM+0XJecCf6IzCdd2
GKa3HciLobD3nuq84C+J4QzshpFR+cgp/XUBnDeyKCuvv00qaJHLLQ7PUJBe5jlR
PgCniK5lGcXjOwIdx28wHJOVtlI/3zI7U+dDr0dBmf0GjGjA5Y1a5Senb95GVqQv
Kl0u0eGPiL+XlUCRHHViZkmC61A2klTcqHnCTI0HIF5aLQ8/MD3wAq0GvjVdlmIw
4n8TFbhaaOoIB9al/ZXeSTvOV2TgNPceuv3MvakgY77RWDP/D8phroiF5UQ2NHiU
CSmTqxV7Oot4QkfDXdXv7k+xFawffRvj+QYEZGlFDvqbACdUBbCwWMiNRKcKOqly
QAx1Yq4OF39bcqRXhdu528Sq7U9a9+DrubwqVhQEcueL3Hyo2CJNm6pY3NTYblku
k24NZAj/WFAlMv2L7kQHrnx2kPdziWtv0GPXUUv9aGWPqIKwz5swFLCF8pNjgcUi
Fl2AFNSl+uOq9wII350NAbyuHt+kCQYyYa/6DrykM7IIxmW0CRRkjDhtH/A2ap/z
7whDleyy+btHQJxoLxT5GlwGQE8wtu92qSWGVm+6vMm/Lg4bbo6OqHEEjhyS8HZC
+MgBW+z7NM23apqPZciHL+mOGIr/y6h/h5X+c013Rwyet3RgtmPb3IbDlCjtrxz8
Nn+9rKYPuyt/Z7uH9dL5y4aOYAonN9uWaCGXT2gRw4tg3PKhTHgsKUaKbax31fcO
KGNOn1y5js0l6VLC+b0Uw8b4w6aGvmDKRNMlNMqreve3w+YhEfGyfhtp5xoMOvLU
+i8u2jU/axic4w5t2MRP88u4SEY67BWIV/4PQF7kOxk3DXmoPmO8On8RwxaceK3S
Q2g8AIcAc71D22MdKmTm9cGnjamMHO91n513pZXCGWlS/ntyVm/XuZfPfnT9nKYy
AP1g45Js/OtxVoD/f9QRLi+KUjOFxeG6DxmTLrlec7WmM7ShWDJ6qS/rgYmlpzlt
eRbMO88215ySLzmFq+3jLwnhG2PE6fdFpd4cVSYvooVvq0lNOw6lrpxvnyYxNDvi
1WIzM6UUe6aEM3rbBL6Mtpre9YbO+h5LH1nBbCpgclUBLkqUFsxRfkGVEF8qWyN4
ll1xAudtEyDChZQBwmC1LvhtqsQf4pIN2mW9MsHkSjAtQ13qxPh0brvHmk1/npOD
cF/pm5ve9DoOxd9Z1G0pxVFxFg+7AwKIVc4QAA0j/hezymHPJCS0HaHLQ6i92/zt
b6PPwPmL+VXVSgBLu4kChGxK4aF//VMEpcnvJlOM+qJfkBl40opU5QWsaXYvmfPA
JW1x48iSHAvInAkh89g/C+VAw5hEdMvxrQAJ39oBCHGNhlzVhtI1AiSf9fm+Ja1e
g5yDzjpETepJf6V5g3a7kwrJJ0WL/oym0oqUH1Pf9XKMV4d9L7mfoUikmpmYgs3c
RDWQLkFI09qKcgEG04M4yb4YRifLYwuXsA/IXY3lRvBaTMa0PbykkdMoNNbNEmQM
5OtYtv2gcJUZ91uyxa7r8y/7A0wk+td08ZfwfpMuPgE6GrndNLZ4K1522QbOmj7D
/DAnrOfUHj5Gp6J4WIkzy07K9RbO3EPmjcKxMMJM8j38wZEXqMyUtZeq9k/tG47c
jIWjGKRciTNx/AFxHWQug/VEGqwu56htF7T2r3LtSQH2VehOqYaFBoFb9v4hSsLL
nyOzyJCPebM2B2HhuHc8bmI8BA54aGGDqBwCKtd+oemTypr4m1nKUEVolfF5G9Tw
okYfo0y9af+afaZ+dkbU5n4N4cqwBWUM07K9+acRSBOq0oRSZX0/od7ADoS//bEA
pBKaKrZLH8CZD2CyiMskJIFqwCKEaF3ceZxaE172w2h23/6qp39Jdw1bb/9ZM7P6
wckcCidEREe/cG80e1g37bkt3CK5COIBUJ5QJwfrsF5lXpxy3SPFpFlg796VCKB5
ccj8W/sHtomGd8zqglF8l8TlgdDGkjrBdnqLLUf1n1/BVDkG5LCcFZatIhi0t6n5
KVKZLbeYyMma/ayX6x7ya7CfRfEzH4mi2qXBXDb6J6L6XwNk/i2SNAV2/+hZxHsD
DntvNpXX7M0ZgzKg4Kjflv19E1H63PTRD/XhmVGgOQHSksV/bYZiLnRHC5EFT+SZ
b//Y0POApzar1tyu2tIDPsCMeAffhmK8RyGkh0AYTLn6DryHMwfvmM5sKJI0/v+o
E4yYO84aXydsAO6Yax4WC5H4ahuKkAYK6CyYTBDWvrGYGvlBikwaKqWxsAjLI1D5
cxPTHB0J6wBg7U9K/YTpr0RZwfZo4SInayyruSoFvJbRlPNEIlXSTS55tq8FPzOl
kqmAnwX8O22EDwHjHax8CiOXjzePlOTYXhqg0DhGslQnqFe14OQYgR/OWqT1a/BR
xb4v0tlaTZLPTLv6lAvITBMouLLRC3V/u0LtswQr0G2LkoxKukB+R6DGlHlnfgZ6
AANuLe4CBSPXb38kB7MxbgVFvoTdo5H9VFUO8vgw1hhEQ5tK6KHt5lBE2zY1svKX
Ym7djsIWUTDgZi3pwc7QuODTNmgg0IKg9gHHY/WjQm5g7VYjvvAdwRrC3rvPexqP
ygXckZ3jMo+jS+CHx95MWPdxP9X8sDBpmxZfKkwI2ejHmlpt50cmSlFXohKd6vS8
ILw0+8BxNu0tKuGw8MI84uKMAT9TRccRIvrbxsdkulYrVJaiK3taUvI7lOx8yK80
ZbnLI57rin90zH0KtT97pTxJzzpEChAG033yFbj8j0Qb8HS1V+pMmH1xkV2Geb+P
OoEKY8enBFP8kR8umqzFmU6XNRw4ySCZFL7AhzgSUfZpmPX06YQtwNhJ5Ea4tSX3
7tMaYRtV40hz24W7YdOQXqBdltEJg73hn/rz2UJwSFc9trU8wM0yZZhtXtHT8pBp
IhwWoy7unuNMiSpynha+I/sDow8Hm4WMDabedIMacNmyrNKG3ZBKXLRTV1bU13Ny
RSP5qY8jS8z7Y4SUY2XjLdButhhWvM1MQzdbPlfIXmNvsI7GNRbAobalwPcl/qh3
Q/kfVia3bljCRyTsfJy2Bkfd3YR3w6amRfYs2UZm3a9+bfGiEVh6/05e8Ft1ddnB
DvVbxaO/pOjsOUxB2GaQ00UZME335w81+waTVWHeyEp8fYFIJKFuDrzid1Z/QB/u
7QbnG09UwljzMSqcCHoQMHNEGbEedyYpZ0/lKVQn3DdPHCJ7Mg/npGrufSoLJ1Yt
Kn2Qft5EsTMjg/IeZEidz56AkduAtsR8We5Z8CKCnDJPiqSnr0+1TDnZJYkwZkYH
2pngkUXa4qpPILyf/8o3nYNBEqyY5M621HAjT69pYqBIdm4fyhMLbUrXkNbrfUz4
o8Rfgb8iJKT1e6vPif8/l0h7sDKibUL58FmFRw4DJ/hCl1p+LWneyDfrh1UsiWM2
TLQ4qUYhoW/rea20KsjGnsbm0Ma+51qBSnkaZkkBS+b62dO6p+hgoOKJONessHny
3R/J36PaEGQvNWaHfLBgdglFC4yY0N8yCpkX3qIXotCothZNkQjYs1ZYAf+wpe5i
9IFNxmcoXVNJYLGedLEH5RC9RAhmwdAO+HZgBzuWPzreVEB4Wdo61y0vHfLAQSwT
d7tyeIySV+/pKjD7Tp5JTsTa4Tme0W6OzH6aBrrdpRkqu/HVUIPAVU2RuWvwfIQj
4UnY3Gt64Z383S9diYj3VEL+7GAqTYy07K4OMJ3sOdZSOQzppvTt3MlNr3AfNADv
Fp5NfzEIA4igYi6ZTAlxD+oGm5WLej/OffEXZEDopN5Z97XjtwGfziQCL+vSXvV3
zwGImLmV7MBa7hVSqDoEAz7PMZEnEuCK4KEccVRQ55e/COwdlvvk9HwIcHkTCNdJ
Bxys4in1IBG2gdRaspViK6HEDjAC1ghUsZXmw10dfuEQVrNlmgoR+4KZcMa/2l36
PIf3MKjHYt5s76k8qlRkMJssc/UjwH4KOCC1cX0svn9bxR0NVwV/dJ2dANnn5iXF
S4pBsWqiBDPOfOZfWT6EtptNkm31I10igYl/fuLQqKiVHX6/qVWRCPpBYVenKsyN
BsSD1Zaibu1R4xtElVwsTgPnQYRFsoRB21+9srb11vsXXk9eNZiolMYBa1YwQplj
YLmIZatsszWuCQ5nywrUYxcWqWVHszESMjpYEKy6Q+NjufPlguF/h3XjzGsgkwAE
PBN53ZokAh0eM2xCNbma/IFt1lGzZYGCuBvtBuiiDtSf7DcRF20cA4XexBh+A7Gs
Kv8hlcncGi8X3On/qItVR596/xIlwuCzC47am+YJxxBVai0ZXaPOfxVL3nWvlud4
2N96nwCqK99QWxyo73kvySsjUqbdFJHer2FQcwj6dVUVk4pZ3aqdxa1+9dAi0DTl
aLJTe7yfwhtGC2VuL+qGBkkjvoq1pq1vEXY7R5MLnBkyMtmuZO2mbq4OSlkh7kgC
bkFamgH54KBp5VArhQyzqhBL8JPsKje4RmmEeR0fcUKlDjoTp5cDB8ZGZJ1wx9bF
19Ca2rQOP2KWB6wsAaKrUFBovIceSsXMJ8PjJ8ebe6AzXUEZmATno1n4TDBxHpDe
iBIctaGCQ72rZclWOpL43caYtLgPGj8nMtyq2LlgSnULIBQ4IdHv/p/FhzmfNikZ
+mwV2NiAGVWSQkKabZ7p/zf0pWvCN7UziZcL8i+ZCdC8S42kJDvYYcCfnS6OkItc
WyYzdJ1bVpaiz5Lmm6c/uaY5d3djYAQHeLttA9DJUc+BksdF5lwYY/dawEMMfGpr
YXBPhgKkVh6AqAlWBC/Juhr2j6GsJH6LIKXGpSZvyvZOUBoqwt3tKCTXTpfKIff7
0z0q15LTHPVVn/0aFvihRAtKDQYm2cqVTL6np8dB2/3sYmU8WVV0/otQyuFqppa8
U3rt+T9c0NT/Uprm6kL6MKbO+ong/YJDqITb42+ROe5XfuQQgX30F8njTQXc+92E
jf7Hs953up93kh2erMqoeK4yd7fVLWS/oGzocA2xgPVfWIBu1AcU5GMnrDJlT+9j
8wN5S+ujBAKW+uelIJnob4L4A+rSASSAYZRyHOdXbJgyNqkufvsf5d9M67VVN3IL
ODnkRew41SfWqnIzv+4tGU0sWeqVAcwoomUzjxJ0atVxgXwoD/Irntbo5Jf/QJXG
ncr2cfIAnJjzmjFvtdBQqbK6cBVZ0qsBngbKdGJPgR28t3fR6yGlqDbqcsrMbUGN
xJCVy1kIUTSBUDARysdUdVc4UAwYmp9lFbFBoEKrNMs1bVZSZMDqiIIqzQ1CKN5U
6gVpmhYEbwLRSpbBJkNlb7fgPZO/h6jZ4mUfXVarZD5huRB4EoRuiE08mD7BXtuD
SUKx0D1Xy3m8pMBciWiWhM2uDBBTr3fHFw8AaRqCePGYKa8800XS6PPe///gjhBc
r/QcAIxc9PyKi9GEkYL6RDWr8FM4mLfoka4EBEpRS74lDRyaYX6aPQf8bCRMXGvO
MWs15holztdfT+0UzFtkErZp5c1YiLIJex57Qgzi0hLLuRFZFcWgL9YAuhJaOa3M
H/mxUW3ERf5HJo4bkTuo/aezTAXw/xRgpChnlS+92NNUzlcjFHpApKjhMtsdyPMK
aOkXh7rFWTJRj0zBS+EqCUt2arU31dd43BvNiaJj4GAOFahfVcNun7Fca1YuvSw7
2bfJMWxNxL/YSmPCx8wKAurlewwR1/FKJ/QUud/suFTocYhcjkek08EZszhbq+H2
VYgznUOGo9Tn/bu7QD4IjDrM71UAT7cWdwIlneHEQQ0FkQJWTXALicBfhltyJW8Y
5zp+F0vk57LHjWXOy5noQzgGjYz0OLn41hQFGZMT9X8TgL7INfuy532eS7AhsLsJ
aRPxe8m4PtY5xRkNlIt26vLFj/79UBSMFUMNNcclbc7KqJmDn/gYOub8z2zAr4kC
QmR4nS7gu/E1zFXDE3NQI4dEfrOnwMdsTPx+VUS9CsWS6sZy7sxUHY9iPeRIrzhI
OHlzpiSnzmb8vlgXeBGPTUCUtro7y6ZK5GJ02jhOkK2Sn1xzHQNnh0a1lJmcuL4V
Ss2dUMeUoIfGRGisaMfiZGqy4s9A6+Wz08xaR2AsZhH44Sq7TeINsmaDePQAMU1J
/sZvWt56nZ4HA9zNlMlMdeXXz1W+VDvIpXt9fslsrbLT9HXbAw5iIB3tOoEzFflw
HGeTAhUXlzLnv/a5TFIX+9saTmA9YCgflIVFuAut+qDPhI1jpBWMulvHSn197bHT
TTeWGZL+klnCUHt2BX+Jbl0ywtVoiV0bkNS59n/urC7TflCx+WCyUVIOPNaUAFFe
L0WHf9rfsx56N68vXO/asbfoBqMHWhBmrw1f3r1flanZBBHJKeCREdpecHpH7BSQ
NmitQqVV+dEcFUmfrSv/DQrH0KjYsmA8FrZT76NfsTMqNZkB2qNR9bbiYIzRRj5N
5eE7qlpRloIRuV6ukTFTF9BOChuKZF/qvWJgpIOJerohCh0DV/PL3fREOK6XZsqQ
qJ+H6Ebsu1cXFzzmNYyQEByI01YINQj5qL2csGMfYCNriQjBI2m1fCHfATw1Ll6y
0IZJgO5LMCG8+oMOvqzReL9k/lzHXY/SmYgLCoRmg1PCciNvbnEOmhtaeHYyO4du
WC1uL/+XGqCv55jxbxCFEKdVN+FiGPOXvAN3n0vqcBZamcCMnSQUrDJLbFs8UlJJ
sSzj+JCxT8kpr3e36hHiB2DTB2Pq58OdLcnKz+GKmC7EL8a7L89R+T+tSPnX6QtR
7T+njCXTuP0LxYHH4Qg+vVQo+ESnpv3oUwl/AA7WguVTRBnOkAmCJapqayirokYO
qvtwlllf3LpV9MKQeFH3yDxyoCJTMbruJ5yXNnZ+di8AVMu7L57Go2iND9LzqMjV
JFIsVb7B5k089kH9ll+MUXOYVyAOEksiTkD4yt9ro/JowAUPhcYfU8YuOb0C4JCz
SR0yGwDUh23lTuzRw3/afNOSoEhGV/K2W552fhdD+gr7pLBbKMdDPa6gdgP7rRiw
j5Q+yeUWV4ELNi/Jo/896NxDm4aMxhXn/SUyAUmG/uqycdpxyRc1qUvNLmPnKgAO
l6hRTUjMITO38vDxRfIkzNF6mw15Pmd41I2POwoT9w1H2ur88XuzvaeILyL4osHD
LefnK2YE2e+WgbYDk3VzgSaitL00hW54nczHWK9WEgHvtxfsie7tDGAIAPNhv93g
xRYhzSvtGXcayTMwPCz1Uo7sXrtZCDj3DXPwdHaYJSCkkIMMuUUvvn6i/TUmba/R
e88HFm5CcVVnxB/RD95tbfW0AOKqDynALK9whcB8rTr70dZIm/wZURo1Vjy6yAZf
AGgCKUoCm92TYJSLAeFkOBuxzqAkD7GS+PiFC+ZWUhMk+9QV633IZdqhT0ao6sSf
wm3PNwevTPnalRuy+nAJadw64xn6XkkfZJfTGMdOUkAopjENyqpcgWOIaOXM9jec
7xeDye3OWgsoGFwRhUrbhn8NM9AqOFFt/jckCqQOtUPkHAPxl2dfB9eCeCCDbvCc
gQWBTpAxnIih+HQM2I0Qz+E42PEjE4GFtywFT5XLAQzFLQqVTeY+ogVRk6STTIdH
ooV9rZXVvXr+Uc3rbHPAkc/0/LHjs1pb8IfjP+o04uVnXHxD3jFLNmk468A8sem8
u96cQoZObW3BCc5+6qUDrCzgEDsbMr10Kq+U9nK/BPIhsFqgB8Hm7aEnm+BBB7jo
g4OVwrwwwu/FhFlBWEX4IP/6nAUHf6CzYJHFRTCW95EyG18y3acwr38/vSNN4ZMj
nP5UQ3l08doB0ugwLlxwWATGxa2lz+ZJJk0jxE1NESevNoALf02Fu3yqqD1v7XZb
gI7Q1rPSHwlI8AkpfUxautMBWmoj/wOw60SAo5Y+xywNfRneRCApZO5sQgai47Qs
4mMhgeEKQsdIPT921NrkpcTpTNkLRZk+n8Bn2rJwG8fNofUvdQo2FuANwqfC3F2m
mFzlucgKbZG5TkNTUU+qEjmVmevJhgXngI+c7f/sa59dmyrJcZGu5Kov5InQbOxL
hCo0y3/o0P5dlDSux7rkzMebnTULLOKtRamDBAban8b8seGcXnNbbK0xClx4Ggxe
PEWhdACCj6ZifdqwfnoA1h+/hdoUDforhsnwaDBfLAhsrQF0r6i3tuergqB0ThT7
brpWvLNSwRVrkNuUhtwHe4HAnMNVrCYUcdVMnhVpnzthhieBg6MacjcOZI5ImvSv
OvAG0DQz341Gvf+ycdyi090FwVBU13imkvsRS4D5dBTRkrmD0lSUmgA6OE/vqOJG
3Gb8voBtV5Skw33gk1XDv5eneyrKnS3z3A+kIUE60vX16+ungL8PfElFlVzlHJiC
r/vsFCmTH0ecWLu/X4cAB9rClno8u7O6kK3z3gbgkTy7vgJBZSuiTedlwczNgjSi
vjBK3ws85/vpU0xUa1g6txuHWCSsRRPhXFFx/Dsx2Xin1o64uZeBOUDSn0KFzEsV
uYdsWiehQ8AxR5GH7vA987CKhfXQKKZJfmAdprQDOmx35bLqLm7avjP9Pz42lgbH
loZx8z/wwlIpRmcnoGgo1nSu07QlDYcY4kp3Qy6CGtSpllGISPffDRheNeL7gSAC
HT1qp93Tek/djTR9IQ8wDvnE/nM73LtKwz+t9h7xxNs2YUJGvhPp5UVnoSLBKd2s
6N3gR6cq7iX4uj6ULRPsM5NaZ7eWnSSVDSUJ9ULZQZ5qFY6MluJjylYTvHv3d4pV
1Zu9SfA94bUkf6tGH8mduZsrdw2gHIHe5kDIqbQ5BoMeaVwGzT9R6y8ldFICl4Fr
eT5EdnvqsHsfNaxeQjVr+xOTOLuFuMgTu9okUAdEy1KjerwUmyNiGIdWhlUk9Aja
CmuWM5O4unPU0TBLIcMrxt4r8pahS9gItYtVQs+DxYyuxn1+x5Bz3zTbC8YVTfdO
lMG9nCLuMXRvGDJQ4VYLYxtFEbXbaIK3f8O40qgCx6gzFkDyD7Dvn5XDclw8+8c3
kO9Kb56Mc/zovtqyNr/0iFnUnT7h8dqikKuk3IkjfURlwptsBFgb9xW2pXhRnF85
k8H7Lu11hxrzhij8mXgVGUxMVKHSpHmlY7zuxKpIrJ+0fi6XQv9qKF8tQ8p2UZUw
btUYREIXNjayMSq3UJjv5syd845uP+ZZTF87o0HpmXPd1Omi7sO0AAA0zmDhgkXv
ddfEyigiXuLkDJ3o/6J00/2AYPSyGjCBgZYXdEMlAp7c22yjggCHBh0WLNLCaOYi
B9OWW4jlaAW1w6PRWemgdki911mt8X4q+VCAJayrWxJxqVEztiVgZHiry1vqlfJD
CPZleFyIPzGxvGt3WKBKFJovbPFBfwI6cbszJKJhfzbdk4vaSg8VhJP/69McXUrT
gIFl+C90AJgWe0JnccrkF05GmaYPDqkNUtJBft0tuJq4mqufk9eGGbdQk+kGywh5
vkrPnKAZIOdOzMlYZKod2AZscqxdEZtsan3+6qI456EKMskXNlEMzDYcUxPp0VYZ
vCIBxU7xcNHdI0WJ/IEuzE1FNUc2doy6uyqprYaGUykGVxjDVVmQt5i/WBFLh9uV
GwzqyQHUQNZFv5lYk46mI1qu2ymWNMkVYn/jLmxOH8oc3+nJvE7/UkLcVchjewCu
tQAQloigKur31rt13KhQWQlqXnbdoye9WJk7DoYiZjyAseBofg9W8zLEV3p/zwIu
I0mbYph7VhmpLfattYxABGMv8S9rIt/p86CJ4vQj0o7L8SyZZU2zJZ1AAw6Grsu4
MaKgZ9KEbRW8EwIik4bbbtTF7lYSKD3Fkpo5HpYgd8Ea2KiuqArnYd6/zxaoXRGK
DhzoCphBhu+vUjKP9ZGo79b9D8GEgGgKI8Y2ly2LZS/7oeb1+xgQ0NEWNYOYHsPG
LAJTI3PdBQF9LFsZ12Eu0ANOLCB8ioyZv67G9POSqivZqIyf5J5K8heywjbUQ2sa
vi3AK7SIe1hXxucBP6fFG2j/PprIe4ubr3MRql/a+MHLDnwozCdUpcaLurtihz+9
TQ/EEDA97AfLqucJh2YkMU3HxLJY4KWSVW/W6d4WSG6ZhKTCSjMI0dt1/OKhsVUW
/yXU6bt5z2dDYei5YISoqBMrDQ/6fnGPo4YUaWLr+SuJjZO3oR3jUxC7mAESpYUR
WMnX4zF7O4B6N4S2dNvstMTj/bvKDN56Os2rW6WJzrb7aj9nOlN5DeqtCXUKq4N1
PPsbwkA638ZF+5IsnGQiXVRAoZTAtdtYMW5r3Fgf4qIrJe8m/AdSPRJdarOU2Y+M
4uoYV79JpoDjjiti+kfTycVUF3s8prbXmWDTUIzbsXIEr5w99n+5cHCZ53S/didJ
4vKglBqZDwZfeIyx/FPB683qC81U20+vpUjq6iqPugE194I8q+cmb6SaBesHhawt
PvJdKrM/Old5sXmrEUkpOdi1miCWBUFP7f99fCGok8ESKPfhatVXriGR4EFfwnjC
jW/q0TxrrrZgArW1206ybL2ZJBN2se9ucAEfvYunt0JW85ASL8m1gA98KDvM3yEc
eWI+NvxN535/LyR7U1LeUXzoVK0KJzZCriW3PB7Lrcrcet1Q9VwOpO4ZtDThIU1c
nGEIIylWvW9dKwFPMcqRuRXzeyeHkySur6f4oo4Mb7q0x95R4FBgEVZruUnyElqK
aTJjRSCjX9KYNMHDZ3tVhYPwFDriGJtU3ED5AjGE4JEkLvM53CalrQvkGElbB9xB
zeVsqLjpfhU98JAzU9Vf7IfRIIEBOrvfHEaXFLi8tO9H8Qg0kbKKAZ5HAiwAeGIU
P+qKivfX6zg9/FtQdpHQw845Z3f/999SE8I87KrDMJ8aSGVJmLM/G0gop2ZaHkoD
v9xdxvCtc7/Z443WoJi6lCEHldclJvkWQ1OpNTFASaptVxSpCPK7aQqIsVQCaIGn
0q8x3erNX0DMAPJFl1c36Amx66KwZ6QdSOdUiyOJ3VxAN+AC0xgegjNb0zJW0pj5
UuQ0y+J0SGIFSZTDrOszppI8lPO9COkxUlNH1YmGNskieu82Jln+SuzQKS1Nx6TE
SXqgmJ75aLqzQbz1nUmoTmwxxq9HiXZLwws/SPvegqMVFp6Bbaq1sVK3L66B144e
A3KCbiTKyo0TGNhKGY1LCtisLz0puG3mmJHy2NrPQRdIKvom/HQL6CfkaZuZRK1g
Z8nu9kmo6AX/IE/7jRSZLnOqRNmo/9lf19hcpq5Xp/ETuTfzDjIdo9NO5gTVQR7/
5kCRbXV2iddGbWndxRSHz8WRv6Jx/ZrtGCbDOXNob9XvyudY7BbkRT7mnWPA9ieP
WwOUWPL3P5JQJxjk0O1RXNDT5twAqQ5wZ9+2xd4usGqJ8fDGH8lf2WQYdldz5pF4
OfEDS5tQ8UJNbDsgh1t465hjHAFAnWwCLFMsJ0RONZZwuON/P6HDobcd25xqFDny
tyEBExHhTdXB1dnqsdk37hySJUxcMdA0pKgZcjQCPMOvqhT7MO8GGOkTcORpI1ka
Vie0ihE6AispT2TrR3ECxBDAgXI1j8KM0pQ6UYunXXfBsqnGZflqmgB6Qmh4ar5R
QqkOnanB8vgUC9/3z2z+vgcxSqmM2sY/oj296P4QvEO8BH+vEQ+VFaM0QYFhgXvw
pmDJ9RPHnWVPk48vGHrH2A8erijBApG7YFgG4qHZOEa0UVajZi7Qh4DZFkoi9vph
hGHnGgA4lwQ9tKgIC2LNc4FYwrUfsICkETIl2Q6PCb1H+5JYEyqS3lM8OLMeBB8C
paN8Mc9zMVJTqU5U/XK0/AC3QSV56+Rz3D2Tk3V99ZTe9HeeMBn74GBOxuNqOcRC
t19qSv9dPTKHCPs3eXgVWY8pHmPBAL42mSFpBVvlDbeX+rBpdIEY8DXlR4zuF3sy
XMhY0zFnCMLWS+ypWKxZ5PNmKBelXb1/jP56a4A9l5tSCMG77AoF6Vpe61HI9IAT
EbnU73it5fsdREHXqDnBHQ3BiQrZIOz2ZKNbm6mhUNUcI0Y592+hPwjET4JQrg6T
3R6UR2ITFfFRhDlLU2kh3f4vy+1nJtcvoJKUUdv+KWobTo+w3bklpU+ZlJoLEWYy
mw6t8txO+EG98POecfjMgd+AN2PSTW7Uz8beMWjpYIuQwF8hdDVI3W/W0gBSZcrp
sQmoczf26a/2Um2Mxz1hrl6KF/1EMCRG6yA1u1ARCnyFAsjpGS8k8R/Sljk1Kcfn
Bdxn5f6nes09D92ah/QH1g8It/OT6R+63lTy79h7jY+SrHAOpdHAI1jIA93yyADV
2z0NBIUqWqe1lIOUoL/zdYntHoMJ0994H7SJ1U41JlyHLS5pIJry+UWmaQUabSli
/ORrOqUiZUVbsQwGUf98WSyaLhfkQzfKDNQ8e0faBnMd3LzZO4zTfnhCHUofTqes
`pragma protect end_protected
