// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Cbp5gCnPNqHbGRzCih6mHUrbVU/WVOPDHlLEWhMagoEb2RgOqpVbVyl8EP4VrP6Lng79kBKliwtZ
cIG9STbS/M7WhybDQR77+EFslgb92Uo4qS87o5sZ+QgA++6NzlV22G02x1qoLWgTa0I7wv84ybVs
plrUqZ2/05rSdhqsBCnd1IDcOmzwUJMP7eXnwnbSO2AXcNB4NnxfGaYSFRfp468rXGQPKB5PPfH9
Uufpln1o4GAEjIM6daq16RZ4aj2bw7AyS64udE08Ykflc/Ippc8/ulTWfPjsLJBi0H92x5fVTJMv
3U4pWwwbUN/NQBF7b9Q5BGANzlic1dR2pZehlQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11088)
pDu6EA6Qa1LRhiVVweIWAZ0wO9YbX+SGLZty3ixDsXIjNFHUP5mZLVrJl62WjmWkw+1ubaDDfqyD
dQ7WWHoSeEqgHjbaPQlnagDd4/WOY/3y54VYXkkm69hfOhVO+m644CEKDQMMHnk9tUkOzXcD7eq5
Yo5Xn+MayKj+5yy1nLq9tdp4QzIWqaCM7q2KMNViFYj7/eaJ1GEHtgoQGfpFiRj27VnmlWzP1vg4
lWeBzhqnX4kv2k04sAlXL/VCEzW/4AFbjERQXveS7IKowIwPGTTTHBOwDxMO0aGq09JGUCqPdyQu
x8a9bNa+pQ9R4OA4Cebwo6UcFetf+38eNeyv9Xfl8MdgpTkqf4m11FWg5IGsSj4EROZ/HGXktweo
UzZQqshJgcxuWPwqNDHXCfmiJblX4j70cOtmEOGeu0G3qn/aUNG/b98LWHBFwvLNY4U/74/RULxC
Qvu8AD/S4HB1yig/otCC14uhRM/AQV4UXPvE7Zo2rHN2ORSDjGU/PKCGjufjLpXfKN5RVj4+V1M/
1vsNy0qdwU8aF98vcC7mBuvShj8r/SyCz3h4LU0yrHwk6hc8fbTQdXFHRjYVAsLs39p5eLVVn0Wz
5M3NsiIMCPWvwGM7e1DByEagDJTI/bELwfO9QMtUlaXso86WT0rGSy2ogB+b6bjk7kG1R7+lGE1l
KGsbfBJwT1xREiLGpMrhER5LaZINK3VlNZtI2EZyoaK7Zc6yyIAvXXAVg/38wUfTeAI74qlZM2CZ
n9ij0x0U7aaR7zParJ2/1rcJZHmfN3zPK6Xj577cXLCaKOsdTkVTVOCjNUueAieBVhG1a6NOPnNg
JD18mhPcaMmVQ2yiJ00WB/MQiz8zVOBvPc7XNyDlXUMv0iW7VRyPiFCimGm/L5kMLFXVw7BL5zxI
LYZguIOvusheUn7AYm5AbEJxPk3SgxBHYeIAsU71++zUTH8WueZnkeAHhc1dCQ/ZxOeIer11v8Kw
3cf80cD/MIJUkIvlR1heZG0ev7gg9WUnTMjvb+h2Il1JcfMmQWy405kC8LPBzcLYO6OGKCqSLMiR
7InKzaIydWDEdNoSAZqvsdhqvQ4Ka7YHq4n6u+z4QzlTVE4ys6ykWN5EotM/XDl2Ji/YSe/MfNx5
mJSF1epYHgJY5/YTn+mqVRrTnGRXQuV0Aa0kosftzQRWGTESCtw6rc7Lsrm0C14KQ7KND1Ep9V6s
o9qTioOlgk6CX/qdKFjrdqyfAqhWMOhYvQhup4zo0+gvlKhX6O6CO/h/RH/S8akkc5QLAr+F0AVX
IR9oeiOyaqYF5BzwaiCtRtdFwwomm/d+RlKk3UYqSN5y9e7BtyQK/nsWn+9dVYNx0S8NcgwXLnIt
B5SiBsoa1IftcyHGTDkHiwYkM23c4GYJHUHtqTf4/sIgKqGgtY0DpQvKkOaX+RXJG1BlkME2kHJJ
BR2w1NgEzDIqEcU1eCOXsFq/W9hAPi1p7jpHfBcmPyuP6Y0hgCxwZ2Am1Gzb3vGqgEYOf1OPdXSu
6Wk/MuOe7Yak4dmWrtED+eBW9SFbo9ZErVerVLllOH0BxLdrGqw+KDriTXKnl/gTrkbQ0NRwhZP1
mfVcJKZHT7eldg6WHWuPSSaoOxU3HAYIxq8Mb0+OZ+hhwr1fjovZI+uZKzZ8D72AmJHmR0PwfSGw
M1qF4wC1skwVuD1EchheFMWRpavLEDJi1K04w/lK0M26W6zFcZlKrPAcKYu4BGOqHab55Z4LIX7q
Zy+lSBTSJPG/m7UgMOJxtcxw5UVy33Clalwoq2HbHVOusGs4lKe3WVlPHoEP4zLYKbRKql18XQCT
3MfzNxgGv/BcT4wyc02wrlpsNuUClvcydhbQ/LwjTV7KrNmPlJK/natTP1VAAAtOJII9jyXP2Ivh
+0LzOirGHPZPmEj7GiH5ttD5CiU2vmJjbrrsT0JerjpFQM2hlJILpPnpCHAvyFPvvhMzwmBD025i
6psfu1+BC3/DjXuez6f5GpF/ASR/cuL/dGOMjxKSxuhdK3xArJu8uznJtp/ASQzhsZoEirf6cI/D
ieXeGiYju9QadBTzzk95zEL1gKMY8ndNpybL7WJdGBhRQcu0ZhhN9s1EeYV1Ekg3Cfavr5OoA6+Z
EK+JJfjhFZsJUQcFCYc6E3wStAgEMahTQjSRQ5CmaFQdqLsJKmT/JXxwte58jIuR46qm2ftlyLNV
8F46pVqXCTY28qEYpV1jKOvM5ydf8kkEegxpYV9IrPRc9SejeEanc8eHiMn/VSlCcfIBlqTahzTy
7AoHmzuTD5uOdOzh6XKQhxgSfNcHXP2b/8tKVScRNO2cGiBSNxhpFp8XC/ImuP7Ja8hRSQ+uVIvi
f0y5r7SNh9A0K+Rb8wHpodAmYHgkyC7o4rHiT+XfQYpUsEnfJq+QQGrUBVDy2zZMvBs5YiZ+lKZ5
FKjV7TE/fgWTJLXk6vHt5OE4L/R2yQtwo6HOj2sx4U+bW8Or1dOSLv6/PJAwVXz/NnpSm9tUpWF2
aT3+rhgHKEr/Ddx9vmZiWyZnGXG2fkMcspiPxYePdhHuwpjcTpzfmuWEvN/M8GqyQYA3l+xgdFqC
/hhrS8k5G8NftvdFssVEhTZkRsqgKCvKa2n/LfquVKaWg0PIqnd8vJgl0x3Ul7Cd6VrcDa14NDbq
+/9GVzIaLLseqNAvqB7j9KBzeXEFPJSAte7e06OBcQJ0+/tz32AtmAeiloL5nyoqSnaRvzRVm9hg
ZCWcgAIdebE9bdYhGrlozTrfXeZoy/TzkdOuVTOAf6QsqehW9rji0g7ON6KpGsaryssEDHLx1oqp
PU0M5zaBWLiBsThxrS2J2vs1/vGWdBkhpeQ9AJB0Rhnzf6x0DxJ5bHd6JyrQIr3M4o7IfvYSGI6T
WjPPNrN7/DUKVHRrHRNeAb4syNHcb6o6LNf15ZahbFettk02ddIHajUbM9WPeu5aNQKGT5lSt7iW
eFWFNDzG8LMok2c/KLevCZlLQ0Y7My+NSwSxcASxqDnpGQvIdWaBNiQXNT+jleGOubcoFWWZ8cLB
5codGZ+/966iFk4JnAtL/eD6qRRjnss0QFjy4IfJyqkbeLTDFmA56h7YYFJ3SB/12l6byRPoMXS2
lJDuh+TQKZsOltHB7T7G3wYSYCm+OOCW0IqLKGmmwstkRhMoDQg51TT3Sm/BK32knGHVeY4Xh1M4
OW4Q+0B50mosoqGFFJG2ANpB9g7DP96+L3vvQhxjZh9jd/wL8V6+u8Pfc0Y1wjm4l6+bYKiHTU4k
9BSbWYQ/tE3fBu5cL26tED3iCcaB2jmhSrx2tUDtNRxmvUeTtWBk/dirZT64tQoVJ4V2Yz3od5n0
Dn0TcwWt1U8DnpfrS4Zt0QkK5bo8UDBLhgmaR1uMkngAKsUUE8k/64oACQ9Eiw4Ef3IlF+3sKQ5q
cDdNdx9eoFUAE9KmytsmfLQaFNN+rfCZSwEIAl0oAqSE0cfWJCzkFMA/I36qNBEiQeS/q1gDeeui
kbust3UjuOX8sQV6VIxnIYzA63DgxVEMakTI3omCgC8Gqui02psy/IRdCnJJVwG6zK4qz1va+CQn
Q81bllfZzY1KePIH+UauuEsR/nW7ZumkjdwZXQvs4yDs85nS0cP+GfSGicKxunmFObHUPO5MDLRS
56k4KOWNYS7IUpT2dCUwy3VuYrr3AS5UKgEF+FWy2JjJjVB3xMBKIpTKjc0A9zbjXwZHi8jpZUT9
89bJzD1hEvwg+ePGpQBPZYUrtjbb2rVC5B6PU8gBED4sLXFFIyZeYyc4/Dx7BrBHvwlbPeRQ9kKN
n85IMIkUc8+xwhPT/UFA+X8sIR9gyfscvUTk8Cq4Bsd8hlyfRNt1sepF0PmrQVIzH2C30YDJU+RF
EYAH0ovnqbbNxOkitIC97LOQO1DC41mcZQvd3kNpUHx30NO5VbarOzhk0Zr2poLk/RL/4fwqiGt5
kOOc/pe2D9wvEQ01MXKYjlHmS8AdtK/GGrLZHI5hVcJoR8Cz2zdI06KigmUHnznl4FtX6x43Arfi
kBssACEc+U5uZaeSTbyqycNY8QkZx4EH7WCQMRY1pmx78Jniw65yz3wV0FGyNQTGhGc+y6g8p8V1
DaIKBzSGYyubUYOXNN3ZD7hFqQevkjqJSzyiw+wSPGKEg3Gcm5jGbmxTxYdV8MqQwMQ78XPrxBHI
JfNAgmjifjV6PhFBGUxThMYLEibdn0uHGR6BeXIrUAHP1ETzvZ5wkLgSzCfQJEhD7OcxZy8LYowN
N0x0xPRGEYsnU2FPWlQozU54/204mAJwGvAVOCn267+t4ww3Kf48jM3TuqdJ39iwdhqLIjqFKrHK
jk0BRmbdhfQvMt1IWP6jUp+bsv7Ya2Ym4XkRz37isrK8RoqhL4I0Zw0kyRSyMPMjWostKn8Uzq3v
tU9YO+qUvOTg4l5uQWbLao/kBMyTV617rxk6xtiWhX3oeNyO1eFCHSjO2Ot+g9jbXLOB1lcHWaMK
nTX7gZXQ6STt06WEcj9xSuysYiO+n0wWblO1EK5qvxuhQeQtUkrxSBKTUUE2Xru663CCwp9a9lc5
n2JdV8dA0YhhyaHRv/IB4HfNbddkCanHxwHnBwsSMf2x4Zb9o7PHaCgAiHURtx5KfING9BozfDoT
sGBmmHQAbTflJervEn0o7ccn5kuWxcXBx1iMXrhmNLSzYfSeOsKWzg56VgObzjtdUOFKndqyS0rJ
UyEkXD9xVTDedrcrcgBfvB5unXYej/lCBNt9m3h70h+MR4nIS6UNwHIp8HPMhjZTLu0BLWm6GOoP
bo1WlmMCHG8jRcDqnmIiMILUZyLXSFILeajsRNrkeHHr3rkhQqrcqjmbRXA9fMKiqZNSAyEeaR6b
YUx2zEYbG+PAtZaz+DG55muY/1cMYpllqRDCMpM8SY5vhmaH6RGf/laLfGKDTNGU6O52FdS3yMpU
qW3sC+405NiwTrwx7Tdtq13TVCAeJENckyzMgpbbLOlypDjTvPnwVJqO+savDVSGrKppw2mhE8Vq
Nz0WvcMkEz3P6HqQfAGzxWBHWaZmoUp3ehPbBVoVpWve8U6ea+CBhYpkTa7+N8JzHQd8ABa25+1U
VdfMfswV7pDTlS+tA1sNlu9/2g2ideY1Lu7uqgZWwNI7LNOAoJ0CYeuHXHVTRnQgRLhhLs8x+0CR
UuZtY2gdJzKb30SC6CCqQF/pLdrSOYGs+mklZgOyisynBqoBLB1qWm+dwEApKUBxhzV8z9CVF1xa
+gBJLmmdgbqhQmLhSJdQU5r90Iy3bJ/notRfVYL7uQ/Z5n6TiqBEjUwVkAoPHEEuhJ1tpK7RYly+
7Uh65j96Y+x5Hi3neGrblCzce6Knbmfyp72iAri/Larx+1pLv9FdXzR8eJYBdhSFqaUtv5tFQDZK
emP2Kxz28IEeulDsS4KXcK/NHUHkZow53tdjGiex4BhGZ3RcTcM4wI8FI29jxOoK242a7n7Ui9Ee
fm/7WaRphzljg1KuI06Kg3ObEHEW7N5rlqXVV+2RiQPjiirdFDDZiVxb4K25aEFPk4ba0V92H1Iw
xlB214D8OvBfpMCgmKgesO7quHHKJla1b8DoqMuI+y0LfcaQABpRMLAczelwB+SnTsVBSm04E7Sy
sx6+jH/9PlzfroHfdoWu+ZPjS9x4oB5rItMtKI5Bo9ZYBpAJofKklR5kVK/C+wQB4eyMwHiC8UU9
Nma4Htr6WsDf4wa/42p7iB6Rgz4ewlfrCzP4bLjgmnIRyk0RPSM/nM/dzAxWOunM5BwlV7mkbNwh
aFI8ecOZoqyVN7FQ3sRC6YTpTx7SpPxCTlZ1Fs+oZZlH6GxH0MEghUL73RnYX9JhUJ3ZsM0nznPE
rDixRtOTHixiBJ082venFrCPluIwF2QyaMUsHRdatpaIb67ongek0+7U36b0+9lBglh6pe6QFbEF
EygUO4xJmkpr3zpLiQ6CD+Yd0sBgrT26t9+nbcdpUobWstEQjEbznHFlOuyWCEGwWPjqqE4rwU1x
ke/fDgBmF437fAa8B6VZwHmBQ9dWCTcxSEr3+wKQAKwK0FYoJuEoyS/wpnGv+7t4ru/zR++OLrsQ
O9utIPU2GDYtBMA/gWPck+6LE6e5mKMWdggrAFx6d6EEx+7hHS4XWAaeecSp7DJ0MvcYOYZV5eYp
gvCPvCkgOrq+2Fl3GrwWMXSPlg3vS7E3hhWYL6kd+1K8jDkmdg96rN9So4YXlK1tINQ11LAAqyFr
hi0fuqUofua7TA69hynGb7GnbnvlHVQYDEPvDZDLtJRin5Lh5snm244tSVXsii1xaVbA1/uuwHKf
EuTor4FThcKTd5y6bHUojBh9Y8vT8LaXr7r1i/QKZDwAC55N+rVcUawvgFmJhxvFv/gf3910RpTY
wGFTlUDR8zMGsg6F5r34GUetfwXHn8pOLdNXAVkZ3G2pwxMcm3QtvW1951funJ7pO4Nv1S6G3sPc
e9Yh5F5+WEnTHBJFTP3JxC5rjrXP5/9zUNCgdoRMFSmEfDKB79BUg5ufXmqiY0ZgVl5kYjbIs5wU
YDkEIApfsroMFcB6+f/sBevllL1jY+GXA+J5Whw7LK378xXZDM1QkoxDHpGRCZuSsPzlXUHDsGhg
mXOIZOPjqn+iIZ9/+IN15iAod/UYyMt+n4jhD1WKG53tmUmreq7z/ZeSsDjnRnUR1iu99QYV5uQD
9Zk3jqQxtqN9VBd/B68rOzN7UqpHRXfMd0NfzvNA0ude1KfzsSB6HVOvr2e6F29USbr61EzhGeRq
AUztt+Vxb9iNHa2U/RtTp6gMGGSW6xC6iIjl3+pKEvpOQjF6VL9yxUipv6Wyjaw3JPiO+g5cXAdr
VY/LvOiW7uUbonUbviJNDvIqp96mD+P1XJ694fjk7kdu+sd+z79b4rDQTBr7e9Ep5boxc9vnjTpm
6tq8hpBJvGnJW6S6Z5t0of2ORKosTGcsH7lA+wyaxjmVs1jCWNmvd14NDAH88bmBWrGR+zCysent
yiSMd+Bpj7v3mZ3gwYv+5B8lx0hhbd2cpOyEWWa3wpCh86Wa+OENsOyrIOBDfeSR1vxtXEerNER+
SKFtnmymNQtzILA4TAy8eoh0EOg8mJPtLqJLbXkXysJyij07ddmXOBCzqmIGmGZKhSB4Gep5+pBV
3RHzWykV/0L8C4Imal6BSi6i3ExRMlx64HGR0BN79GTFUdoRsO5LJks9+uJIext5yJdq85QFIFP/
VG5MyZw1Qc1yw8v0cXRUrp6Wofy5GuqLKxzSzzt1dPhOOA1JJVWULHWBPvkECri9kEXzoTP5PSRn
t13gjLCTrT6FT8n0SpARGoKR3tXkDmRtufcR76yRo2IIkelaAKLKG2AmCeOfATybutGcdmPUmQSe
2aGcDdSKK95PVdqH4K/FCc5frAI2OMUVb0wThT5P97KoRbWwoxHsjrpvfu0p6C3Z/BsE93zm6bMd
74KsEmEbTCU/mifMoKCZ794KR7+4lxN3Bf8OyMm+C/3LKdqTFH7Uz0MdJm76x+OmdLvzkmap2Zd2
E+zVSc/UKX3N06GN4M6eKKhQh1SSxxT78ST6Mu37iZZUmNlMsf6tPvV1bj6tbOk62Uam6gsHfJNB
YcYe8UktoStCrQ60pJK+Yy6oXI9eWtD3FG1hZz6s4sMNCnkPTYAOv/d30ThDped8D4JSAIW7GJSW
XMYLm40QQ18Riwg+zn5K6tH0cMYOhe/m+Ff4wa/43fyN8ql/ayPfO7mTULLRwU4PeFAar12d2g1c
0JDKXpleP1a5vWebrbMq/4TBW+O9iO1jKcMGyehjakW3fBNqdb5ruV/glLrbzRgDDJ8tqek7M4s9
X5u/yd5jPl2U8qcWu8jT49Fkz7KF9TNgvQXrotD2IPaoJ/ccmzq0o6+pxwuQobKxjtszpEXCHrVC
RkzajbhWjuqUzwTR33sK+omnsiXSrd3AYGaiPS1EaUG9KgbPPYZ/lr7SGSyD+xWY9rlWZEfXST8y
4CXl9nXndNNf7THwWOwoJ0EH3bWXecM2fhbdvzMG+h6M5+tBs9tx4Jza/vv7626EYgxJOV1gNuXh
911pIafFLdVYBpbWBn7rPhxJ8owBNK4rWO+DI/FV3Uy7ntB9tkFEzuHQN1O+UzusYhizGJZZqpAF
gkeZyR/ZnF+BqEO03hiHJq1MXiTx5hSAfYktx8rTmjfTxGbyn1FA45xTQAAFh4wRZXVhfr3ltPrK
3nlG0Si5G8nZZ/5jXpkY1d7lPt5KeYKA8j1T8YtzEzWaF+CnG2uAyM369k2d0WhRi+WHrIyF7UZT
wtWF1VXhhcuvXNCoyfc2ELOBJrDonE3fF+NB9yWAr4wFJ9rl10a/peV8feAJO4QOyvSf0t63yiAp
5bWqfK8EtMcMul0AXeJorAK4T1lIcZkTkHGtFRN/enw16vo/qgGdTLCJPqX3MfgRi+1/yDHx5Z1U
fGAKGFJxfQUVVvnVLSO/iOv6RwYa3PDsmk6Ugv+d7npZwT+F4tLvd6AgMwVbQtyn1stt6KCp/kI6
IPFyGGGbQp+ylVD0QFL8gBD4cEfXVL9koojOPY4wSKrj6ftYv1/pE0WnqX9ecZK91ojD/GBIqPFD
ZilY6HltTTGlDpafmFPsoneKpKSBRwsTUBZQjkB7fdyTTEUIxvGdygEE8NF+ypSZJ8z3Qwy/yOdR
vpINz4awvz1sn+k3UayFLl/fyPeGISDDk7bWG3NakipJNKviPKn1bbnk0kycTWgWFvVH/pXQN40n
Z2THJH4aI6qvacFpvgg7NyWrvkTSfnNNZ1hdAvQA+M/wdG/nUaXK2Q3ty4iafamLpXUWWueecmkC
JjBwvIersNRiWHsp4YriuQp+pEa3sDexuKVXi2eQWEufBkwqpSkLRWPuQ77/HHszwz6jsYaNrsqz
U9q1ByNBaNMkUHyf0RMkKKZcstWWFEAQiFgNscYdgsaz23kWWUNiS/NA286+SG3ftM/YogPcePqB
CBoQVlkXeUCpfUW/+XFW1NBO5o67PWgVLgyMvL+5Nby2j2/rSI3PknGsVPDpiC/D17sfRL1Nn2oA
jPP9Y1j3susqLdOZgQDAoIsVOLvV/ve0JqJOH0t0sI14vLDf+2QC5E/xHlWpt5WUvSq2KuGGOJud
6HqeCh7hngrsfqIOx6DhUKhNWPjZN42va6E+uaxawnf8gTUAkDD7X1EU9huxQhjFRyoIZkHV5lC3
q6w9SmD+0EQYhDlUOQb1283y9FQzWLOMRwn/sd3Cf86SmPwI4vqNFLqRvxl/olcvsralnVG3W2nw
oMZLWr6ZNuerKkvXnxibSyXSVLZGyZP90R4WmS0txCAi4OFJcgDxkWTsuAHFQerTgbpBzoH01oSp
K2y4LiiNZM5mbkW0pOL1SueUdFV+U8FWG48GAhoP/abdLxyCV8r4FtkSMlerZm67UpU/f38bTz0w
JjPCe9gBVbU8FJw5A+aEzbXX862QvNnyUHj3tleGu9vbprYwfsOtj7Pf+iUs7ZzKlrVo9f16GVht
4jBrOR5vzOj+8rnvIfaaId/K5aznQrBUscBQGkElgNija2Nxw06W6xsucdDWNoeAhOu3Ev9V7Zly
BdlBvzoiKiHAK58r0yruFFt66okh5OroGKRKrgeBaCiF0v2Nz7puzCtnjlGEJSMydiEzBPqKqqQq
X0DksFRJ5/cwUkf+GsMGGNGzNwwkUvD96O5TEO3LMSnuZzXzrRDPitk684llCEdAyj3es9E0YIGh
NEXWUinYycPtkf4vOylMYhaXNCMd0WTSPoR2HbPP8YDZlpKsUG9BIfD2aIdCEdW4XPDKc+LOQuTa
xTWan2I2oG8IcJyK4DH5ERkS9tRY01Mnd8R5xMM5TsH66pWJOjL85bhMF2PxtfpGT7RsEPJagqi6
LMZvMBD6H99/ripQpkqfPsJjtq5k3DaBJFbmFDA5eh0yfsW2EAIpOFV+4UYldDo7JJ7HsoxOhaDf
n/b7fS0fbPS91/ikD6/XWKBkVsg3UqXJOKqFWPnRsMVSbjRdGva8OiJKaL2fog5aooQyQv6DJ5kp
rcHPpj4p9mJxpytnKmpzhduk+rHPom/YD6x7eav75exl9ohHt6/JQb0Iq8YsB2E5qE29tYdJQjOe
S8Gq59tP3yeaBjxC8I1xwYgLxceUpr+Jic0qfrwF3ebUZZFwzy0EjuDF3nnnA5nWUzRvVl9/oDx8
j4GXafJrK7l4IAiMMqBYJXGlr2h0C5iE/5c1mLkhYVvAhVla5LofOYV4iVdL8S9Z/EADCqIIUEni
jZUY9RuBH9/cfNc/VD/eJHbamn0fQHa3eg443Fzufm6NRH5cLOCBrE6eTXRDiznwprH4kkhXdkcs
xXdfIWngJLw3zLtPX7mKTxwBFf/CD9nyOdbKZJ0KZEy5HOsIiH2l+6zRCo1AJeMXuW+sjAaLDmTd
YOobPfP9xlMJCgWrpjsJjzm1+xfL0nVMwC2m+d2QruqOV0WQt/XzO/cpNUc9iBdGCJJ9uSnYCJ5O
tMdMgKtmRjlkdGX+Tx5GM80x1ylij1EZkmkd7nXV/XdHaR6a4X6ay+qBiuFqIjdB0cTunigf2gyi
O389I2yBJp/DlR82Kdzh9DAS7ggasW8yChRZDQEnN9Yxvboh+AqsTrWlrEzx2rsn/ibHCSx6RaqQ
eVU0sfBr8vtiuuUR9DkOmxeezBUiJi0+DUVgC+8fKsNzi4vpgtNeTFv1XDEbgl60nf55BvJjuuD0
J5Hz8feYThA66IgSo213vsA8jq7Yjm6zSui11C4wVkXwkvDgXFU0U+gwvVm5gO78A2dhEax/a1LZ
ir0wRoEPOrwbZPWJzgeXb/z4nLWUm6fHlwrkeHaAGkMh+M6Li6fwy+sxnjZKb9Sh9aOyns4e+5UV
hfmbkRKGq6kiGDCxDqy2a1Y0Hn0+sdI14wCwqT3Nsjepr3rjKmfUXUqFTc9uhEwzEHmL2s1M1lFX
+v8xWtA8fbTCUqQufCZmpv4mgz5lY62b4FLVuG/EaN4y6QFePxM4/0D+2GqPiHXpvaUGPD4k5hOa
7LwXDLHbJ9iRTAA+OqoDKIFUXgcafjfyezJ4DxaMgzII8pr/jxZenOUMSN6/1hvfvBYpeX4LC7cp
VeOuzZm+BUORdiIyepVDpWyjJ7PtD/vIkQaOcBmfhT121UsxgWFvi+6b6DShDtLEuOb+RK5ikMEt
6+4wtJ86BxQ96+4N+Z/i1L1gGrDdKB45zB554Of0aPOZ1s7+u60m3Ri/kgBWPFwlgmL3noFC4C3a
tVSRI5UEZVtoJhLcK58BBKajs/JFeWDDwDDopcMakA4cHq+Fp3Bj2NcqZQV2KQ4vatQnebTIYeC/
66Mqch4Yu8/UPEZ1+5ucEgYhwoA7buBrVPtYymPEma5Z6RLkokEMcV2FaFwBbCgGI9I5h0uofUF5
/pwe2NOxSUplncB56DTjgD/vHBUNUbkRni01e3QWuzmKIw8qEF4uHRKobtpNiZFQwfx+Se8qwiGY
7qDtBWVot2k+r1/bnx5Dfd6wa8nvmEYAGkto/B2hz/anNegYolgpIrFuXnLWhTAfvYHX/8DYuEAn
RUVxXJLCYaTzjFoWUffnQMhU/6Zaf7fYmIOO5txDEC4SC18tsvoJY8UmnAaQ/dH88722I7qEWJvk
n/AeLwFQKcIdqEE8KvagexovKvXDXLky954CiRPmT0VMQ4ewScvG6t8PUfSbhu1XEkMB7oboPl+V
qRgsgJnGwQ0Frk2ObyiK2OvaV174FVoteKUN1t5YtHzpvaWk2n2G8E22REDtIoObxM7zBO7UYXw7
lZfM93fE2CfXf6JdiYEN+Cp3zPBlaRXfXiWcfPVHwaNDcafqLqu2uIK5We4EoSIrLQt2ClOgl3LN
yPlQUk5S0F/QiFLuxxMuEtQQdMDzS69iCA6Delazl1QPWe53W5c8LB7OV+cerWrv7y//gAR/5Lpm
gmarr7Vo3x9OuIKiSx9XdfC3Q8F+Z1oxfcH8TYEgGR+HDB67pcCMHzdVzf7gIX+PV4EYOeIAZlrw
S3Rkp6NNb7EroddIdlKdhPkiFgbP0AaB0iSqGDbrV6dnHKuHTjoMZLhOXguqJPdnwdr/TE95Ip5a
rJAAmH2+0SirJBKTk1FJZTdcRIY5/Xj1BJ9yKxR2GaucRHF8AaLwhiRR/PtzZGbxZdLnd5M26pIr
ECyTMlAnO1E3ris9EtKBqZt8BqUrCt53jCc18tP2KLAfklrN0kBqIBu3gswiMRB6hAaCgiPK7GPf
iibKoGVDKeSW+X7Cuoe/J3Godit41BXP8+mxWTjsXI2nxgx92J1HgDJEA95hjLG/gEh4RZfmGOxL
RRh1z67L4gmq+AXWtS2IuAkXqssx8SLLGDy2Fd9ZISvKB+RAY0irPKWX32nWQTMxgfX5bWiG3OXh
iqW+b6yrEonVDCGby27tG3LObFPvyOxI9k36b6Hicgyhamc8wRjh3OxkP6KFuP0M4y13bId4qjWT
J8q3IOGUy/t9NLq8p4Oce7HefikR/FJYmMNodSlnMmB/iAuFNJCngPDzPv77Ujo1P2GBrxMDEpon
nDQ6xYnQ/SsdOi4Ejppq1AjuYVFDFjj7iLWN1BOF2lb2r48lHFo+stzXo+W4iKlyFvQd6f7CqcYk
kKWI77PTwQuuwvdb1l7OYEfgx1SFqnUjaR9ZHIDtHskBEGNJr73K3razIM22oJnOXQct3M3z2WyA
nlQzwKyTi43afiF9CSRcWrbtENniJrJcMlzd/LQgYqVrQwHThzlUfs1+OpwaFOb02ksp51nWB5Ry
/qqJkM3PqsYIJG5OfT7HSkmaLdptFhiUS/K6rd9BFoPlGbmtCi7ZCdEU+HoksQe4E8mb56Alw7wJ
/TMY7IOzYHoYuyKnSWYyXm9sdJwn1rj2w861nxtaRennmAbwd1GcU5xZIsRGMAUBPZIfcZENwa8t
b2sgik0dyfxmH2kbfa7xl1asgioxbbmF7H0dj/HMgXZVfYRyDKDzGOcp5QzDr+lyXIH0M4+7THox
qlKKT3w7WwsHtdKg5YDn6um7JssFqS5kP1hgoV26Am1UzWqhIVs/9tqV5LrkiNXckjuNP7NWjFtB
G0knbJCAA9uMf8LWu+ISz6e9eXnrGsPPle9DPfdkF5ZETAZioh+q7MfR00w7AHwIekUxiIeNQ/bj
R7EcKlZ+X2vbZkB2uY6hxkI0rY70DAeq3zymmU93cvf0xVoiI/PVJ9ocJvPueRkTW2PFBfO2zs7o
b7KirFP+/5/XgPnWFkwgpDBlvqk2BhRbalTOu/Dw6Zz/za16NbegEq1Q8mGPf8+6PHLyzEzgWMXK
VgHMBRAibSohzq2c3O1s5vuGm8uawSIqK6cNmewN/A3GhC1an8ONdMQ0MDVnqN6kvAlJMHmV1AZm
cSk1inJsdl2uFZ5+UOEdx70Z9eg2t++ENjXnCAstU2XyftXiJe6zi3CQ47WkRn9MMqim/UamZj42
gGdESKd3IrqzXltKXnjaV8ULSppq1E2D0l68U3QR0DJxJgqNltWKkM0ACY9s9ueks12zAvcUrenp
xneux5ibQ0P1QH4+3rAYfmHeuWtmeGmb5VAQa4kqkSNKQpD95gwS5MpPv/J04nFueJ2e3W/Zkm5L
ln2u9a2yO1LZi1I0sMfG6+P8s5I6UTgA5r26L/KVXbLBYAlhfnRckDAEuHKkaErYI9gbYiUa+0VB
A40dRnRJsqiMjt7V0B1y+rOrG3rZ9GDv6rLuow9DWRFzvkTVBsYBBIqpTgTTUkfBHUN2E56ItSuz
HtOEbvJdeG/8qLFpvY+6p7WNmZBgYw5t+iwUo3E4c6KyFqXdwGvoy7aZ+oMxJ7Kc4fdRhjWLWxn6
Hb5inITr7KSQb2MfCuRc+qE4y64C6p4yXrM7AMRvDV+hclNqnumi6PrskRoJ81RGAMzkVxBtplb/
elwEL3izp9IyNCYtn88iE+WDM0zwwnmY0nQyigZpXy9n9uUBFeKN9TiBalpFdjeZzTAKPnZ+7YRf
H6Qh9IyRHnkyYXyERyRFABv3Wz7az9+ZlZJzJflwMSq6WmoYlLfF5tbQAYtyBLpx4UPayHg/5hcM
fdqkau7m0FTs70zd1VF5/rU7Ra1PW2hvj06cyRoR/F7IelJHOqQ4zIDtQL51QxVxST99arj5z8g7
9iAsuHipipZZ/poqQTq1Po2yRSG+YkbKxs5H+OpF9ryuNcu6a8yqTIFDQHZJIbZPned5Nj2SRu78
6p/MURFbxNy8H08GTyMAuGpJK0BltxOrItdapqAEe5pQXnemTWDRiWTVuE6YXdiPFj+iBD0HLBy8
JFvNmGaHhs8vOZfDY27N2qVKTX1ER70y3TA86EEs1mfmEHwQiBwPoiKq3M5OzmaEB9892RCYsJ/d
cqGrIqmB8+W3SMo3W5aC8ZMA5+AUykZlhgSmwRHMZfkRaIai9ht+dtZ9+874ryQwvH1MWnfQcGcA
K66UeTwBvqc1pSD3PGS3NPOHdZhEc8ze4EBhNpf5AU1Q1VPWQhFyoM0TXNcHGav/sWCrD0VdhoQN
4BjNVz2e0dtn/DmQkFd+nFinAMYZaqqWRW/CWUNcUtdvONrvGkF2YYSpoAxTeifpbEWV7OHTdE/m
hhFjTbDHUio4wdshtHsbPniJDo8PZvKgy5Iucdw2eJHi33wlVrRBU6/bUT+2EvMVbJl+gREoZhZz
d1gDU+Xem3dorcYRcgcsWBNOdyEL+n0QBN4PC8WLMZg2aJKcLp0f69wC6xvrrdSWu+AfMO7YAIy5
moBVsp4AX0n9OmRTF1wW6jguLYZBNLcyc87zQ8Ax
`pragma protect end_protected
