// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hWfwmWKh7VZnLpUgpbMKCXnIztBkKsWxSk48z2OL2nDwWUBsarDXweZ23KLe4mKG
dlaJj4BWEdZzpQHeI22Z59WFWp4YlKDQ/ASlKLElRxx82I+KFysTpTSG79A0ptEq
tjuFBX6jd/+5ACL0StclPfhggyVKt7leABbfbtQ/u+8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20416)
t6WvMW+khdpyXvtXPzSFHMuxcR8z8Wq0qlPHfgsqEJ+o5zXtLeDrEC+bR62XhYYX
szpOvw32X6lzXuH+7rmyFMOQJXybzLpBBgeECqg+mHlAqB5AiN4uskfnUuNzPDzy
pEeBnpEHcaBk6jtwKousivcbvrt1kW9MRmyWY/lfirm9QpCKo7hkHw/jtYeglqMu
dm1xL8W5GgzpcRIe6vFne39DJ2o32gIr5YGoO82cg/pQbeqRajLCWVJ6ztJpNNWZ
6OFNJ7MPWpiqOsik711duXfQfYeXktq34vF5QoYgOyJOA90KAUhxSgNnj5XDDVcO
6G8JILPrm7ZlvQX4OoOtPCKiDr/dCiVudJ3y5WD62JHT1t5UfR6lS2g42oloV65J
XjQynOeekY6dgo4y89hKnuBE+J79a/hAjBITBVgmfX8xayJ9FlYryeKG0zmLtcKU
S4eWd3H3zDfdcxgTzBd7EzhSlJ3Vk8qIhF5PK92tpvLc8A5als8QrYIvB5wCI5CM
5vhWk0ZCAuukVSPtPlE6RZZXcaPhcwj4FLpiwytMNPbA9UQ4vGsc1JAtX4TwV5KN
RBJDcsBthxK8315q/zsBscivDFi33SeCW0GuyVswRLPEaxt7P7IvrBXRPUomMQXF
Uuo514/bUAyYdMQJIKx7052EERXKy8s48/Bv69h7XoH9JjeFCv+M6oZXI8IzTCxQ
iHGzki0UR6K+CkfRvwTz/4W2TQZwPulH5p3ARkTMvH5FnlOELL/s8iUC64P1IXrv
h0jY+Cr5RAzf56JxbHipnVydDfT7AqZz4FdUY+5lTzm2hy4oQdVhEa10mRPogM+t
Ca8ZgIWT6trK2Q1L86f2S4SqifYOkZfb+QrIyAX4z2JPUw1ngVAWM9+nP4I8vWFn
Lctsicy1l6dVfNkqsv8cLfhAxRxe8Bdp/5t+npeIMeM9qsUkQgZ88luAmeo+ePCJ
pslPzDhxjgpeXgMcs5h8OshOk/AaM/LU5ejqVWu9T34pp2KGXqTcEtOdrdsfU9Ez
0RmJcJP/QL5BJHB4Aem9JWO09PTIfu8UgKDuvyCM5ic/axbUOyJ+1UyTAVkzWWed
29z1VYnO7iwl77N/rwCsab4U2ec6kaec+Tojcayfn7+WSZFIfNr5HE97YklsAHUT
H9mj6aWs0i3Y6pZn+OVfL0AMoNd/1oAO/mQYMLFCRtosL+r9CSJM0hkSgpi33kAy
gmhqZPIyERH4qZKqA1Se/lhpRv6nAlPlFFcbXSfYwcMIV6Vi+1IhLsZHj9wSu389
C+dCChFblSYHyOTXvm4puu/xd4c2pBbBRTlNPhLS4Mb6KGDU2+12QHEfpARoDR82
Zvk0KqkSNFd78nbTv5ilndAzZBn36tqMOoBEnpwP4KONvNHH6Gl6jYmDmKVQZ6oQ
grgVVApFiWEoYYgO0PPPNuwduaMc9VmYjf345pmsWiEvockjVTlT5nS8tevIAqGO
9SwJWOsaGDTyCxyXMOpPMrOaZ8lxktXRFL4kcpQBlZ+WivuMuYpTMSK+IN13Vl+G
9ezTkPa73dBd1BekOwlHVMGFVyCAm4PxGYa5FI7w2VwV5ScHB55qL8XoCWSvy6ok
X7gUjEZbGWKVM6hAKQ1gVgar/EC3ufQaLOaW4yWbJ+wAfB8p9mL1Du0k7jrnwdYM
DEuFt7u/oSP4TRZ6/5ica7GkM0N0AVAKGQxnZHE3VF5gJdDLKdsoB26xHO/7JOkq
M3MuBZlr00oC4JeR14iZOzQouP6x6GVF0F0V9oiFzCr/eFPGYmHc6rDa+cgkb7Ed
C/lwyq8H/89KzwqEp2GyAONwQHSo+pkA4HMXOBIPiF1+6OTRGSZlEEbWfAtji4IM
/nUv3bWazevPANRTLv73Si9N0gUBk/gBcy2s3aa1ionGLJEBQ89LexSS5+w+mWjq
1n6DdaDRyVPdCNOeTG7Ri2N4IWhHERjeNIlg/mra2P1I60xAS61J3Br+md3yhPT6
4G2S+arPqhy4zndPEhgiXH5yFIA4N9Wp9EiLIud57P+w9qyTs06StBqecMJM4rTw
ZWXeEOiz0XMiDBRb4rHnbou0mXn4+UwBijR8lX6N76QA4CgWllLRUmqTCQuHkFVo
XcNDLKJKJUxlAyg1i7HVw6X423DyWGFT/jnV3OZrmKXpJxeWDI87JmKKye19RiwR
1qcbMM5lloJl2SLD7VOt4kROJdUDV2y0lUpVkPgnAHmvQpHYu2Jb7uaj2bgNQlKh
Pewuu9ujdpHSuUYq/MFSY+2MpKr9eAyorJRLGfEwtUa17MVAIF6AzEUj4bw3LZDU
K8EAvyUy9EdEUDRhqRuZcT629BrwYS8rlqd40a9DXz9HxC1LWtoPu5YJ2P5rn02T
hoamyeCplkig2fKBBN1rQiZjnqkVYCWMPsnzTBkSxHsMAxbpBYZdHwowp9xPMgRm
xVbWry+dscljvdeNadBdX4nCSgtqvQYVgYmk2N+Zgzd0inY57IKem6bs5D+b0UK+
PepzvExW4HoFTiD/XvjhfLLpUb/k0PlzD9PU8TZAQDVlMHS3NCRmoc1Wy2ld6PX+
6HLNlJwNxyicytJza1D82hLwiHjK70Fd8/nCrrdX9NfkQuMQtXyxnHXW4W6JaIZI
meJhhIelNyE0jjMlz7ogP3qehqNq/7u7L/3UrmcPZdMHzapmxdJ0NhtoCd63sKjs
XnzCToDck/AuDu7n/Q9dLwyqLSs06q77+4XJWYNOmYWFa/kPn/xC1eMPslNSyagX
Q0nwx1et94FDa3GdeM5iPqDhW8/1Rsmz6zj/3/hsIQ62+trowP0xG4RyIskrhenv
GH7Ble8JIPboMGTwTF7LuxK/1nMekIm57jlh5VatB3//ov0scblKSVzq+yYq4YFZ
ZO7NRZSYqbjUGtJMNrqApdVLNIpi8L80wvaCl+U0H1QgDq437emnZdmX5bnE72pI
pTbPl4trObpFuaCzp/214AkvgFkCVLFWz5uqSAhozE3SKIIEBGzF9Kg0V3dkNtFo
EYYvlRt8X/2zsUGpg9aY8wHLbgyRc9bSAn7Nvktkxwmrg4SuygIbl17IbsezKOJr
Tp/J+3unyNgv8+w+0dmkaeCHwBpojc4LZaexiSzmCRuzmI87Cdh2/YN5ZPgR/PV8
hN4cOKH23GHYrT0Yxb+twORgJ8deOso8TxV1BlwNAgEczx32HltPycNPp0dnHy7k
EBuTJJrr0d2mha03tg+JIYk3e0Jixsnf3hxZSYJfm3GJhhvGmQ6S969CqNfN1Qs3
kHNooZArLJR4sb0qwqfCG+tissSilU2q9+bXv+lObZZMlvnE1DVxY6FynWIremkB
sOl8SBQ6qkC7aUwuJM21mwW3hpcM16jDKb18U+WkPD2+ZlR0OA3AbiEpxLXDGepr
Dry+blMNjctMYCckUlzF55W1Tr6ytyj5iUhwg+WPDaywRfb2EVROmn+SnavLBGyj
5moJ/eUCv0LVqBdfm8Zm727Bl/0FYd0uWw1bUepO43wS7TnxNcckYQMVpaR9Wu4A
+JkUjC0G6PgreTSh1kalrG2zgW8SzHWUpgyDfd2+Oc+j0Soxqqhk8FcA6o1qWNYq
fnUGJSA4hjNpd84SXXpfjUAUqBJruJgUkq5dAkn/ZttjTfTYI5oFJYXL6cIVyNCO
EJH7cc9/n3Uq2GZtMnGzqORg0IpDLQQgbUJ0dll2W10KIgWX7aNnwgqbD++A+zOF
QVhUrwhZBCMNTL625TV8/pYyrRH/l1oqMNSADxd9tkd3DxR/aEWjqgmChbg6W1Fg
yE0ybij+vaRggl4PkjSBgaRntcMoqtdwrA5CT9zcH/sLCDGmPiP1ZX3xm7rAW0Ul
Kcn+3Js85WtIGICIaHQYWCXwMupMXtVjNlmLtm9A1QLtS0PApbUHx0lz9Gb5+pG2
pVSjedw3wHxEBPO/7FI8yihWI9zBGqYJ11ZZmpVQJ7KWGgTpSqNVt4VOdKyqrn63
sqklNQgPNog0mC9LRVdOm+8f9DbsrJ8KNUWK1MlqIP8bUI7HPR3kEHJCu4kEoyq6
Thd+bdPPhMqi4PoxdjRkbUsVwDSLgO9rPnjPyJbfUlLjESUDXFgOWgaqYKHUicLz
RmJqn0LndCVlPPeIKQVwiH1LSgueE79XivvGSEYhQZjiFrgPbtW8mle1vu+FOK6e
B4Q4ySlK9GhN0mtOnUmmt9IEQRzIExZvmz1K8A4mJxBLFGoYDUXf/aUP8X9rjLws
o06SXOcj1mT/WcXy2Sz+Bryfzcm6ovtfqobZCUtWKlRSOTOljy0bCrEB/a8eLK3A
7yRbyUUTBFXJ21NLEUbBlHmXBTurPBTl8mHCG29h+/49kfTgzfaWPrqmuBwGsDPR
HSC1JjUZpmLFtoL757aoBlP6zi8VSk/H+72+2vWQSfzxtVLyVeSrs6Zh22HjSuYw
oLtd3DjUp4yHNENgt1CMDooNXMz5kOA0KhU0lbZ/D7MQStdaytIjwluECsiSgwKq
RSMB39fCURKoTvm/hhQPhVF1RTLDVDk51kiCwmzJAVUHvmVPTdi8RglnYmVWToR5
/OYxom32hbZlBLB+QXnSdx/vl3pzqF+kQuL0R1zNTJZ25H5+m1RsHx+fAvTZ68o0
AdxwzCaFP1Ybpb9PeM5tZhUaVKUNWoRaOAERE/tsiurGBERpLqAqzh1oZ3+XWjyk
LSkbjjnqSUk3CTOqpiSGjIB8SGuLHMzser1fNwIX7mYSyQzJzNvBS38/eH27j+We
PsOBOHf1Chk4qnti5wR140gWdfqLEyvbkmgG26To+8nZX+53emJafTr7Uo36+R2u
6ieKyaHPx4wmQD50J8l5b8do6ngGZF5JQg4zJ3msBmcIaHS/h4neeJdDceEX1Df2
KxFi3FeGu6No7lViNTiuq1wJltSp+mYBGCzjavSxu6lfXKCPyY2ebMxo45Z0px/g
3qhuU/nUPh9JtGcDBsc11dY7HQj4ReVpsTyFn2VEl81ZlaxfrVIX5KFKdUyixOtf
wRXnHFCgl4P4D1GMfb9/i4Z2m1f/hrJl3n7845xoWpfDLScRdpYDe0Kix81wUIq6
tYSQ57B0flfV4Dh5D4hVAHiE2F12bfybyEjPneFrymJ8iKLdB0lSnurapZhXSt1B
lCjZ4/6wYlca6NB4XlB53yGEZ8EIwmew/SnqkKsgjL6VvrfYBG1zj7Ik2yFk8ZEU
a3J3vORTdjdIwgoVhsOz+1Cn4sCdZQmXUuwxt0oTvB6cWquHHY3PxrJhaiMtvx7T
/Du2zwAxbr3/GsEx9TuFh+NbmFLCHBXkOsAFOze3KUnTGMcqFG0Sb773b02YQtGL
Jt7ImBCwLukRAExteBCkM18nTvRybT0cFduzhc9Ws8RBiTFchWb44Dhr+I3fXUbI
BMX/UxaxXvF4t96c3fcaQUAkQ7wwZPVOtA3FcAOF0E7bBPx7NHwm5WGZAxXWGn2N
koel/wH++DXEJPf9nwWJ/QS5ojtRjm7RMZXslOZM6o8j3OEb3JcI33M7IQc56+i3
717FVwqoYZLvh/q0zSG2nFmTaHHajkpuHVOmVUUN/S9tpsg7cBLCbYFF7DdYg4N7
wUfTDp79JOkGde2ebdv8btr92G00RmzvwpA9FunuHvVZM/TgJ64v0+Ox5cBDs66b
OTTx1sJbNtwMJ8TAchUg5cT9tkyadXFyAA8WApxsIWywLXeaKEH6Y+f1Wedx44kT
zr5cU54ST9Y8NhtWQEOrzekYEIerMpaNB/N3ATuUsb4f0ShTPoUIah3/WbRqzaM5
+sLPBLP19AJiZjHNh8w4ihLijdAJGZwgJFUs2A9lfOSO7xRknof0WeunaEJTmye7
Sr0CZuPBfTyCaFUJKCDUZ1NUdGjalctWtIdUnxhT1V4l96SxGQ3StZqAK6XNtmW5
mpwM5U9YT6S80Q4inLbMX/My9uu86kk828ygGXVg7eetxH3F+0yPH0IuTW9crcYx
vZpVxkZp351K6tUu6LCBJ/HYSvn7LvZ8fhyn2NCvLvgEvptNBASM1vN6JUjmVtYX
WneTPczc88qoeBhCECdiHdvgQ5lqANqzjpCp4QbbMrEvwumdqo8jSOX0XIH6Dlxj
W809elZp6+22sr2U8W03MzhM0TgxuYaIdRCRKkflsPFLnhdrN2Gwv0NU0cdoSRqZ
L5Ev6nepHwJfI78hBZvxjsnBBefNzlfyKHyRtkiZ/bSkS/ps1spKzfEsFpkp7J3J
4rqEhaOygarahZ9dQwahshpzfgX0+75yVdjHmRKBHJHJ0o0cShi1rSX3HUO3r7Lc
U5MVIz0ooh8msVdd4AL1R3FGmbt4lhHkWzvLUjEC/OePrQF9gNSHUEOGVQbVHGNA
dtWIGDHKAfj/lUWm9M6tMolYVHeneQYi7wwCXPkluShzpbZ8fwNibew0Pvpup1qv
6QK711YnaTvXDXPFMvx9HrNEV14kW7fYWwsZ7ReY8zcRlQgSqbFouhu9uXA0QhJC
3qB15msCIAWPJs0LVMrsqYxqCqAqKiwVPH7jRp1i6lk2TFOk8ksU2PTE7kLZgPcj
dKvSyKJopyPtKMC2B0JPGrsOQTFLEBA2jKrHP3BmxtSCaZa0alfGOmFB9sOONLxM
j6WHa5XTS0B6LwGjNAX9XpEF2Kwaq0lAsG5REhpL5pfJAVx0DhY9TFRb/O1jlnH2
/9iBIYSEp8sbs49ifkGQdsPBH0FPmcZaP5b7tzWW1xI9ILR8wSv6X/Qju+D5/d7l
JtqanYkBHbghY7ixuxrFEff5HV+px+4lAb1GMyb1aHqKrtG1z8XPz8xN/2BUvnMO
Mf10yiVBDL+4+r7/xWv5y5Jpnw/hF4RG++ZMDTXxF7kN73CXiCU3owoAZNkm3H1+
xNmfS6wCugfBcwbKkgOcN9Tl5S51X3QqEEqliGlj2G1EkpY/QARwuQnWE3A+7naw
SLUczuzHZQOG7gWjV4Y6bK3hM1SN1Jd4rRWh71G4ZPUOhVzJD0u7XzBCCj57s8FD
1/BFHnIOgq0zDjmQmY4t5ZvFmGKxUiADkO3792e0PgUFCmvdpJWC7bUzwQVJe+im
qMG84IYRQRivt785VLwq9smuY8VfcxWehtXNroeYQDo+x5CEw/FKQ9ztRpKO2SEP
50p7Vnz7+hgnwfho9UOgVrm0VuK4TOAIavO1y9ur5glvU2aRWyztfEkd/FZZ8+Vz
vi8lwTKUTRfYY38QHctGlkQ67YTm4WVopSlx3XrH0NGXscFPXqM9zUPuEASiSx4Z
2gcS6UQ2MaQcKYUwz/EI2cYXr49CYqNJqi33CzUHaY8de8egr1hVuyfUu04WL8Lw
xBxmIwUpbw2gab70kdRRoD/5M2qMSMIgsqV9+m9mHtndHHiFLTgXiDI60adtsL+w
xr08N4EOr9W1WXGGWiZQaYHkZOHV/roj1rQ8g6rfLXJwFO+vjWG5O1H3NpHHN3cl
3vUT40HJ5KMAjCAn7KP3QgK+Ah0XxfLIa1BcnwluQIarckwgtFAoG3HgO9Big1L0
wnK3PlblFYwuQ3bzuEsBUoxG/RM7HXZAr5V7BE7RxnZZbKCCbTOnvz+4UFu40Ek2
rTWLmUdQBfYKnHowYkQTf5CC6FKDlGMIWH+WaqNYOpRcIuFe85dV4RLF5hBWv1fk
2JqTRYE1k8oOjOSU63oNKFf54z+gIoTMmsFXmMABZnvmKMWfZ5E9/l7ljL2Jo+CI
6LDXYzJMw1HPAqMxyWJEcyYwoG9eJVPQMcN8MpigxiV/0ptCTsv/1P7ojcEdQQhy
ZxSKUXCt0+0UddTt+WYe7eipNNLiDN408QMtAYCi6CxRRHIoiMGitZXDG7CYwYU2
qu5TgZZp5nskq9eN//5hC/xWLdA3vcjbg9qA51XaboN91Vqde+P9NPgrL454ppkd
Dt8/nJOXUF80uG+8IVmM9qDCXNgWtVxaws5xiuGpW+vIrQjpTg31l3CP6b/lWFfQ
Hr63c7ZXecw8/+OYVe4uiIN57B5rqnAxqj3uM6u7i+okBZyQ0/YgXKT8az+2X4n7
CecQGpC3H6AQKST6ko3vVOVPoDOi+FZnfgveIzJ/JQbgfMmEuxeL4ZBsk/SzvGYd
lnb2nEPfqa+UKbCexRmmTKY6iQxIbXYKCta9vwPtvP1Igq2VlYl+fehVVf0IE8ER
6mJ/5jEnFdhwFrYP2Y+V4kq/ZxoLIZXdMtiV60eFgtLgKQz/3ROa+oAGCVxHOL1j
8XPVyuQWpSmW0e9P6UhcCMA7MYbzITe3QzDj2Tj5Z91x1OWUxdVU8+zE+bGD7Lfe
2IJmkTa12TtehrBUHEj/nX2f+EKFg2EpWmz/CVtbZTDoVhLv3ccuXPBagcJ4+KkV
ZzSZsbYDxPQ2CC1YKqVTcertLJtFV2Y4E1mztbAJAuUqAiDWZeuVf76WhF6GkRn4
ImJfaQ0iBYfd3T1ykBIWR7qW4oUECVkrY+AHG5duPFH5w4EP9Fw3UwIqzRj2OXd7
grWmM5LUHAX2P29KvarFaLV+5hNil9tnyuAdVOIo07Um9iD/fkaxHllppeeHss05
/zCj1bdY+V/A157sd6AOHe5IeB32wfzOqZ3Yd9NL8vyQ2DgeTyuokyx1OvfKB0pV
EqMiaBVYwRsGyAipKkOV2oMjA5m6D3O8hTD9nO5ePDFqDVYzrTOhhrKSplMr+S1o
tUrCYpsTxcFao1B4cPdxo3vBf3dzY+imjErwMqPj/YYJllAdTAqLz6PJRt65RSyW
/XvoG3wKR1GiVuFcNK7kcOrTAx2GbCjZF++4UyqBeX9FceqnGV3OvUUY1B5PS0Zp
kFiAfr4+v93+/RHN/8bIr2kDswk8SqQyLAL/yJ409Lw6HozuMpzRkpQfheeacLw/
4OvKFiQRSKV/f/gl+5pjUkuD4+ut3WKeQ1kr7FW/ld0CjkmhLEnSDh/3YGYRffMg
SIrUAuYGkZT654S6KJTMPEOiTB7YJuVGgtTqmfbKrmH0R4aHQne6TSomPxGvilzi
TuY8dCF5CkgRIGy4JNWsyRbk9KgOwirYm5tRtfkVKydPSPc5LY3TvQq+42DCEm8N
u3mPWxn9zdNvuUySY6xuNeVHLUPBlxq5FzNunBNHry+bycqM9IlewbpBxe0G27V2
F0CyUm+KYSWB0efyD2XL4cxkGfamd7h5EYnCJBaK7+CFZyUyyqGLEAFhApElbc+Q
xB84kBmMWHKKlmQM98aBy5nVO1FxWrgzyi6V8oQB1bO8QH9bEAamLbVjphKmzkRv
sX3xW/K+gN2/TzQqSQKhc0+fbyisviuMrQfOtXECPtUyj6vsJgJsfstMvXQFqE4D
Kz+1C6E+fYifFHiydi0RC1DB6xvGBxQ4hDJ5NrVBy8QTdxM69zs1pnYS1cOA3hOg
gkxt7R1JFxXIwK1R7q8N0iYOXxqYZclmFCJH3b4Kb8/pInC83qyy6O/74iAOeCV5
2pHBxDRdQ1UCh3DbHJ1txh/5ELG4WWgF2dQYMiZhuwcvfTKYEWFNd46lycC/RyPt
T+IcjMzox0FcX6q+VQsVkS+ZqBB6pDbabzYq8yYwjVnPt0LL/ZWmmJIR26DhDw9Y
Bs0Fodn7Y4+6jS4EIMKWVi+osxmCCRGQbfeWlLLAUBvgId7dJzrQaylly1FXQXU4
X90P9sZUaV9T7JVJvvLYps80VO+a0q7ZwdSzgulG+ErbWjuW5J6AgY+couFgtCqC
CkVBENDzMmgJOHTeQQjGmZ8kgzV9GnkVrOMRlsD9HsrBMWuxBUCXPLl/hXYGu39V
asDudGJjGrCabvRSRMG344UouNk77Xl9q40JuhdEnFlmJLb2QN0mlgFxwYBemQiD
oCnKU/IdorpDNRLBlxmcpRI21+OAgwVZfQGQuv9G1ZgrGX4alUllL4yVXENYCihX
42yy6UyWgtwBTjeR/qkZb5j5QYl8xhN5y0W99x/6t9AIDMSVcab/PNY4kVAgRw02
RFg5mzr2Ft6l4fFMjDyOOOcAULTgRwt0d1RICmmZkNsx6T6/0MevxCYUAhaeYAmd
N3A65hVdLKAPxohzq6COoxNN/j/8pK72Dz9l+vMiFgdSof0cqaGUMD2dgQ6c6P1F
83HLOaWD82RNt6uaFExeUEdg+ulTcVtoujzccoPmNa1NBvR80K+S0ZCFKGbHmBqp
nVvr4dbeExUSXuaY89kM4QrwPzvb2Sk50HE0JavFXeRPGIQzaVsf+sV5t9gXXPqy
DH8yT4CBtRKBcCBLmbjBYttPQt2m0afSEMirO1bf1rtfmrSs3Ly46dd7lKexJJd2
6vej5xX1bex6Pg596VrtNBfTLZrb2TQZnXi85QOY25VpaA+5/H06PHabx44Q+Emt
xZScmbNBN4HemzGt7yudCsB3A7EECmB2t81YOZt9ek/ibPW5QQR6qYt1e9gSfoOW
493kPaaWHI4Kc9AIlYrxfCp4jDm0V9jDNq6iA0TM1z2SCQWyr9WTAqF5xAnFzuJT
XkIO+Lw8JYNvcZVaLT2En/5wBjpI3b6hmvdZADQDnF57Q+oku4ix8WyHqnnDSHgk
khogTzrXQtlUMptZN23tBAjiQrgR+WZmrxp8bu4dcY8qOeXV/LlRUR8oo/3LhZhk
KSbvc7ozYnb34cbe2R9RbS0cD957SxhpN+U8k7g1L3MSfVf7yIkDlYplhPSN9h/8
CGWosIB52FxD/TMPpT4rSMpuyGeKGq39/ve31FMjHQUPzEByQM/ylleWNoGoWg0h
ZctJo1+GORhL5AJAfCh+zTzX7EBDJt0l1rAUUCFqBDz87yRpL81eU6tf29HaSHzX
XLZvSzHD6lxQjw7CN4HH9cY3yLDqmnxOPICx21FXmtpwo+59vhO2PqlpuqAbMBd/
B/I/mABy0BHtXr9oOrPPiXxoXGHNEcmdOqzDV2Gjll07clzgo8zwg/iwHx/AenYH
mZ5nElXg5JUKnhYycMzuw74jIfOSDskwK3szb2JCArmhkGcikjTvm9L40lxs/6fe
LR/JeAP5t3i2JSVF+OI+icZodjBL3v6s6RSvKRBNBWl/LVU+5yxj/P8oaVefAKaN
66ma0UL1Hw5exEOR1tF8G9ET0NoLT5Gmsgm4LIZBqrQNAmf9AnalJX6+wzc1pmrg
0uxMeFjg1vueTvQVPu+WwhWaBo9qoILHn8miziNLRXAv6i1T/PJG3p/OyaMi27Wu
bCFAgScETJoUjOaDXD2nG30s1c2X6vvPQaYA/SITyuMEG0xNEUh1dHivJf3x/8wH
jQhQ9BIvAUZ8m6MSF116rvg1skp2I00E1yTTO6Q/ViMJVeZ1pjt4foyaGGUvkKg6
OLHCo8HmMFYMFcqIemjOxP/xK0vJrfSSmDwf63LHbEe6JxriV7RNMD9I6sUGCb1D
kU0RTAf/SCu1QQta8S6/gvz009URAbkz1Ip+oIRgq1md9xcH4qvz82jGdjOZCmuI
xBQTPZXof0aLH7r2JF7ngoYM2awS/5EgEyDgvjTr2uP+0tHIk3gpAa+TPtHA0mYY
fg6QnIVbMHn/qwZntkbTtLtAXUrrdpoZ9lFhoGDKfnKZHu+Oc6diMZzL+uITQBs3
+a9drNXkE8ZtAL3+ezHgkOIDZrxEYAXFVMfkuqhw8se3xCHC04kjQGPHvketGWai
TbP6ELtIAAveackXdaTV5+CWS7bBob/XLYRWXhqjLV19vN8A3N6UUw1XR5lJYFlR
43u5pyUzC+dBtdqCUT2AN/5cXNtuRl/kWpV1RJ0fF21wrvkytGdH0WnejYiaiwU8
vFUl6l+TvXGU/BLQiXiBZ2s7ILauVJnF/ycHGcXIS6+eirX26+lv4unyGk8k+dlS
MlNPJjzj5mQUaeBGBd+Q9RiL26uiwO1uvIGtA8UGZ0lDw6G2ulM4+bJL+UGV1SoO
2NSGxpUEOl+DeOcuMe5JmjFNkWtxhpiMaKApPwnBlQnTgk8pT9r9GinsPfJo1ztq
9IVsiq4dNrIS8Ctz80tfpuroOYywJfk8D+dB+TNjb3PIU9Vc+HLUMzbuww28Np9/
Icz2GRUdDrhvkPsSzmj/HM6khHWfm3KEe11rCKaUhSlTN8MI5fbig3rOya402TZT
Hu8myMSNc4PkJ4WCtf/Kh+PV8YKDko7RQJf7uIZh5CJf4U/vduEqSbiqfKfsSOUd
9JNeFIeUazroR1nTVghEvhqdmvWiV8Yg+6E1uUNiyAnjAkW5/02v+rbuhItAg/Oo
qO4ctL0i/rEHBVx/+6Fn8sxn8s9iEgQXXd8v2CrBY8mq/DHolWR44WQHZm6DJLMw
sj3iX1lPryjuBU2f0ZAPr9Vly6T3+LPHRviUNCi6Pcqo8jJCsU2P/r1IEt/xiWfa
Ca6unkS0d+3WRj1ckYmIbzuYqWm4sDp/Pd1sYtVo/GefDrT1/D4FM6QWyhPFFdG+
mEEA47yJ35Bm6CtfydVZ4nYf1sk/48t5qsbqDVFhk3Rz+A+weUW0O7av5kZAmPWI
TNNQ6rDuarmU0OHGwYUHh/pg7Q1pKbECosZcV1yDJwExuVOvGRk+1kl36rWA3JHs
hesyzCZltk28AmS3NS7tNEu+s3MQqOMSiS6mLRyt3rxpe7XcspGpoIa9gCXKDOJm
Dy1kFp+Ixqu5pVb/x3HDBwt4y1W1PtLe6cExoMrl0mHjyqG0wKDw8mjg6x3AHKoT
ilHZ9O3x6n45gFlnfXh+kkYVkF2kaBauf5PkqCoW6tMVrBNjnCjPgKTVem4SSfZH
vmZdLwG7nPTeQ5OdRL97Yx2Ge002h8bg5/U4b8vcLjzfrfnMJa5LESKDkDuBo3zm
T+slWDqaQBe2jlQ1dxPl25vkP+Oek1K9M4ixQuzcm5pFdDmbxQQpCP5XYv7OWNXF
oqUV7AGjU2lPDkWn22LXURvHdLj7ofeeTjOFn9UMSUGuOAZVH7FDL2cGCA94NmzW
NvKGqyNstHBXzrAgjF2VZuqqp0i6ncUTUsPunvaytl3kP00OdWWZQ9vi5m3PcLDM
7pn+uQJEYKGf8EJDjkAH2g/1VhAaiwZ0S1eM8lAqu+JcvYf84528Tzw/WBO351pq
BQUDYHBSdcLXrZGil5iM0SJXKz2LL1mdD/6Ui9lbYdpsxoXNG8XkMvzHEv/6z/Md
8KhPZENDcJsPy9t02Oj/vFXg/Q/bXLwsRhfsq4cLFi7W49e5jjfUHpzbhpP82CZ3
Mo3QFW5dfHtc2mr85xBesMqHtuQ4gvfTKo8P6u8zWLhnOgEJoG7iqJZDfV0s2cVc
tbJK23dlipsKfOdNDEddTn3illfQnIVrYS9cLqsXSMPFqAlhgTkRX0a+gqcqfTpQ
Ty9qb58+yAdMb/hTEaaZPZMvUIy7racr1/qKmZkio6CIQz/IKWfNjzFlgxLV1JOM
x3x9Z+GcGIe4ddpvlTsyTUbNknfdLAVOAJJ3X2zIcHDspLA/9D0R7dclkgBm/ysZ
2V3U07zuW5kkuruh6mLzdymVkHJJzT5wAOGMC+BednqYFh5Qrd1iTQJkSHV9eD6W
XSb+IUFsLsE9hI6CNH0F37l2utEVJs7MoxxxtXtSn8EBPhA8alf5tDidMaJ//Q8U
y95/TpRQhBoySa0Zh79iTXpjwyOMW6z7tS9bRr45vlV8A6Ow+QVYHHTnQsAULsAh
rrsiOGo/4hRzA6WEAvor+yeUDoNZYHjuLWjGSrMVVfghKhacp7NiBu8wwukYRJlD
C/Wx0q/Qtu6EqmaaFjpvPiRPDr20NOwmRsL1H9TIVerZrZMuFzBNypbHxZfUWXM1
cEZ1qASfdSsKCMJhqnHI51Eee0TVzJTQqhj84NtM+zQt4t1uu40J/TLh0hcSe66M
o7CZXBmwOgctlzVMXKd4nTFCputt+V1mPwvojAUHT6AItUHxbr3vN5IORn6sjrwY
6c2+portnoyUdTisbvnxgPwYTXikzV20YcVWnOXJZ4bjiMSI+7DbwABZxFgWf0z/
yd7os6O33Ofp76xW1B3LM2Det7xiepW76TpYMsAzfXntaTBJmJV7POxgFbSuLTcS
XKO789nJKFkEFzWSmlW8QZYTIYxnXP9dSsPtDOHNs9eL+xIcY7KMijdY3Qemn8vQ
qWX2SSqYn3NDfrkl7Rw/JqOsqhHDz+j5GZXv94fY0LuUjUyaEjqLieCb4qwy96dm
scsLA6cFL39UsEPEq2jkcbZZ2CV4zFA7D0z/uWZO4XXthsDic66UMcHZdnhi+CrN
9B2qTspKcd9+ughvpBsG+p+cemZlINO8LWDjqKEKiVF+Wi2p8seEf2tQbE+gvbNo
wDM+rgnWqvbO5DU/BSbA837lUpwIzLp4B5y2f9gkrg2M84g3vPQ4tMeB9izVAIha
LnGgXFEiDkk4fL3xILFSJxAcg7pT5NPHhVdYOIKW5RtbVWuUOsrlpPp5IM9Aibmf
W9k0q4mUMSHSzTfmX+eayDQkuaxAogHwwO5L3IRSErAOaiL0rp4AT6eLkGAy9FVe
S+fr6p7hF4L+UHUQ9Gd/VZUgx2DsI2Apw5YdtONw6hYbjY8VhJ/PRb4FG2YiPxeS
Z4C6IDe7GFTSUzHSIhzfUTghpl3mGDe1rF2vplQ3jCT6PDl0ZpMv97LJPMXLitLb
2If/ZEVT/ObwwWySnQ53lbl9OW7Rp620w/L9KN09K08wiuwpGrFFL2HFULi8B+wH
ojLj5UhdvLN75vHtJTQzCTYq6C1A5Fppt9g8u1zC21a7aakwFD9U9iRq+bhc06f9
1MBqnSnOwqJzQNf4MPUtGPZQDuuiBMquHvl/SEB6TNp3LDTbXBgIbuorwXwuSFJK
bBwQl5l/kTQGk7lcF5eZpUBHnHjzbRdtBleQccF2/MpQp9knDQURJtcvmTbpyRJP
l3WYFQXgBSsPPgbFfBVVj5kWERHmNhEuHA/G/22ayfQDeW+7AyD9I0FEyu/uK4pm
PbKwGfdDMDW1DFGZEjJwDIIT/+x5HiqggprVMAmzD9zg4M7WsSQaYNN8zt10huR6
WVdSt0xo8L1M6y//8zvTqBbelyXr5VKbXh25xMEH9TdBwKh50mvdgDnRIjMLCpj6
pSZMMFG/pLp68g7VB6UakLe2HJhMxbFabSGbRY5zYFobWiF9NYoU0vBUJIL/90PQ
q3VQsQQeQDZ6a6jS0v+0G7bwRVO95N2cFNz6IENQoXx6JLF4XoG38ZWJXX0nL80D
VPSiWMK87To9p56/mGsSSZDXKm4hMnvzeUvFpnoJgYyIUdhmiWcAJkr6jDZWxVyj
N4rwd7TdiYImeoF5cY49R3D1L++G7RX4SN698LLIMfI3xSC/Jg3sWCqDAffmWPE0
eTGq2bEUhn5VHD8w3NovKcPe/ftpu1r+zDU1u+zgmCEE9Arcuamh3cdzJ+nhfvNK
zaSN/IOwSFAkOYH7/Qi39c9bRuzoA9xws9qxBbnQLPTLEjeFTxEqrpJylQNhoJOo
ZkrJ8bQNS00rKcSkbFKvAL3yBGSKAbGOWNShcCNO1QasMA9Sk/KF618Pcwef9v8B
Xwa3iYC0QDITdrmD4b6r2uD9iXsLIyoOszmmEkrWGlRvYV7z3d2XtbgmvFmG6sJw
srgDQKcEmfO/peIh7QUsMEB8WC/eWMsqfNP7/BcFJuM2kIfTQFS/lJVJbXSthm4k
vj5187c+xWhZUjLsqmh4ngy/KoslRDFebumdYv/SMWU3DheCZIRVVGaQsVKPFHYV
E5a3cRke+vCKgo9XsZeUcxUC07JhMT8MMdCSWbmHHJ69qqfpw1DDq8k3l1Zc+1pB
a5FO8/mK/QR8DBrfTAedrzh5OkELrp9v4GxVV2kseWD0zdBWdNv7dQh2qctXXNyb
iG++Vl1vLK6yZUA7f7Dd7Gs5JGVPZUAp62pNKTrvYTZtEKj6Mb63pvQHkF8JiRow
SUBVWZWFKn9v69ToTifUSJPGjuRm+7VLfOMnn4scsYM1M5dgfmUW5tT1fNq/n6td
LqnDXPDhdt5Y7mRED4sP1nggvsH6WeVKBVappizbdxag70bqXjtbmlATDfBhZSLf
oG23unAUvgX9FtS/362pdSLTZnHNsawtjJquLVtfJOJo8YZVCTMTX4Tf9y6mrreH
1jgtokw7U8Cx6V/h7ieDrQ94joMGywzjZ0gNDwkY8pniWUIAtTiP0CzBPYB/pRKN
3YGoIHRcsJ87p/DBlNOmmBqDe4opDuhknLXfmR3mDkxBH5NrwKr/rdMsytTxHMHB
55n3CHCxp9Eee0sd0fCleGf8+UwTzhilFLgtiiXIC1MFROjZi6B0CkF9yOYbi+AX
UiEv87pHPDGGYaYZp4iTUfXmJIe1WNV48OZ5tOMxx8PxGF7VKp9JYIo5bSJtXOHe
fNcbscf8aVmco1PlCU9Fd2VOQ5w+OeC2FB50E/eTYQqMjRP3jn9+vSoGfksiijcY
H7sWpXYQucq4bkjaqm6WQ+D4BX1+lpi9ZrL8X+mVSdwlNGL44d47vcy/ekHjQMVH
O4kXy5Qm//GRKXlF0WUyBp55lW0S74eidO1df/on4dddfmtxSKb97bKIEjEQOYqQ
4x+yWArec1Pi4Ej+V8gLnTaJ+FiPFvwQh7KdMvS35xSF3AB1IjfEeRVrOl8xDFQp
mArnPzSv2WCLBB0xtImP9JWoOptNyYwsz2Vo8gHU0zx/C8rpgyxgoCbnRy4/liPi
q0nfwSjrIMKSDKvRAXdzIXjeutWPKrJg/v66bBkbZPUovaKDOh2K12zJOdi36WOF
fjEwl9cklFyt/2ZP2quPqzgmYtHuJLJSCWJTwqJ7tRSTA97PeoIqLDSVQtwffSWI
5R4XUv4EfewhhqGsXxG9oZby6dUn/LqXbCdfi6hPLYXsQSm8GUApOkkwxKr3yrQG
ki5mJLCuZo3Lkhwfj/OvJFnGGw6fZGdJvrukyr/vEOjRoX6PvaMOQRUYjkkC3mqe
JIA3Cuq4thYkchmvkcTbxctK9JhaOjABinttXMkl/jAN6gbHlRsg9WJV51FrmNhX
EHMkKMVKAwckUf/RcMCh+wziYji1SQjuREiecCWWx0C1HkaKSDG2ULaBj/CN8/Ji
xiz3qcSlbY7O+yNai9kth05i7nw0dYe29QCKSFgDjyadSfInmdH8q24SJ7murlpN
UqGzj9iSdzxU3Se0JVWqXrxJoJlPUSo7r9o6V9FDA6rcWtBhS5hecfOXGm/stxq0
BgL7A5BMyLK4HEO0e2uXkvWBiW6TtmGaCd/LSUT6DXTCvfr0WbqmeUPuULXEfKV8
8YV8oI4wCuhagXjgKwLiUuQxLnEg1MrsvViAsFk6ceIiYbVkhF50OHEXDt9Q15mc
zjSXcKciLYhzZeGGzPq779uAqEmGDUEFrTglnBGdvkpb9ySfLGaRb+gXdMka231z
hRjKDrUUuyzsO0OQ5tB+U3iTlfDMJ+puaVOfV6QLob5prEKuOYVwqEj60XK8t5Wq
QaioWRQbpsP2EB/YqfEtY6/2CNP3F/n+AE+BmtLoIhv+scpmEIy/WCRZQdmJ84V9
s5L1wilR+Gc4Y3hC+b9EPPaBoMG56A3yaadUkA6U7kEDpTrl1NJwInv50qIJtTVE
K4D57wLlTeR2B84+LBnB+Wz9X9/ougsiMAI4wpJ34ShR9fLVguiSinROyJDsYmpU
N45DGCNjxbAmmKoB7Cyjiq7600g+vLbE6x/Mv5RwTIN/tyWi5Zp4nqgFCshCK+r5
+igauM3IvsbAH7dZ/axd8m0GofmDau2T4RnGPCD4M6FN+cyR3pDtMupgrbd0JdBK
Yr2uRKFuIGWJW0ccojUhB2NSTSndKC6NbYwtMs2Rilsmsva/2OofMTS2XGigXttp
P0yoysIpvU+p/SAr/uwynceChm/eDKV4T/joOpOP2JEhoXWkam0Q9V+kK9Xdsjxk
NxWyEa28JSw2SAhzujX5Z8NHboHK/mnoXeiWx21PCTh+m9ShxV0Q4wbKWZmc35iU
jIZ0wx7ecqhNwGSQium+F+clfjJOfPrU3Ta1JMWxZmI899vYsbEuJmuuJyq0KcHV
gVHxkDHGF8WTvJd/20xPNq1FaVcq4XTSdEjp40dLr79uLwhZp3FxH0jRaSNMopYg
4SliovT3wRXIO3ffAB/L95pRJKatd8BpE4w5iGbEgWgg/3prmzAl4IccFVJ1qxvP
dCz/arXM4bM+ipxQ04nchrohepf+O/BA9YWKvzVn3lEOV4gVqsPpAYqAcTy3u+DW
IG/tdhDGrimmOtwZp6CH3VZWQRqnr6lh1ARO4xeh54Zo+DPHi+l+Gjf1slSm42a0
l9XAc7YHVDYPeTWe38cBp9JLfgpV+s82ZyhdFmjCiXMjgrcBGCv2PvRDSpTyPUB/
KAVINbnBTi/uLeSwr0wmYISqZ4fcQCquK4X7Y1DuEqyE9zgj6joIXKCh6/iAqYTi
qFjkTluyglf6wngxipf2HdPRkQcNMaRNet5Ar2cZqsxtj/F/7GXr+xM1WSWuYkYR
o6DAZ/IDU0mREXkxORa1f58IfCnhoPOx7zZPCWHqr8gwOKlF4DjUnnGkTqtJPM5D
Q2iPM+amZE040G6TlrdIhqi/e06vxOxQZC1Ggt97DBVSLGdwEyWL6/vjz54ZFJG6
tt0X8fBWgczf3Bhoc4+I3dvvutbwtVl2s+xvkd5iW6Zsuzew7WxQNV53es+2GMP5
Dk8MNciwxkK4nfgkqBtG/eAcu070sZJjpHZ+JZxYiBKlQAavcPgZvsBvB6HvxTM6
2zgxvUM7rX/Mc/FhsulkC9IzLc8Z4yFaofj7LCxGl/K7BTiZdfPE8HTQV4WCTr7T
dnRnqel+ptJxw2t6tJa9SLHLNSwXpR+l9e+fSb1bL9QaDq0dcDkTR7QTx6l2vgSv
aC9rjRyEJafhfZjlOXc113SACD8y/RcYT2k9zJabHc/hM8EkXbrcDuNLQAWBVoyG
9KAoiOh9w7wXeelKnBX5BJwRMqEkPlS9tbWOcBwd1eUPGmVLKPeMCM622JZb9awX
giOmly+aL48boKezMgad736BjgBym36rgTbXGBrTEn10jHiCLQG3/YFTP7gNtI1n
Wpc8jqLoBMIUKVIrTDCU6IOZ0l6+atLJPOrFyfUuduEY4UeRMHFwuFOR940cdu+B
BztWFi3H8xA7g7BNymHaKphlxSIcFHzGLWYLcJB17HLtAYGcNq5ZXLOKTCgW2OgI
hVdRIVZcXL9wgLcx856gFWhs8uarkb6lwKsgnhpvXZ1gR/M4ucvJpmEnm4hLgs4P
aKpLwhJANTI9JhaxrHmIC+GQLXvtdu2aWKMPX1DyUEoNx+Yve97RoOpu3NCMFrhq
mNgpBmz2tKSw24dLNLQWf1EysYOOSpCqxfr6N5MENs+tqrE3FcI8NxjgTv+3yPjF
9sGxqz6W18ZoGMpB0syZ7GD0XL3lc4KgO3mFrfLN25zYb2dUpnhLUqJpDIkADTLh
XHDW1CfhfOGgbf8Wn3ol0ftFZJ3r8+MaWDM67VHC6iddDCXv3F/0q3ow1U6EDyR7
d7ct+MXCzz/oq9/J/9zaXqDqbEu7zZtprZXfj85sg9aPmnTgUMn4ESB6SQVP49YQ
Ndy5BrqZbHzjt9KXrsFhvL7/A9LfXxJzlmZMsD77UtBEFp2ky6/y6so1e+7tTbH8
HiADAM4yBwPqNGJ6XF9vlRfoBy+hnjBsstci9R6z7NMHaXc6a0OJCnINkooX4ZUb
yze3ZGqz1krWHG/o9jLXJ0AgBBV9FNUg26vWADlKPc7hoVLtE5DouqepOhKTTFIO
QrC0rDOVUhCt7QK/9m/aalM8Jnq4EQcQcJhFaIri6efw92Xupw4RPHMibcaaS7au
iMX72oeC2H0huSgbdB7eMKc4er6mudakfs4CaKU043hr5nMaPhHLvlvs05NVlxQq
AA5Eg1ujf/X1KmrCOYEdlrNuGCrSd8ltYbEMZeqYyHpNB10TOC2gBcnRVqkz2t6o
bbyOXvpicbM30h2inQIeLCIVjLz3Y/8TJOe+5g5FNe9bztR3yahvypPJ9Tt8zIg2
BMIAaD5PyOqUJ9qU8jgcmpq/NpU2D8lMPUQMjDFt3eZJJibetzxWq4sZCdYkyuAd
7Q0jeRHxtQXX66DW/c9eqJIUUU7BJgJRe5yKIdnWpcMK97aoAPK0sGcsSXy0YfHf
P5QFMlw/4c3PW3ItG5PlGDtemE+VKGuFd6dHG8AbCCe30+riPy9sk6JwMRt5ztEi
oi0U39yX5cG1hFY6nKbui2s8zsCyoPZQHPXwJX49X9oq122mEFbS3L8ikSWzvwHv
iaQ7hnDYpllCth6rTKAzybW3c0/FjbMYjF36OJ222UN6zJfy2Tafa3Dpav1RqXOG
UYGKPvI37kxcCtKGNPGygtfOJx0lNjxg/sEcQ6/PfSjvK1uxa42OIczcjVm6MVkL
paZ1C30LH8OjeloUGd5fXZbXuKQKQyLvkjRZxDrdteeGJyrb8qNTRxzex+mplNF/
/oK0WEL4nj/ETeLEVvilkto0CKPbID7xPeEvtPp0va2RzBLjqUgbwMxX5yqO1bin
XvT3YxBhBhVTmRM9z/N3SiLK+Z/4EczIOuPfD7Ldpi/m/8CG/Ig85RKTBV/03b0d
UUJxgzLoykiQi+ncoIMD4Ja7PV2MPpVn3Kkt0fy1TlKiwsMcsxqUp1vbtXbk4b0l
ai2orcPbxdGB4Q0SjM0/eQMQdz1oF6rYP2Khm4WFX7n1sZ6AwJ+/EihwwIpEGacO
aoKTeTeZu2odialNCuSOxcJiluUZp5Cpb0JBO8aUFw7a/NfhpmRSQGzb6ud0mtEz
+puQSQVkULukLgn3GE//biSq/m6Drhtrl92+vXOMrZHgybxy1WM7XsRWEDsrObEs
z0ocbOefdt+JRusG+03PD1uiWjC/dzzkPFfbED7rLObug5bzrITb2sl9hsAoRsui
S4JbvoGUMY3YMtvqaumn5ZA+1JZWdpcQfn1K5VFNtZbUBFFaReoHydvJCoFXj9Km
/bH59DJSIopwNnDKK7yjk0MeD49tCRPrWzLkRwSkmrX9qbmgUuTj9m5gPsMsfXlX
zvBYdvFLSu8gcjIOrbZ3Vk9tN5yUkRAKt3qtBEUh5xF29Haz0Q0Aez50GoWPmGTS
ft/sEib69E0UY9fBEhryHlSNPuajTFUX6O6MJqsC/Nv+P4VpKQHz1vgF8cqBoI1R
Yjp/gK94fWQDHYBpgkWzZto+ga/xsYeZKFn785wyp3lvf6WH1HnO7fiy7vswyuX6
2RmnROjkLNy/KlfUa/9Y5cuPG3QEJRxFeVRs/1OIEHdgFQ966lgLoP8jy9tB6IMH
ckvAQDRrp+ESwLGYZQala6Sq1bCByMmkdk9Av0ZZksz5fzXURsS7Jyly0uridZEV
85XqKjMUJpxtq3A8mcnBeqc/P6jxnPAwCFEee9vqxmOz05VIQgLdIjNts9VFM/j6
DSrdZ8hJsYkEG2Bc5emIJG3q5MCMk40Lc9UoRV0eeeqTYACbr+IiZMNRd6JSUQ/B
/cfEaVqnU+tpG/8UTdY0qkCQ1GdtqQQbtvXcl0qxuN45q5A06sG4Qatqro938N3t
sMNs8949brufmZlNnY1R2+4ysHuv5QTvSFlueGEPfZJIWuRyIbqCuRQH9vAZQrZ7
LaKkMw5fepRIiJthBXmQXVFdnBQpUl7e+4VvUMZwaakso03usC1ou+PkD7mi6Trp
87/DwPOuCbWGVy9WL1qPby/WQZxMuHna5Vl/2UdxxXJssFUweeYEjc9AGc0Ojd+w
O36/6w99TQvM0/oTQKZSxFNEpNCfF6/vX7SWYIPbCwn97M0hv+hlRvVb9V/tjE6p
QnTG8YX7HNMYZK2sY4cvh9UKDFdd6Dwc3B+hVnXlQDU7OO6v8vLPEayPqCeo6HNK
XGCYnN8LI8MoltrJMsIbLMXlil1h6wn1kU6ybeQeBkIZoCU3IStamjMSzocI0h1t
NkJnzU5stcVkktdIpBYbzwuGotfx6oOqonh8GtLt+j3G17PWAuSiNBU36yk8bvgB
XFopXgLOMrR+L5CjFxRyv/uqqWS3aElmRlKXeNOZmnhZeV8oaX3CEUwley1DEr3s
WAcqHgo9CelAybZjIPRApSO5/lI/HsTnmvpoFFFjR+nAlJNZhHaZbVhGaaTX7S8e
1glvv2Sh7/E7WHdmGwuRaFjsdxeOx98cyfVgGwAjyYzT9xeXwW7nKm0pbyx8XoZ0
bFkJSA0sp0tQCBwW/+QB581SQ1pik6E0TyQq1SBBMds9rMDSdkpOSYIlezm0ILMp
Q/jEfD+3H9WNUmbNsqF+QvvLPBmu76BNy11WFbQ8ZsReMwngSH0835ZD9FVsYp6q
p3RrsB4tWkfSZxkpoTkDMoogxp6QFi9BPBt95kIQZCcOWZadpTH/IhdqupzeU+3o
jS130FUY8dSibwFYJyuJgJvYzluAqtr58mWVXNfHjuCDsV5BdNQs9tmoK4MoWFZi
ldD16aQJsYIeWI3X1O76tMq5fs2o41iECOghLCSgktulex/SJsbBUYsg05IPcHkL
+i7XpvNPdNwcXEcY9iqEg3o1UDyY/R9yO5FWD1Kw5H9Vrl6ap1u0Z/MV5r9cysy5
iBf3Ckrh29draPgwDXGXctc3W65y+IZ6aKkPeF9ja/mYixp+ojaVQooqxmjO+mNZ
l3DcHReyuhW6m4bQ8g8+9ZUnk62rG7n+dvsu/xeRrzSVG9x2mfgOSXVJ7fv6ChcU
k0aNtS2i+YDww3tzqbxSuvxo+sBQKsSIcxe65efXkok05AVaK//WJTDMQd5F7hMj
tPysHU78qryW9KvaTll8VKm3lCgN5kuAutIl6f5wwv+fI0waN8NpxL5rq+PxE56x
/9HJikvHlbLu/UaTSu4KNZ2t8puzSVsE3BNlvdhWX2X6GZzr4WQkzj1+0mhzVd9T
O1KKgh+Ea2ZwkGKrrN4UXJAo5FIOC1Q3cMWDKCzEE2ZjP8lossfw5hXFf1vSR9Ts
Qo5PnLYMjZNuXcnW3F3KD4Db8zX/lfLw7TxWbkbat/QVEhxRgMMsN9sal/gForoq
IL5oo2phmRKOyr2uBAK81Q2EeV6PUuwmVtFE5tPYY/yGb2anxbju+fEu9BiSyqYG
7cMn8px2smEHMiqYAQYciwA3HJwa5GtLz2+I9PLy18PUJ4/MOdAz2m5qWzkzBHK2
7o+ACdsmG2C1tHRx2iX5cfkzpjn+l08L1Yzk6lQx1xz3AKEhDsaYc4EZK+G3WWJH
0dLn4XxIuDlCcVX/6FJllhim8K/VVd1zaxodOm38CPSYZpdA/Eb42zkBnrRIUpAh
1jEi1yXIGEOp5VZtARwXw6l88qxwZn2wSJLB9njW86dCuL4PKZxBAPFb+6yaWXgS
t4fLbUtCDTOfZnRPvwPy/Kiuw8KgdPvakPIl/zt6TYKzbFPrCa9JamkU9nsVqHPQ
4uEwHO7qwzMxyDIwOmtn4CVpvJaq+DPnMECfeFTr+LCmqHYCDf9Zyv5pN87znGeP
0jKMfVMLF+23pSCK/zjJkjXvpwna0UwSgOCmfBJ2dWXhR3nYU1iObYqGsRi0+xuC
zwcRC2juy/u1Tccgix+dufN4ylpAAa2bz/yTDLAio/AEEJWA0FYoMAwcVp7se3ZA
ZvjViTLkGNAMa37OnbbtjA/JjcZGZzWC+KUUv7Wba2nBIZVmTmp4N0NyVifkoQq4
+udDn+Gy0xKxpNTBOrbnYvogV6Sc83pWX/XvJI/AouDMmvvSK6ikcFCUMJLkSplH
nbxVoAY7YUWCETIwLqA59l2eU++YUWHJ6btSARQwA9Uuj5Qd6Pme9vmgqOX36/ZD
2OzsWJfO8rG2OtpLQYsUW45n/YEVMJh/bv0691NavVqFIJFInthZZwJiQgKGLr0k
jKT85BVva1zBkKqA7EWtIcg1NNwlnHoL+B4CBqBakltVw4zXP2CwQsKmb0oR0z3z
upH3z51r+oKT4EipciqIaXDbZbRsTvnW8ream7jHI8ta0rszra9APx6KtTN2VUDh
v//mlrDOkOaf3J3r/JsQBJ1jtnLB8pnGzU2wEO2f0k2eBp4c2RpUqB4dbHC8bIr9
ga/K9ipgf5omotjoy26U/cM3xjmlGPJOPtudlpvrGmpCZ+sJvlgGnDDuWlNkZrvX
pE516A0/LwuPNlMe7dhfpbXgiFzcR72WhkgOw54MBweJHsJ9U72YncdyRE/atqdt
uf4XvnHRfZaKLOOzR0bo+aRMTYFfy1fGBwE4pFowwxEXS1QgWg/6IFppJBXwTkgN
usLThe58OEd6fzYlsjmC+lgowKK7/GtgmGkhyWKWRAx6gku4Wjgt0b4a5kY3deyK
zwlG24Jrx+tf0hC6hhUJoEweKd2YxAG08PbdpRhib6kXgt8m6XbrNIHNiVLMbl3/
rzF2lG2pnbMWEHZaGY1xuPUt0UEoGc8g0MB0yeBgMK25wQ1sxFiSQz/uHjyd3FMI
MFaBe3wIFwXKeSwRpT1ZAXCxAiXMVI9qFZ65c+zuG/qKzEgkGW73wdj1FOMpdSCw
a2ncMxp9dx2QV2pJMAQA8iQ/Ou7GdBL/HCff+YeYT2q/RYxc85EEBkdW5bRlNcJd
nP3Ffz16+V9ufXdD7uLuicfMb0I0nE4xwawwfbhgktl3RINKFxPHJMxgdDhV+3aw
RctmvLNDXdSEmFMrIpeltjqrHg5yC9ZnfjyL9xV9D2HCfcId3cPeY0R5HFtH5o+h
x3ze06KLJ0WiaAPrysV6dC63zdq73CIOhRqkNHBap272fujFTtfVf3HX1kkrO5bg
rZi1Q/ebM9V3nb19970eGjtQoC3K+yYuTH4LcFKC5P3djXqOE/AAVpwz7/FG64IF
vPQTyw/n65tNMWzH6crFg9f2F7hXOZofqVEuYQ7epKJjEhytWZd0RhzFJbB2nDlk
aLywSeIf0L8s7zFCNg9xcPr4eo74uIigQlpYeSceAfBM6lYbncMRAKqWr0yk6ixq
JtXKbdMQPz0ghkcqeznkr5RdliU1o6BGwEjqLUqIsIbi1O4JQ9LPkTpFL7z7I3L2
Jq9O79k4BG1c5MxEAO+Kwoy+M8CyB5vmPgAfUOcYoRJ59AyVrRi5TYpzfIkuDs6q
R/w4b6DaQPJxcF86HqoliH6IzGzzYTfARRd9b2hVo8CaHSaQbtFHWtHzJw6bTwG4
z8xglAAI/pTnL0OTqV0RrVmatprf79RR0/plmO041kts7kl6Kjl04Ks9q/uzK8V/
IAg3hbw3Z6f/TwuqmtaP8asPsV+BbJfE0Vkjn0fy9Uy55D5Hjoy+l20lEB5YHmZl
DIjAiTbYq0KCpVKKg20ytfXJq+KnoLZTOp3sl/8j2wOhNh7KazK+IYBcq/VRBZfN
CNfyTCY+lsy3VlmNFOlOvYG5F1TCe4Hii8sQUkoyg/wCyLybO5NrBa/zAqFUHX5r
mfDIFGqFosxHGmSTzIpvBQvGjKS9azfATCxjuA3n07daRbPwxsV3snIK2i43GjBN
iZw7g7kyJS+0C6udyVzF0L0V3W6SwhIv48HPWSodW/OSBV3zMSt/C0TLzXFhc08a
rZNG/0vbhB6VT94+2yFbaZcjZsdbTIE/4Bdb7fqjZivkh7C/Jtd7l8/as+1xgC0F
fvCEUi9XpCoRvHOtOD8Avo2EfWmkWHGsPlpw3ykqkIBMRNpH+JiRdPuTGuoyca1h
sOPLKDybboJX1Qy//YI6j+5+KFpVALZ/ZJ8Eha8a7WDGu3c2Zc5a/k4r06rPB9XO
7f7Twusvrnsx976HZnfvQsWSsNEQ2E9TQlJIyTCv6J2c3uO23Q9YmvhVFocIbSTe
SKqlwQxMlsUEYb0b8r1KU0WVPbJ20/RgwHxYKYhRXRi/7yaqw+VsZnlB8L1yNJVx
SAkpZ5nVi8dg9I1+URH15lldpMWMQ87vx92TIn7hU554ZyR5tdALs3cXG1jOV4hu
U/94MhRZTy0zNTEhfkGr1fVrrxJ76ZY4KiX24ZEcTvnvlgsyDJ0JxzCY5BIw0gbL
DS3Q9iLroDajn2RJ7V8t+ISWbTiieDBKMen3HVPVng6K8HzRLoWHo61d0CUXoAU1
KtciuTiNNqMlyeXaHmlNXT3nUfe8hJkhZD4ypF/WKNE6opJALQsemKVSLMwygcoi
k/a7RewOSZ/Ly25Csl45JpMgowH3WRL5iylPa4e3SRnRg3KgGaK1G0/zYxDMORz5
zZ6aKDZSbnHYi/z5cXUgGrRsJvTQgKyD6I0x0Yc/fVLDWmbVmazeW5EdQEotryK0
aHTN0aUo8PufKW8cpwn+0fV8HQ/rci2vkdhJpupMsKX69HyX3e7ANOthCwKD9IDB
OOrC5eGjptJ40/9eNuIycs1waia25noDL1ZQBJagSms1G8E9SY/WX5MIq85noyff
2tVQ1YIeJimE2eF8aY60BI+MsHTNVKhQlRoDITzuiRpdMyYFDyR9ZQsKlf2mQHT3
2w7QuOhi7l+xqAIC6SLzcnKmhRCZ+JyCZF6bZ8ODYr9NMTIYEzuSl8Vx/Ij3UouU
oRise5KnPHhNgY1B0KZcr9ipNysVlk6aAptf3YIugkXPvnFtomB4PltNr513PSo/
lkjCww115gA/73MgEMCzwTDygd8UEY5OySoh6jWNYO6U7nob1KvkEsifuHcqXPM9
KWAYeP0/hkzkRN1fomj0S59DxGPMYulExf+wvAx1xdgC1nXPhSqik55oagpBxSIL
qmwMtnXqtJacyd98OE40DjS2KYqOGtnANsTMMoi2Mg0mbkpg8m6NYahqWqwZqzWC
hA1+7iMscXGM75Wqqr52mRmpiNtInKJo63O30sZ7Y/3Zvh+SQro+7s2MaIDK6DnN
BmQ7BHh+Uv5gTYZHM45DRIH8HdPzMYI/OSlMOYePh2tsIHs+HaRj25oeB7Yh977a
Yrvv+k8omXJzbA1nltq9KkLUq/H0e2UGK0PCicdLO9isjiGlIQqWJUiDnMEsu+fe
tpBm2zR0YelQsl1zLxk9Oa/zvT2G3iCdCnrZcXWmKi0PXovP90jOL61BW9sGnH/i
fwqVQu+Ih81RlwCXF0dniDSInUMUk6BNMab4tEe2+dxrsECwSPNO7imfux/pIu2u
guLWBJKkLcEeyHMwSUaQeIQhZAEd1O6wHSnzjdGjwXu17l6qxo0LdHyCI342z30F
EX0gsjC4zOAtMso25+CuQb5sYht9kkFrhlI36H2cJ/3k+JYHnaZGhVcLhg2hFAgi
n5nU/jJ1vNyetOGmulJClrbJrtyyK1Y/CiGHr4l/19l2amspHhFE1PxhqLQeK0dH
fGr7O/vGfUIuDg//I8qO9/Z9QL5Xw6JaqWTb3s3BpuYwBwMb8kRn+Vw2iCBIXNz1
kWB5LEiW0eY88CEeBdjfzg==
`pragma protect end_protected
