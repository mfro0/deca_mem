// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F4C5DQpAfPRnEAL2fY5Cut3o/CuP3xwQKls5si76dbd1yIzgn1UE4uRvA9fKP83e
/DENr9OTYfPqdw6syMWJz588h7X0mzpj2I84MPQudWC9EtUcmT3Z400Gw77B57d8
cQd78EfyA9x7s7GeNrEJbS6+K2j9xQsIdwOilVrfp7w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18864)
vU4lbA3zNOGLN0ysJaYv/JGp2upmX2vgjFZPR5PU9mQWX5O7MZsyDHW8ukMhMtm0
7dxtTZJomad/3pZuzQkaRSA5JAwHZhQ3PkJBQOmwjt2kNubhmtqWdY097bpYR1f3
pT5PEcnRPc+fO8dJAOIbNIdKjqiL6h18UhdoAX7bkTDouVKOapNEfaFvB89OLI/o
oXQGSHj2BpKfrwfcRVwdsi39kGApX+QITLa2ggRaJoFtIvaL0t6ypMtxMABYyaYv
Pm3UAF5briVOyZHqbOqS8wAmw0w0DlyUq/4KtdqT4NzFpzvr+u9xTQaOmySQ/SWg
9BWtK96Lic4pjznSaZJvvlmsMMpnPT4sMrT16Sm05bTQLSpoebd1AoxoCIvPMBAJ
BD+MuxsL+1qcwdSj1+4H9+nBxFh3TtCV+g/UKBgAKGFSXWI+70wq+GYIdl9o8qm1
hDO8j7addkgmh6nxPoxY5PdNTvuS1iMpWLUVMTXqYLNF8pRNvcYQL3sh5zLC2Tn/
/7qj7J4hSd3FjALDGXBmV1Iu7Tlqsyc/Onv/Z6T6jprTYhU0r8y/JUSushX6oA5B
QQ9Pd5OYDgT1krSxF/Jz0UeJ22u8uLSliM/YNspJHr5Wb5UXIeodokX+a8xKv3zy
iiQiCa6DpalmokOCHMODmrp6ViwBGGC1YCjFTaRLzF9O3fY1r7JTjfFtGWA6W6TK
Vdd5GJ5gmiMVFYwZMpyDHNVKdWbhWOIMXbodffIUzulrXVfo9xyK1xgN2dGtaTrG
5Tt/X1lkKfSy3BJ7i+ieQxJye19bbYNiOwtln127BMvvCnwr5SSI01NEtC/1VaPq
oGNi4MpcLHqXCDjCNK87jpN3WIYLksqwqIUAi2QZiRuAXsk0CuIIrxjxPczITLy4
+FBncN/1e1IUbNtyvw1eUSkgr9WJRU4MqGcmljxkvoMqml15ArsV0PoOj3q7hwH/
GtLNmq7TeA2RpaI2jZ6jfiPJjHTpYuhXfULMv6DAUjtQzxV+yluMpHsn6UrJZRB0
Pg3tWAMxBEA6p8ggucLIRlTx/jLgt51C2W/WYM8zlfhdeqOWg4YMaY2kmdaBZMbc
5RsmcaoOmappVzoQwFtdqlVsTa/bneBZ3jEW/AB6yMBMsEn2+1XDZG+80wJp+fDu
ZrgeYuwdhRBBWHNeZN+w4npZTOXns3LkSPC2BxFMxkwCiqU+w71X2inFJhurCSJp
xcxSYhgC7F+JH2zWuOQuqwwv+zDfZAr96cAoXU3XL5X7s6Qe3f+TcBGZ468Sv06o
QdaSWQnBf6LdjiRW14rKXubqAZKrEGapI8LBYijbDZfJrxJLLLhRKKz02EirHqiF
jnKZAJHsF8YiDz9KpAU8hpO02ZqWwjuIBDmdZxq3/+5Hj9I9aWhN1B1bJCfIVkoP
v/o83+3cThGdbHehxEbnt0t7HEIc/klI9/PwRJY5HYX1/gbD7bUAjo5KluOo6GLb
NLKFiQzi25o3ao0t+meGlxN/6Yt3Q13h+RpfshTsYptdIG9PUtGfHptW8VNO5jAz
dPLl9Yq4TPErbK2koRkuE8ufhWEwXin8wnCKnLM/JkJGag1ywp17K0ahz2WN1Yew
rfysEL9U/mXw+5ivdZ1+jXrLZtLiZA2mH8J+B3gXqEyli88GNhIq287S+rAjNmdL
BJ2EjxOLsY6/OyrpWp0zFABT5QcfygRQKkhI9QarUm9AB8HWjVrbxuCz+Mc/m4ev
NcQldIrPKb8HKr8cSI7povZEK9M2/L7yx+fDvq08v42lxtT9IYPEwtb6H7c1jtih
QGbO16evC9orOBOfKwYVbNBdsJsxvz8qrvT2sut2VrIR2PpslMbz5g0QZDx0gOjY
Qm3IIJgSoLgSkVYo7fxHE0xY8I8akDEGtaZNlTICpmAajkSmgZD7VzHi+aGVuZUq
M2DPt+LF+l/JxQPHsNn3dnvAvdql4dN3RERb+uh233MzsltUUXCyCTn/BcaNDLxr
cCFrVsmXLmN3Jo/XuprZ305CJOTTxnPHserYgFXJCCcXRdORRWYmHTZ2a9WVJyMW
BicEact20GS0B/YQnLjJLgfIspEz+YCyvBmgIPBjuIZOJalKVWrQxJDeLjxfdAZl
MlNkqldehLeQ6qqH8vZqBFyfcHCaZg4PzjDIMsfIlxHExiBdzjN0eNWiGUqQs7bV
Nk2DbNwGpXiHJGXEECwYiBbnar6dd5plcLrEpLzDYXQ5mj7xzENmE9EK/0VhT5qr
jtDi15/HsL/sPsayh6OcmcxbHWrlFYGgKccZDwU+LuXOS1VY6S8X3QGCEEnU8eC1
APDBiVbvnAKHI6iMl5At1BDEnLebg9sd6FjmO+m+Fsi96c7yQP3lB/OZ6ptD192l
tyJkDWRnE/qtzzCOmnbKnH87hXyP/Qt5/TMWJ+okMqn3h3jWsRQMhZzMc4yu5iNl
bj0izEu8CENBlDj463HWnjaIfaAVVCNi6eqAK2Lfu3nRhc3CPrkplKXN6//OZW5h
GSaZco45V9BDDm/E1D8EtqqYTtJ1ai0ChUkyAM/I41gV4FQ20I8ucMbSaNE9BVwq
JOVAMQiqT9iIKt6pG7mKUVBs4JHxOzBvClngxeUsJt9k6U+nIe9iDGstW3t6CZqm
KEk4HGkkwysnZnisZe+SjbjCAl+186PhRD+Gf/MmdW5/HZReyTTx/xLXaJ/uW6BE
Dx1JTuj9wVk+ris/i2ZlumAufGM2luTT5YOO63CFpOh9T5P0updTWBJe5Ff6CdVQ
07Cv7TygrzXtCsbZR+WbZrPH75jsSSQlGMBuNwdR6h1FcADXdi51hoDBIjrbahwE
hbxSPvGB2aN8vXwtSqrDlhT33x+6kh2pq5ELjH0TkTkzGznhoX8JTwMA7RFbFr3I
31ECh8zyy0+AR07aUVCTo9IuwyctZ530aAgLLanCyjvCpOcpJjDCnmk2M/0TSggd
LYMjmL0nx79/Y8BrZh7z33KE24jbcMdCsDFuMYWUhqHtmQW3WDRlWrxjsWsIvRPx
CVO8VpfrKgoJNcQvoWRky2Z5qHoW4oPKJicL6MnLq3hSoa/fYMSGHh1pYlOois8j
XpMoTJmE2ocJxBhpl0/KvpMEBOPkz8N4YSEPnoegrQD3gT9Qf4swY4puvKN956sZ
pgdOXvyDPirK6iUOEocO35UfXna5onwipJHhDKi6OS+FPzyOHue08AzfBnB4z032
EVQy+gdSEqJQ79IZSEusQ5RnraFAhSStWxFsXcSVnWR5Bwc3e9r8g3ipbRU/RHq9
SOmHxU5OGJ5HIs4Mb+r+xarNh3kLo3RomTMqFCaqkwUlb9iZuSUqPMPRI9VnlNsN
OSF65kroVqpkPhsZ3BYdT8V3PJI3FQ+J4apljtENfxCRFijveZXZvv1rJAzCZzzW
/ghQPHGhFtKt0NXBRbwTjw56+Q2NkhG7RGTNSPp2IbBFAdLlBQjKWeFKYXx3DL+I
ssm4QuQae7vOhQ+e8BtMb/Qu4yDYv15j8ggws8JGCSUsjqezyizoSN4A0CX/lBk7
udcUf0HcPcX+EsdIVSYKr/IrZzq8KSZIPsugANAJq2Mdq54THoqAr8HwE9bh22+E
ttj64aqJ+SJqIG9OiPeUlOEFtrbxwZPS+vzUefa5TSTNhpxy869tFkyJj4RiaykY
9Ivy8W7lD2wWgX6p+AScNI+9PCtwJq2LKXWLUbfWnSOA2RRCLT0mGtCZuKp7IUMe
k9Y1H5fI3n9wZSTm+to8a9RDzL1H1fcwHxPDTZMCC1yxNoHgR0kwwLg770hzQv7o
0OY57EhUloXdByoZz2HUUrM86mf36WgiaCi99D/kf11OEnMOUPcpBpX8Z+P6O1AX
xcnYq8HzBJN+o6OjouJzwYoND0SPVGckkBSJbSh+Zhif5yLQiW5sklXX2nySV+H9
v1mMSWYXbm0Z5iCdoGKMJPUMXpyjgKPMh6iSMO9RGUlJ2SZ5czGV7QgtnBI+RYXE
4BdsO4Vdjp+CPV/GreZOasL7GgMhNZsbYRBfyDaeJfuTL8j08myImV/9dx2q3s9b
SBHITeS3NiMD0EUapLsohUjdGVfLw1zywJ9BLjF9MCdGQ+xThQ6nQ67PqDJm5Rl3
YPviG9s2861+PYT/9ESCj4OYgWBKnnFPZ3U5ngnlpaH+luxxb5iGbN+sqvcxyjid
oqDm7mawM0cb8DZFzd9w4KKe0/9nfo7tPFLrTooDNy5KNdpWdmK16oJJ5+8UpCey
wwcUBluOPqQiSrE4viQJMuZ0Yd8qLNL7CTqwOMkyleZMKEen7FZRsFRaarj9929u
v5A3gx80mwQKw+0vipNX2UAIiO3PQjV44Amh39xvZzu0L1DjJsh6EyXfumbT5/xI
gFvcLlyrfWaZOmmYmMV8ATw97qk2esmOQ8kHb4HCQpWuBnW3Q6UjEMCmB3Udy2cW
NDyofY6sd6rXuGpBIW6h3DoFA4+QuQ2nga22V1f691Vn8CD1QfyCFf1pZHMA/c7g
oxLQbv4jbOg9IdQPppWXkJ4aJjQHPivNUveWYYJmQz9w/JZ26rrWzahadPU2KY2A
Xh4gqGzLKE9EgGiJ9+QMJ3KwilcOWEiME7WN9V/dIV+m5Ky3F3Y25hcyeKoI8sf/
YCO5rHQZ+pdSThM6BLtHzWKwc1aCHkACPXH0s+P+6eWwe0EN0Os/5pj55t4AFlK5
UkFGK+Z4VCjkZJ9TvZgVms1j/PKZcY5yg301+8DsZaum9/8QjDUXAYb+qJHQ9I0o
2xzIWi+kUmu4fvKFkUVGrlFwB37EWdAawUdTVeRCPmgpli7t2srQghi1ZAaoMNav
qvrh9ZgdJ7bmJas4dwqFM/635+Cuz3m26IncGmNJ7KQ6BLe4iLhkuS/tOgj67AFU
iUlRDmPavZJR2rSH0sn8Qr76h3NVau0lAQIIZpz+oRv6FYSbBSYjn1kkndPLPrgY
ieBm6zvTqPFIGhqBcSIq0QGFUxlv0+y1wruinrpbYmb32WhHB3651UNtdXbWnvPe
ea00PNkujAU+fZxTBtOEoSzuY9neR/dEb/s6941VHHNpsC2RjoIBrCdkAXWrUiWw
zVLM+9YZ1aPJnpQG/Au3DC+DcD51Lq143YvNeLQXxOtxboQSWnlasP9Z8rTnOq+Y
4ZzHdHKzn9ux/ZD6aSk9trSw4wqVv0rruxGUBtQ0XAKyBVmNwEhfWCGq4RjQv0bq
aL7YTFVaaoQRS/wJCshZgWRTfamCF0QV7S8e8k/I+8TlaKUYVIAIplipDNemV3KK
mQdwv1Oa/RvWGDEcT0YzWH9vILrdOw/a0LOTQnV1Zzh5zGsa9UpUMhFGPdxV7PRs
4+iGweeOF22ybRcfj5VRxi2sK4VSUP1OpNIqFnTkini/fhNF0A69Y1QamIpF4b12
1/URMpj2r+YGP7qrmuyFDXrsLyojsxTXNbTkmvzIayt0WlFQi8CeFA4rRwKS5lyD
Z9dj02enUxfQ2uF6nKxgy1ayQgrmSzaDW2bwi/DnNUmL6fNmgYSF23mEnD8hLwrG
sFsqDLVsJqJdU+tMXbreJxnAU8RRp+5lchUV4INOj7y+G5XiBh1xXDXSfDOFIsDF
fcMdaxs3Y99F69wU/rVyVYzhReTEQnt7OuQYqaBMouyEqREihBJe2P2uSEOzspNz
iL08fzzNP0DEGdtOaMjzhXzUBBhIFno4arG9B0Qx0DDVbW6pRY99dQexqVNPvMwj
UYq1nzpe8zFrlOhOkg2QDPZNrQNXyZRGmW3C8zYrZghjHNzv92yG0h2ilMm/wnDo
2AmM+yzcoE93dDMgiqxOjmZCmPWgXokBkknBA7oQtNsLLn4PIIrBcGBN3n65Wu0D
ptt+7sieVPMUkIm0RmT85YjVFfTVY7U398sp2GUv44EiUcnxtydq82t02qGWmqMu
JHEUQh4s6XlTBooOfmWB08Js0yoXpeqhwWmo9a/+LdVeOWIkqyR6MzW/4DyBoEWe
Dx1r8sSrpwaPLjR9icBQUe56IN72pwuob6PceRd5vb+EEX5pLhsX6wRlLGHf+OS/
ON108LmFrTewH9B/QO8k6zC089bpBj47g60yW915EoM1DgJiG/127aV+4ERhkGSZ
RBj+cZCJQ3EOEbKa4e2/INa12rHXZfu4CcNiZpTi8rqnTzqCm2tk8ZPxOjf6AmL3
auC7lfpJL7Tz9K5CqAg0S0XvME9/UyxVut1W97LsHgwZpoUdrlPzk7jAlMdCQ8NU
1kvhwbNBKXF230WIMnfDb2hzLl8C5ubwHQZyGvxgrfEfQnNr+uP1jvLJQYT64Yls
MwqdKo4YSK7/sNfeW3c0850IDNYC3vV6QXCoe236746y+OqeVyueEbZFz+lor1jm
g5tMqh/s046qz5wl3yuYqJ5/3kMmJnY39Ry2jfrAW1fjMzP8ICzTEZJQaShTRDu2
epYoZ80A8KMPECh9GF7K+HtG8elTY7Jvc8D9V70teQqQdBqT3hL2Xr2V+YB9dcGu
aLeXtnc52LdbDHDaVDWP38OF+Df4XdlhR2xgZ9fmV5pYu/lHqcgT5pEucAky8WhS
3SASxrRQv59wbfejg1lq1/XOpZRawFx1XWdt4E9lyyVY7phmfP6LHaZubsrBeCEi
/3S+huZQqmO+SQJoVA8w3XAiVwxKM3kSvMyDJbJGyxvwmNxQn4X5REkdsBQkUTXW
X8+avWvkieg7+yldxfYIXZpzjpB3AEX2zFh5whkZF355PqijVlGJgvxl+Zq8PLEj
jMYlvTqBPWAgzajaf2dAVLZX7nXtmDs6xdM/iJ+4ed5ql6M0QsuVahP7qAuTdhFM
JDDrGWnmhPEnkAtR/wbyOdCzc8KEBSdNU8UjHv37fbJkDupsUZEBgBME2SmmtSCo
YO7f9YnQM0bO4lkvuRSFz0jjcbWn0aHBlCG3fisW8AmaMmkNa3XHlOZMW23sGciu
Gy3JX3X2o63sRvZsYS32dMkhiLNtzH4unpiT21cwjBxYQxXGpLDifXHwSfQ4X1/E
66rk9N6gZ7ciE3FnddqUf8/DfkD4I4kOuaHBT/Qx4mcx3+c0bO9gza9KGHl4zkJk
/+dPVrbaqXmxK65t+Z+TdYst/GtPaAEu49tpHxJfhFfkM/gKSw6vzULkVdQM+nOS
FOlp85xEgpIDbtx8jCwMTPJI0bipRaXEAwhx5Yc6n6oMdy5IiNDvJBsqT0wITp8P
QLkSUb7WfnI/kRJhQcUgifPQAsso2ANhG3qG2zBqAZDVvG32RWr6K0DkH9afWTAQ
pC/2u+taMt+++wFXPiLmzYfCkdA+Ulh9MnVOUdQgDikbzHfY2ugYapBqRHuOuj/J
6VqjtnahX65RC+ErdVIDtS4fosZcjTUxVhqlzbdRLWf62Z7Qn04iFY8dYf1R/5tn
0ItLRtEGZEcn67KrXEQN4veFHD/GXiAOlSug27Iv1ChUx9sObwVtPM0TiHwRlI7R
l8CtZmYeu6EQWSq0gthTApe+xgJ3u3WShiZGpGKRwnH7ZSz7sqbCJtsNhn7GJw2T
R7OGtEZHDgt/Ey6ef371WLyA2nw/jI68fV9usbrRJpcw/uTe47spCyy14xhXvfqs
kjGBby+BJs9p0kObXmu9RvCnbdluKo1s0TiYhgYu4lwKJlVGZ61C5mAaLuQFDaED
qBIUquXloBCm0EiSasIvWYszvKdAF4xtU4SxH41Id8S1XcNRxBIwLBcQ5egf+fvr
ingh8ouhLJTCqerDwNNi45OM9gZrzEi31oH7/UuIuD71VCrj9ADQ6P/4RbGLTckW
DfgNlYI0ctky6xfyEDqjQiMU57Q9JW1ofUZ/EktOFlAJCf1WFUH4DdwUCajqQeom
hz3ZXdSZHh5TY2Cne6zFou20a9AmPQP9b71d9gxKmAqRECw+gCxeoPQ2w723UTN2
+9XH3v1cBfRs79XZvU9N7sqNrRzuGwRdCUY8kvdbTHfLHpuX5i0CdLWEPbAy3G4Z
PziyGuA2yjG+dryornZxVIni1Nq5d3DO2hiy5TIx0xjISJ4IYCS9O7XNcNovu7kM
r147++brWpgzK1hzp51mSN90yYxsepNzvYsD2JkXvv2JFW7Vre8qONn4n+XA091p
BuIcCP04j75j2jLY+mvrWDQlU0EkTeW8n15jDTJ9RW1y8Da6Vn3Xad+5Qs60xP96
wWOWrgyhakSsZoBvJy4KcWabAFh1O7dlZJsCBmSXwoij4Q+DLnzHvPv5zAmEpUqz
RK6OJxie4fmQ0ME0vCRjYiYhwQva2AOMoNcA3Vsp0nLXOJjW3G+w1NyOSs+lKNkT
IFF9+pACMw5yUidDrlFejuM+abwJj5REOzYckiAOelSbuD6nAyLIckAMWYOsix2h
4Xi2hecLEhENXjGn/1rNN5mLuc+avCJH4Bsv2WQ6q5cdVOuRCiW6miqh2Pj5kKc1
rgMkju4xnRnj+juQO6UmL7ReXS8H0krhVgB0JLriLrmW5L8IyySpGEG2cM5X4ovk
YoPh2MGHw8Oerpl+zNDaxXy/iKNYlQQn6Y+61oAQFKdZw7ZZFtJJdxd2cNuOAjFn
u772QZP7H/c36e1G4urjTJsokM8BNdyaUSVc3EOLgCAhZ3Zz9I9gyIHG1vik8nzX
ihfAUxX8LqCDDQZHy8yT/QZ5N4lOOqhRvzq2jGSpv9jEokP+qL32m+GxKV7WaEQ1
A9lqsc8FwH/FMxyuVTr/S5EeyXf6P3/42X4rKU0zlnnSYrw9YK4OsXyylnQDC3yN
n+zeZdGjw9FDeJirQGh65V2M9LvU80CAlMEwLynd1RmTQBQjnMUcAAJrFLvhvhGa
q8KaFAJvl0DaN4JZEOJP+DOBTmFgMS7nATJZRlpti5jPa1cVaVp6xrxe8XiJu4nz
aVTMtDm/zD9lvr5/nZQ1B+Yjy34/B5FYsJOzHtFjjbanWyaUK8lQBA2LpBWm3KUY
JnLAobKCjxB0lfZInJUPFz9pghnu/aeh8VOz98L17oUK5hvavQi7vch0QJWXdI3b
vUfv4nIColSUEs+lOgGLHqePBJS9fUKqr6IhdjzKGK6nRqDux7JfmoR+3RoxWat3
voYLoCfGlGUK6Q/is5jay4hJSzRUK299JeZHS7Rwn53kQo71ts7afMlOk1ju/BcV
JdxxM4ssxNZRcQKo2G1tJmHKX78EvMAnUcJ0gJZnJ3GmqdZLfkr7jol8zlD7KPWa
BGozBLU8wPLqVQ3ZtRrz1g/TAV3h7M4Rieczr/weWK4KbBq9A+SKlpUmumrEMFJv
IldX1fnisH5skRf+V2OvRLKdTcq7ez79g5txiwY9GcJhzHJPFqQwRblq+3RbGweS
mqVTbmve9mEkNiu3c+pB110skZDwI+kVzU2KIPH1Y1C9FsdUGG74WoPEd4+7r7sH
NJw9p7mbco1kSZV4UvKVne4CgvN8uQQ+70nZwpwRT2PYH+9vOnnLTsrXR3lAWvCE
rjqTxT1toJYxRD3aRSbKA3zFv4QcIiQ6tGi0YswX+KvRvY8hPZOKPuzaI2pzr1q3
K6NQSwMtbkFgeZ6JisifMujf9dx9dLWDwpmvmA7Vb2fMzrvw44KYC5GfyDgk1c6B
/0Pm2n/fIOAnI5R6DfPiK2n2sIlQvAaAX/mLMG+hwJztpXp3jlkU+6Lw9nwTMZ6I
ILuOk6/aHtv7EZMlqMEVqahTLUDzb99c6CfYd7f82BAO7mKUARu1cwuyWsCVQo4l
LTDW4d27yNWj4SjZcTWoLN4/+3RaF6LjNv1Crk4yOn/SgAj77qDG5PJdIfgKEPxQ
hBvGnH0BGW8lZjJf5+DQCekanHPZi6pVjbC0Gypuda1qV/RL9EkNkN8UUbZh7Ayr
i8Sb71o8W++Iuejum+HrOnE3JFuMvrea0+Hq+1PEWGn5y/z/vR00R4OuAnU1Xcfh
Q88Ss3Qqp7u7M4BPog9s9oHHpcYcqlUaWHceg6j/BuNRIgw3Bo8vzXe07pKyvV2C
OlY/dCd3ENFgqjVp8KGqTpbeg1/5gf8I2ge5I7/YFfOT73M86Mt3YY/5y0mZEkiR
o4YsJGjUDU/uei7Zl5etscKzB5wy1o1o182bE/TgOvFT1+jA0Lclr4JEGuaObf8/
9lj/iKaA9ka5PxJZaX1L4NH3zyitmP6m8UOogR7jkUOr6dGcazv49bao+6clu6Ym
u3QvcJDkDRy/vALamapXIzY4Qb+UO/UaXdisY7TU+ynTYyJc/IT1uCtkpprtuuAL
dV7MBEUr8lPrI+jf8U+j9s6S3BqllRlsFqTAmtiOJSa3dSdkF27CpA9sEey7K3Su
SsOGY6GHd809k34Mq/jT8VMBK/RQMLMAw6uGYQ1qDE5acRUJmEVfcmvDMicKBrV0
nDTXUsbEH+9sTbM/GnuRE91IDhfEt6TYw3FxeLLa3we/v3WmdaEF5ji/hGHYFpI4
redyguaI7wgzcTRiv2fnFavEMyewDje9jAHayRHIbPYZP1MF03CMyZqVuoDRX57T
9MlWo8mspXnrwCIxSpnf6ALxf+778hApZAa+7hzXjlRc5rQl4gFVPhHZM2bjPruO
5lcbWOew8cdoO6sX2wLsosk1D4qAKfwqfXmFPNOz5HPEwsTq3EyodTg8buH79F+F
SanmyPVCxVesvnzGWdekuc+kLoVMi//zy4pQNMmRE0dRReHcup65wPP4uczf/tXu
gv7PxihCSEW90EXffeQIkyOczHwJQH9ZhdHJ4yDNngskFJUqVlEp9tKxsehanqlj
kTKJuLTm2DTZz9tJW/ElftyVqSfiJw2TXRH96SrLJ4nvQtgk8ogJ95aDZLjPa0Q4
YsZaf3p18w3+hyQZILPJ5vmKNEluOLhR7WN7c8ByrFvK3K5eXdf6sSlrGITJSUOw
VH/YxpbaGMsD5PqIz+wjdrIOrh6f2i2T5E5NIOBrH7StxKXPwBhD+e0ypobd6x1b
hJUMbsuwnE7W5QOQghntemdRc8AGFZ2VxE9ci73WielL+5f++4EsxGKBDRW0qtmx
q2ibeKqo/a7nFTW1cylpaewcRkRBBJaIVw1SOuB1gMFGfLEVlNX7Z+BQYZl29FB2
SDwgigeKpQWbfCC5omZf3Gxj3KHnXRfItC5RcWccqQDsKkAHsTqgfb1fpcefc6jn
05wi4PnqXdMe0mw71fhqvBnFkRFZm5ryTWljs+kc01977BKhOF7AIB5j8t2wLHeu
CAC/ttNoZSqErZ/gOunWaZIwIhO+IY3u8NOTrrIMp42wHgJo+M/hBr1DgpSsBHZr
9PCI0fnRKJpD+2u7wJJShi62di8DVLPD7mnLZgF5ml+G1twBkHVCkIMKeo8fL9Ut
qOu6Y3K+2Z6YgT5bKVx/j9OWg0SpOG3zmzwVkk+noUboRk/mtSCTMFtJeJ+AvpfC
CD57OFVvJMIsXZgXqFUSkHYREcdbtXJE/JcgYkgAdOmsU+Y9eIVZ2De8TtG3vsWP
Ck8dBo6eQ/tJJO2qS28haDYwzxYwUbJa7SHBhoWbNqg0B6Tu08GTPsgeD8eHLkAL
IhWAtwi03NQKDtotBI29b32gTBp/lAq6msijXEZuYSby/5nf0zK74m1CohJGNM+K
W28EjiNunyJVZxkXWTzMEz+i78SE1MUMnZs9hs6z0ZGu6tPrv0Yj8ty4FhiTgSyk
jc1Y93XhTxnaAgHeneBo8wRCkAy3EUg1tlYwdTBV1MEzJSZbnbN0iXNsvYftTlfF
L7lCFCaGPJv6Usn+FDQJjfLTMqvW+jz86S8w5lENixRCRJvmYHMqokeAbX3ttVRi
0St9x0pdF9r0z3VIF8G1n6in8uS81BrGwIBoL0HNlrqntsS9WgGcDgpm//ZhY788
Gj+Id8FMPyrzDvRSY8z89AqPz+/01WXczDMmhRrN4DhqkMpnl6wgJA7nbaBM0UYi
eECkoxbpL3ZJNT1JgPGuJ3TX8YZ8QzmMEnC/m5HMOfuVrcVm7cx6A9ZiFGubcpjm
lJaTdA7eBZWyJlCQsYC+s61vWTJZLmKb4RIYEgvj+bugZgiXo6JAqAUAYSMcyypH
uQOt527PjeEF9LKq4Pm7AkSo+snV9bEla7Gv6eDV/1bnVfbIHxYYf1QDKMLwf3b0
0M6+wFN6IBocFeuD7EPAZz0EWYSJYfniCsxm1NNfEdvCGV93orvKSikDwQdjj1sB
wuRBuZQ+93NeZsAm2yhJfS4uJdjAu7Mv2Rm2R5p0MPZ5LxhOcz22Nc0lbXbzEoF3
2l30PRLysMlIuEDtySSEZ06G2lnVP3PGrbApIczmBJ0UZX+g0zFzjvWq5CdbZnAr
EZ9+eh5Zwg5JvuTwtFJMOgxpviMhRgzlBCrX254PS9L0hE3oB3ZdAGFlK1ABBa4y
rWTzrkR4+QbGJHU48g61LWerTJSh3O5JDTbRBuqwIeTJ//L1cPek0SOax0B7KtmV
IhIY3t2VeaeHwcRjI9uYJI8dOABqZdy79BSPo9bMLXaOdoFv7lM2W9pblAiDnYc8
BAa+G75lFiU+CKMsUE4EQfX8oJE6ctzL5TgeM+ULoqXUVkgzSJCKnUJPoVZXoyhf
9sC4iHNyrrwEaBpPytL8T6F2Irz//dkwycFL4yOH/KOeA9MO3vLRMYA/dSJ4xHAU
pLDnts8rm8Won55kUkGEnkg6/sMtJl7NFmWVOnRjqRZWkfxufo1pbOhp+26pBE9Y
QwYZPG1B+nDR85PaHwqFvEE5mdaaiwWAvNzj/caqJMP0kSnNG+ANK4stPcXS5lyx
opl1S4BiaUz+84/NTJ2IxQI4lN9UUex3zvXop2wTg84E9axBPWCz7EEa+YnXV7gc
naocpr2O0U+bAooAjpCCyi8PEDSgohlPAr8RPshPlHz5BFXymI0Vek4aJm7FiHO0
tcfKHXlHNF4kTyhrJHmkKZoya6xoVMPbRvbQLhGrrJ/HUhK2rWwMdZbOkxDLC123
OJA9MFPmzjzJOzs26yN6XgqcKsCwgbjHZWG/5/YTs+3Jqfpk2omaj4uB2427A8CH
MI1djNRTbVLWsLwj6454BfNPBGz/4rrSt4vMxXkUhksbT1J9nxTpmLIfMCFfHwXP
TwR5Csb13fElyOFz6/m5F8c6DUnOYFFkVu/zw5148/64Ge4Cv7UJmGS6kUmVYn2h
790tpLAov1dTuRi9DFB1q6SNrewD9oYJVGTHSyAflmJFM9vw3NDG3rSL4zLk30dg
k5rQ0LPYZxFOfjKoDCzH/hJctE7HwysjegUxQ2GsY0/U2ZZ/nPUMRiupBnn0Z9dl
Yl6fVWPuRNVmkCvOe/oiR4FAiin/lUJMmH2h0wZ8MLEpl2rtw3fqm7ogOZIuklrf
Gfydr+tW0lK13OqXjI3P1Sh3sEhGIPeu9PNl9IQvxZWA4szX3WKKSqeT6bnMEzss
Gx1F700BqSoYiTgEKfKukI598IZhWOzekAY0e4/LG0Ea6wBT5EG5e5m5IOgEe99E
XHYzg8dXeHFBsn2mhCsR656oD5RCxxvtwqE0tDt4IpAQwl/hySgeR6fQbddfMkb8
aiyIT3CbV8CbkA4fWY30f9ia1mc6EyEBiXrUU7lK6YFqIOMlStcxG2yXqpaPwtPT
udcW9LA3ZHKeAvCCSn/SZ/SaE41LHpiWbxujExVhOiLBM+4UtQzKtB69V9Z44kao
hBGvLKMV06SE4DEo1oIj5n8hndcRcP85J3f3STRaAR8ScamPc55dVnkqhZkzKR0N
eXby6zX78bkf2YnUbbL4jXLpq1uMiYRTPW/9nvw+4FTw85VL5MN4R7KravFRUqz6
JV8mrHGtGjoHC5h7Lb1S4fULQlr8UsBAn4Pcey3DpO3FtxHP4gdi4hcK5p5mrxUq
nX8nZUTh9knI1U7++25FuVk0vYbqDtmSFegAZlIpQEL3GGviDoS3gLfETW+SovhQ
kUSek5+wiK6MYfdvCOVL3Y4Ar0XDeh1qXKVLaL5nUfefKL0KGvqRXmQiRyspciWi
GVmWJw554TsJ6AQi8FOKxbAWCKd1Q+tYfx2dX+P8Hg/WMcgIlbonNTPQwcWNKTAQ
HBL2AkRMyEGQFm/Af/pl/oIa+663H9GfK/IM5+uHo7o4XcFWAwjTsmmZygT7IqN9
AhhALYD6crPlCbatPXfnY6UHKGiPdqjGzJQmnIZsRo4fzT6THR2a/23VpPx1AHda
7VaCDW3SpukAKBz7PzCuQjjj6YWDEB60unBCacqqULovfR48lGO8M3HgObqVoq+i
8Klt0bNWrFAJkz/04kS7lIzDBwXOO2tvq7Kig3+UPneyOG2A0ztQXHWk/5WXKwYI
nVGXUiw0DxGWundO2sfMahF/fHSjREjmFc+nCC85uAfWjFKpxHboFbwbSfHMpjlP
f9JJYKabWeokHZf9dK/BRqw5ZF/HI3AbFciTITKDax1qtH8qEJ1m1Yew6bz/QAcv
B/XYRbD+biFKBrSOSal16e6wuOhTkNT7j3d16kPbyl3wDLj0eGTUuuGFHY6D6WhR
IhYz2QbeSvTXghrUT6Nb1IytsUzlHQ7c7NVSs8xiInEp77S5XkKdJxBBGHHbhtqd
Y2dWIA40NrST0raNUgHqDnVpf58uWxn2HXbrXCNO5T3NgfHp6gwNmn4HiaICOGXi
C89DaGbHcG9wusB6Kt/Bq4IFSsQ2uB8Zjkx3zO3/0ZEmaZseM43q7n9KYQd2W3NS
qvmez3uUt022scBTQRqoC1ruHHm26SM31p0hFtgW15GvgBNvyT+sdbtvrO2teBu9
Osp4sACVKajbhH7GcRL6iiwZNCSPUlZmL60zOtPa3kJrSfJP4nNjNEPdBHtJExrM
Gqp63jqcvVPKiRAdDeH6wMPvWIXOVoLNuPYngdWx9pE/Cfiond4LqWbBbfows5Kl
QaCF+DUhm1gP6McPQDXvooRr3Jns8Zl2fycqCkNA9mKnar4NZWt1KEiVuFPu5Y3H
R6u7DdMpQDz0hs+Hj9pP+wYrYAHOwgPRQFSZw1Y3uGOhMfEXjBxtPyILnlbpFXAN
Mckp+qN/DL82dfJg2Lo3QlSDH4K2LQ83F+a84UAiEx6MyRM+CiRT5a/P8A7wAnIM
cZl7XFnR79TisKInIWUabdIS4PvM7y7NC7tzJKY+K0x+v7EJ/fGKMTWGt3iaRAKy
37NKItYyeaUvwbI276yJqfDgE7IospXs1TOapPj06w6wfNxICpeWGi/X3i7jD+5W
0DRBviF4rRwVQqXbPbhU0hnI54UwI6MhNpQu3p2ajhz6Ng07iSCAJxe6i95X3fPq
IGwXMDQayIUi6QwHVEi5Gv0kMpPC2aco0GveAKrWz3XNAwzUm/w92sHItQmqJXTP
UstfB1QWsSWsgTvt0Tr36AEQZJEtgaM5ipMmr/XXyZjqC8OEK+Vr2C/JJBRmIxka
aFl1OXlXgCyxGUZQ4F/lyFGXllVtWLcP8JO328qZCeXW/D+jP30RRdJJ7Bghcie4
RBTs56rQkFEs6h1iXPG6ef2vAV6lPA1UhOvpIpIhNdw6FIqtA5HXniaXXCQSNHX3
JXOVCBNgyPFNcQBPUah1dm17WzK3vlZBu2H4YNYlKBoCqzr75s9DIYLOHcBlN0XH
ymY1bf/8f9y4moZbkz6HX/BwB0WrZcszKWt9M0DubyUpdU/+CcJPLKD+XCtYvo8T
1l8iWktCh5gZRgayUwXzGwXRyYjuPwMNfizclySQ4qHhvf11LtQhZTAGkqiudcvp
WgNWE+RrKYm0ra+Jq+M7B6ik7wQkGptVvkvFPCc9kPNOsbCmfVdsNM/tg7mbffFS
rJGf0EyQ2xRPNgOQxj4EpIbr1OIWr5khFw/CtK5yq1VvMV3P6iBhVUkSM1NyC5gk
GqqeqfBMKVAau5iKo359j8eLYdcuCQOwHl2Lg8lRm4QhcbJC0T+aab1tFhaDjEZf
y6XElZT4JpHHmXtKiLcNXQ5GNs2HtgobMvxinqkbCtTJ7PbMA8lTBSNnUj9ppUtZ
vCOxAGVIRSSi3CISH9z3/2WFMZCLWRw9+5YWbZURTcWZm+mV1Rk/U9mEVtyQLQUj
lW7dXkjGMnwBvNvg6kGOVbDVPUHPzQgvvIlJJMkjvU28+AesTZoOqURMLP1fYWMy
5S+l9zGmb47DEHpNzUwrBDZTKRxxd0mtJSnykHWDfjYKViAe10/xzYo0K9WOcNXQ
iwqmHWYibFMsdmcKd6YLFf34GO7EcMXKzMJDhgp/ylSyxYcxFVEG2lc6eL/EKVY6
4tYaqAUROQbWY8nt2uLEFE0ZqoblLmZoqJDXCjOiwiO/COCoEOk0ZPaARZeBuWwq
D8l+duCDQ77Hci5mo2T8VV1zuxpdz97K22fQk9S8Ij35eSkIw/uAoCo9pmL4RpGI
NmdxaT9rINLOjJqd9auwN7NeBhWULvC6e1be/rGo1gIPHQkCQMubkVxDTp+udPsG
3+WX29OWhsbROeyLX6HvE0/5XCXXOBr0oMcAWXCbwbVv3zpvxkZB9YNp19Ds2pQ+
/3xBxTjxZiRV/OCfU9fvWDm7qc3kuFGXacG5tKoXMELWtPehCgB/05yyYSYxgRYr
movZs9b809bT8Ug6BW8kfzq1qqEIJh6a9hNg1i7+nWrCBveCFlqWr9Vi9j5rSmJh
M5M30ZQt2aMfwJkQKfsD29/KgKqJXNSgUGq0dvdv3e+IBW/TKYBQb+ZKDec+SL8i
mDhTRu9+kbRLkL2Ks0c4JIPYAEWsgsJ9fgsOgf6CkUGaVwv+rdCvY/LGJs4+fAeY
81uuNm16iy3KT1mfwHkSwLg2m4HivslPamAPtzx35ycMnZtTF6QUwEg109gwzN64
RTjaDFVsPieWLDzu6ovZD7rN6Vv6XpnZxuYqvz71IJdLN/h3Tmj6Q46Az27KDfeq
LBeXSlTdBZse9Y6vGfu2op+N+fcXndk98AHUCHjaO6Ha9LAnOhcuCYpm8k5BiRlN
9bSzHoh1RYHL8ZLbqpw4j8K4mWr5O8ePPSxdkwuFE+6HiG2kZyFC2cuMuuiCyRZ5
8wZ4WWg7b0uKNF+mxYTOxmi2D8gqXxpa3nmVMpV1ryjVNG7EG4UVaw5Dn60FIGJ0
J8F5AumR0HhhHKW4fqEPp7aP5EzsxO7sjjotYJH9CsdWMo0/7TChEN9HRSLXhara
KiCAbwMH4pCLjm2RRkDYFWy6EIZUkrby+fY9j1fBlKrQxxo89urJcfe28n3TDRWm
5+N5DjlYRa9NjgqqIcPpcw6MK5bXI4kONlRsQLA/WUStxiMCjdxKe0EMoAJQ3SP9
wTfC2HS6CFFXmk/dEx2wp/UV3UV9HPlZIIK7CDvHJ4u36hmmea9Lx+SvOOURaWKf
AtfEpLXPKeYPK4NFXMTU3gUTU7B1ixaMohtxPWNIcWK3iCvlKN3XuXBrWxKBpTyj
2VqsfSgG3C2EE91awwGrfYlmJw/t2gHkDSvz2M4nX2PNRDWcCxwHW+ieRu3jYu/m
+MbeFAvG+mX8PaVTcCGZuA5WpqSG6SUABrLj1SmR2mmyBbfI6WxeXDHcyOqQl26F
jGfPgktUq6F+T8wgwVAgjOmFLGfMf9MquNnL1Wfa1NlR/CJPL7gNe20pug86K0QQ
/mVY8/XMbCLoXFpMUz8fjsquusb6TP2ZeT1CnryT8CI2RUiVeTnA6uP16UZ2ybN9
HSREavF1QQJG/gV67eUNgBY3jDu+FaUkqtuAbQokXbvBtLB7R6x+YjOiu5dw3v4o
2ucF4AW7al9/8akONE+EiRtpCMOgndOqINKsVrzrWGVh4sc9UDnSLMWaFIF4CZtD
tijSMBSA9+v6vhS76hFjG5gauNmbVqLfyw3kARwF74SqBLAV882Lpgu/zty7jyur
0XtqyzHEVSaUFkK03su1Px/+w6QXw1jjIHTN3NbKF28Zfx6a8Zbjl0Je22rphaAX
P+bwlpiL2jh20SDcWcKVB6XBypjxPwIHTnKFoALTxvz+ZX/omxu1P7HAiuGY+CXp
ihltYDUDebnje9fgA/sIzOn0zc/tuijdK1D1kt18ERgZiks6G6JkGIy+fpTqEo1i
L1vLBQ6ltWHNEj2RqiY+KMIhQkeVda0uUpET8wDJltcVgw13EBYeUNsiZB3o9QJx
17f+joOLdt2K62w6InQfU6pHajXuTcv6GeYv5g484qAq0JlO4A5CqJEdz/4pjGyP
PvW4AZXRT+XOVVab5mcnNdgKiVJ3XnLXmptFgx1DDqsgJOzusLcXAisqj6mIRAWW
8vJvtn8YvDh9LKFPLRdCd1C4NbvtR6W3lpyZ0LCzFdD9kelTCNY3+wfr5mxMKoa7
efcVY/RD0ngkawEzVKquc8ben91EXmRFicVtPGx1BH7TkIdxE07QCULLq1qhzwaq
T7bKNlkDpGDH3Ac2uLPnICREHZYoZ65YYcPqK4ofjlqEPa1bcILkqRPBxJlCotGp
kqlaqvM5h4IE7pwT1YxQCh/Bzq92+Zt51DruGpjX5hOzU9iBuwe/90YUHRndNDjd
IOukvs9uWda5hxvVPVxr14HsHBWZWvXBl4OEbPG/wLViBP3nkEpOuLDS9p6BZ1d4
aLHgysazxaawUqfWPWjJM5EYBhieUE72fQnKp0XXzo4FSpmmPyzmOfAqEp6smMDl
331IYL69mb8DlpP7k4aY9Fcl4H82OpD/9RaaIQZV4eUMyXeoBcmxX4oybmx4CYcJ
xl87df3+VGyXAPk381TnJ6860VNBfFcKX3qxIGpSTXje52KzAfnrmLRtQqC1DaOc
zr9VeGWOV4kCVJJ7v9E7E2f17yulK1Rhn67b9u96ukk0BqCF6hqQji5SkSMLy6wL
ARzPcHYHyz/hc0vK7znx5s78wGxz0paB9LUnIg4/NyhjMjTRlTpf4Rm/VZzxM7Qk
RpwEjmoYUNKSaniA58rIT8crUFPaGQZsakRi1hjUB4tcESyzwM2E9o+f/pzZYvkD
jPa6dnC8TLjCf418L6a/HhyJqQY2HTxKN2jmc3adIKHVOjzV+xNCftLaWYG8CknM
GJXRRHEJxx1UDCgVohUsJCG4IDeqm/alx5vwAATjnGWeI/JHrXUd4X4nc5cyIabM
RHy6fV2MsVNIc6s7h6t3OEUYuGNHl8MpAibp32+LmwaC0V4fkzUB0CvUzB2TWbxA
0jYzEy4YZd0cy9VA5JPmNt7Q6+eSaR4U3vCWmclMxyICUa0UNSa2e55Z8xcmWJ2U
Es02jH4uNOBBZJlBAX3IGUx520A0rDqgvy2CJnOMbi51IM2cF6Nbym/X+3TReMNS
QpleC8+ygyWjzx0VAfDLRKd/sRkwkDyM7dCwnX3KAjCblCFB10R/IMGRYwMc/c7W
IfZ2BNI1K8zNgTUJYpfbHcDwtPy6qwJvjeAkv40SPEj69QeTZ+VFSVQSOnX6jL57
RXmaXGHwmvOK2wC6da60yvok9CxEMH1WGoBDOOLoYmON7SPufp2a2VA8c9QrS/Hk
hn/eZCCnl60AxjCNA5I4mBtGxoP/D3yZbsfPR+7ywrjuSAx2vNDC0gKVw/PpfF6j
luDxdG9tKUtwhao1FB7ocd943FhiIxPWF5EcWezNsjqNvNqcqJcSQsClwG9+Iljv
fEL8SBgKRXqT6PIQa+xfBXIarc+271ZGlua7/xH4+DRBxakoVYm7TJmpczWCjbzD
UuotjE99mLxCcdC4+UgodyS1iwS6kLR0802jQs65C9+kuY9QD1BR3DpdiNwS6nhr
jRxyf8H0z4lYW3MSuGmQUvO2pTwP7sRl/B1GgPCNrAJFTy54Al+2WOcLig7URNHI
UcDDEhO/0QzRg7Xv9GXF/ejSUEa5TuKNdbHlFwnncN7AbvMtghEahLKmJSxysqfn
/TSlSXoib9oaUR57sQoj3xwnj5qFRHJ3y9MqZy8iYfhMcfwl6cj5BqAkdvY/uIpD
OnWZ7MmNf45VeiY2F9pIunw/CASr2apGODSCcS3MAERLgcRlemPySs/lh385IEyU
8k/ufJcytM7pRbcc1wO5BqNQ1+qPdS47ON4htPLa167vWjYNuLWX3RvHmRcpsmlF
zu0xNOWBn5me9dYbpiXyEJp/LLyDCY5WlBHX0COjrURNEf40nmlIjga8dacdnGSL
vSpe+DhiCfK5u61cxPzxxwHv8Vk3hs18oKGnVOrQ/y7rUVNQ2mBkz+JRTTQr2F4X
EpPkkXI/qo/15EAwzImyWmV6A+1R+HtaC+FWMIpTZo0KuPQf3zoSQWAdlm8D6Zhn
qFyRPiC5zebKcGxE6qkvtP5MVt7sb2aJHvySbV1s0qtO5RLqFh+mfz/FJFwPR9H5
/EYeTXVp7SEPyomSPQNr41cMzPrK1HEsQMe8WTQDhWRNtuKt1la8F+GxRzhFYzfW
fT1tMdQVPw0R06Ot50o5EY98imNI6UW0QuXuD2qWtK4T1jasUyrlQLRgROzdBINs
YvmfiyxfcuyuO4416/kYeZMvuSmxyr7uowGN5X88ZygnsSTW6WZXu9INRxYeeLeR
9G1+Gb5dwl+PYGfslErAhi+NZH+v0W27dShsstXZf8NPNPqvhBsX2adaB9dxgJIh
Kz3dx964p3ZwM0PyLS529xwfIrZXmSCxTUyMlEDh7mvoxQwc7spjjeiyilEi4/YZ
NKIMM6PPXkYhjfaznw3LLCG74FC74B0pxH+ylLfDB8l5QRc7HfoskJ/mnVUiPu0F
C6V/GdLQ6fn7jX2/iu2KCDKI7GjhdeMWEFyszOf/ttlqp8r/V7eUuD+lchoKxluA
c+90V/7JlPbx7G/mHiyNWiEmljRZwX1DoAQWwh4eyDL/JGS3qyF8R7rcIY1Qf/Fz
SZ0ZWKx0x80RykW3h2dx6JohK6WwnH64eKzcVITakQDH9r0MalVi+/ZpZjF8uOr+
RpuIGcKQFNPGTCKExREouiCQgkvvlkCfOvXapvOqHoKz8bCRqtuMjVgjrsGCNvXA
RUdGd2TvTQvsNeeJ2BcPV6xluC+39oTADktUsXiyU7GkyKfzP5sJUnOk0bVLwk5f
W8pBBhYmS5J7gCMXt+HYc8FYIqR2WZOR7WIVmaO6RkwFlv8SvOMBo0ewYlFXldUr
gUOqfMoooe/E+Uy0ytXlNTCaWeOTqPq2d/5qb/DGx5NPt1KY+7UC+hrA44WPYkP8
HD3JZQKhHHZe14mlWzh0AiESSqR9cgXc1b/EBwWHmf1zFafvfPUVVObdasb9bd/S
oR2fWe0kdNdONsb0fcyNJCfNHsnCvPDGzK3dzysgd40WujWFaK8wGEsl51B0qfDq
54vBquWSUE1crCxKgjm7coZ+embPMRVKLAplY9mOYSgs2DxRL8RSy4Xr/1xVP/kw
HJnRsXVakCNz1X2x6QMIQU5zqrDqk0ayPb2OwA4ZKH5U7ettJii7MTBG5SEj8rmD
MR9+BxIelYINNG0M7aFJ5ejNsXuwYbvPSmFb8WZjMaj5JVFcW7j4O/vxCPSTboQM
78ZcKSBfrbSa526QUhKhyVasLMPOsd516oPtAb94/yZsYSzJ8N6Rz8Fsnz3Cxspa
OOiKpiln9aLG/KqYTcDbX98wSvfY6FvLbsVk+3s+7IpN8Um1xAtysSPPiS8jQKif
cTNxsxWFmywAzLW19MW35dxM/9clTqffGiD8p6xccROtSh9BjTYX06FUPebjAYf3
hKcr/Aj53VXHoQi0dV7Opdl/Owa9ix8DQOIomOKFq4UtLxaM4C8BMRxvpH9GlKf+
6xxuYnYQFzbC9m5V/pD71Bx3zXfJu3xkornJ0VtAtDKY7O/pm5mCMKu3BbNAI/wN
NNzCfCUZ9sNJQNlANbU+wGo/uZeuNyPOkKkcql6CagwpXZ8rsZ+KXweL5e2hQssl
yIlWyb68h4S50vS4C6LGs0Og4Hp15b0hMfULxd7TP8TdDNpOkhoc168CA5SdCxuq
rUaq3pE+H033qneIN5piYQoNn8rJXi1jL4txJ83r6Gkf4ID8FRMmy+RqPUtypXwe
0+LG0wb4a9iT14497aZ/rZjdMJ+dqCDgxEdYqcvEDIsGw+oCh9D9q9aIDk9GfgjN
U7i+g8mnmG4qVjGnrlGZZfyaTgv+jlbRNVjmZ889/tQa+CKRojh9Ans97GvexDuf
G6QTJZrBicwJ8f4Xu/Z1WVeO3b0ukCT8siSUh02sGIX68wWwXmlBEw6TYrhJXld0
0khgMh1lwtTLpN+KTmRtMgddK2Fn8ty+ySC1avqkz3Fy594+r8CtSiRbHUi5QtRe
QsiUxnRWeylDfYXpkD27/qN3vROLRkKqQb76l23ZSAl6hq5Jh8jrJ8Pe/FillJvq
KQz2nodIiDvnnnJC+dfCYCHBwpWKheEs+HIa2DtktRb5mJCNRcitm94EbraYbTCh
qyyDFpc8mHWJVKJjeUKdgAlh2ceMZXM4GxmpqqKbDh7Bn9JdVks0QIURNJBwIyoM
aJ4OSS5QnE/CLKE0dNfuQJL8A6Hezb17lFipL7kF7pwQTnc2SDzGtBakfWaBrCTD
V3lw5PxgiCwhz+huvttPTWjz1qMayCWwqrleab5ABNNvmwYUCYRRmXPb0qADiLPk
2nIjzwJ0JhQTUx4kcVyHdHBnWYIND8CJClirx1GpxCNpqz19jNHTNC3Yzo7HYAha
rOuvo5I9VUrEdU4ongziLjb/px/PJ5d9891weuyZCYvN52BFCQ3GhyMftImWe0z7
3OFegZlNN+q81jyg6J5c5m+sJiM4rTnyKgnMP9O8jBbWnbLuiZPTSQR8rgc3c2of
bJ/+KhkHIXJ0oWYXGr0kga1MPb89/1oKjf43DASRzVCSQXu1gBwezgi6jiSXVFKR
d9OHSo0IHL0SbD/BlOMqyMa0JSrjBvRkD2i0OvkXbcJ8HCr20kVa0wDJdH4xq2Rr
qu/qeV3SfnSzTt9qm9dnbw7OmRLIQwt2z1V7PMKr6zabcHK3TlclX3Vkk/wcsdBx
tUGi73McZbWtngxYnkepBL+cHt7b4GqT4dVh8lwQocLIPPlXAAggBHRN1HCnY/IJ
Z812sg2ntWXINPqscT04qOPqL7VU9K214Y686ZmSrqowemNnLVgmd0YQ1GFNILnG
mTyhOC++wrwJi3ER7KheCXU9aCu+kW0KoeoHnrzlLUEI/9fubJr2WjRY3wCSFKpq
fmv53Z8zG3RCGHtdRFt409Q72OQVC2iWRAEf5pBRKsedgqyW4PosHkcgTmqufQ40
EtF4wHKDCgALVAKGmpywsxDt1KzQPrvxR+L5W4SLH3704yGY8T+eSyzFAs7NjFFm
5ChJ3Qclo4te4q2iBg/ItqhpeuBd4gZyYkpITHih52aLaXGvUVmhWYsKD4RRQE3I
f5GxZrPhr6mpZHURBnQaZu1OiwBYWJlgwYvTZ24sbn7hTpAOhQGKy/IyRVHBPPuI
7eTTGmYG+3h7z0QYomBykOWbg3y+erNPq4JvBftEF5gushQGnYdmngRCjR0T3GxN
uLa3JSwUg0nlwM0TPwBb9O+sK4k6LuEsBJ1SpLqKnPFJkDhBZ8vMe07X0vcc1VzG
yABRg46uOpEkAA0hvX7/kE0FMG3IuHaSpt48aKhexzgVNkfjTBV8TJB9M5X65SX8
ZeglR2FiGHpeLVHLK65Kg5uZj697zk7NwLn0x9Z3zupWRzOv0dlUAMnxp9PmRg51
22INBl7QnpooztVwznLCfjybXq6IKfbHSrfaMMBKCbWAU3flTHToeIawpNwd7sjp
p8dHWndekpqTSRC9BG49jswM42Pbcko6S3/rfKqv0jsOjQEo78Z2jxPKE2rnlLmB
2oCHDmtbg4CWG20qYxP2YN99ZVlT2VeyC1asoHjIlk0m/4uQ8CS99OnvkYs/RcTC
JfXVDLRiEWXfgpe+3G9j2BZYr83cu86t+Ad/Nwsc1vCyz3IhTUCV0WczLWNj4eLJ
jm+Sx++tKXPfXGSBjvjbMG82Zsum9b9IY/18DDn0B0Jo1u732ILUxz2NuD+iPRh8
8IJPGoMjr/sMB1zXr7DtDdqyiRHKHtkByyD/KhHwHGjtS0WTHK8mcMI2AfxiNFE3
MoFM3rnXyZWPjJY8PJl7pkxVv/yKPzSlXjfYPYBAhJ265kUqqmp60PtBzrpT+PeD
hlZKTSrSxQmJ+a9/KuURDV2rQXwWECAMxdKFjLG+6548RzrDVMIW/JFcMCcGJqKX
SYfeJfJoLp9dx+2DFlIapRHtw7ec9Pvrvk8sT9iMCf+Uzu9Q3h93uoBZAkJsPH1O
51fGwvbMSvLEj/ZpuYSgYGewnTb2pIRKAqvIO8QoLqUTj3Rczd8y7qjB4XyzIfWd
NsxjBnrnQboJ5lkJQgohTnlTaPcXeFSN7nyPCTwOij5kx9oulJUL0mtA2fJM3bvn
DQQi4DWDJoFdnpvUwhmr9w8VgIfWgD19ffP3C+OHkzZoLKTYA1WC+vBIMVmBWU0X
LYQ9sd52y61ay4DbOir0nZbIPd/71A4Gm9JXiJfCZ6qI6/hwOzKw8jcAKVPQ/pNx
9HYf8i0bdaqI+hySjsWSGvaD8LkKuYCRLUuNuarZl2ldgGtZCmppBmT8V3JRon+8
djWFG3rgJKjEqf5JZEoQOkG7Q3IphLDS1l2XOtkwnGPLmtNCcTgYnwPT2NkIWUI4
hl84Xbh09Sx6G3RB+nh2w55B1lGf4PHPooWNc5wD5st+sBb60uqGUwLtNOU8WIcB
tik6T6qjruJy+Xpa4x7ic3AHnAELdLcfqekpZYHmBHVFW4d597Cx7oPcpdRdFkqM
SnGKj5IOKs+4LaeUyhANRodprMsBImZxQWR3PyTmqYZ+EPqtDrC/HPIWzvHTtvXz
m4gisaRrZzJ6IgWtalTtN/OlmHm5so0jkF+Jvg6BtVDb8TbU/vRWdQoH4s6hAIdb
yKnEarCoh5f8akEeq2cTrD0ekP3dmObSvuHmH9pnEQo0rT+lec1a3A1ny20UWe5u
AiAjzrcSxsCL/B7FliNCSaorhb840uzv5+Fb99Lcqmc1nMFdjQTiL/slCyD/5Y2W
gjZYQieH7DXVnxGdJJnzglsdGlu9s16FaV8Ij93vREUhbzbhwkUZ7vs/iv7rO4RX
Mc/5PU1kCcfhaXY8LezWZdkU9NKEsfwvlqNC0IWpt6TwAf55IjBBrS7uKznFyn1i
tHRxU83GE7gqcpXZ/n+wl2mMu61rqUW4N6S/BFetak5ZEEZm/dAJcchpqHkewZyc
PVvxBmfKCJZNBnFPvdSfgs1TaxOgqniNkLcLhavGTmeLzheg3GI8Ehq/2kTuz8aT
8iQBHQGIaFCZmc8EK/r0aChzjWpJl7rIS+pfG7aqYvoLzrqfH2agJsoGSUuGEtsG
`pragma protect end_protected
