// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HNW47R=A01$ZO[MCVO##B2XL&GOW^!3 0?-9&/;[9B0H7#15XV"MW/0  
HL<,=M>^9,?*O_>_.HC/;5F5!4H:C? 67:$S-,WV+>FB2/&VO 6H=M0  
H5%2>_&4IY$S83*!9NMUS('RD?RWZ4\6]VH/%'J$ST!6D@4%L[':RQ0  
H4*717.#14LQ7?\OI*IU@%;%E^5M I$HR&9E,^V)ZR$T+AJI4&!8E7   
H9G/+/ROEBW /;B&8DH=EB8PM,"$0 >B-J=[U;K^F4U$Z=\:#;\&!?@  
`pragma protect encoding=(enctype="uuencode",bytes=8672        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@3Z] Z[ +? 9VF?SLE0?%(2M0O6JNI>BXQ8'@NV/E'X4 
@'4Y57SK''GC<_F":I> Q[,'A%"8C3R@KT&#A28ZX1G0 
@A EGFZ/B/"@0-C630 ==M#D!+I E::*[>)XOMX_-\-L 
@_,V!?IWSR=E.^^5]Q2BI97/'BU8LGIZH8@PF%WMN[6D 
@:DVI._Y9!_0T<UX#-JN49FX TP6^D#7,WA.3%KEU9ST 
@KN J%]KF:"\]P"4/U?=/Z+AQ*% .!GY0&YG78+-N#U( 
@2V?N@9PH8M1+Z^9UOA7C S<U!;3HB7$> ^PS)9PA<O  
@;49"?_2X6@^/7,9RW(3],89Y*G47D_KN3YT9VORT&W0 
@YQ_H_I%)+[*0$\CD!KJ)N=DVSS&+NES0E^&USVAA_M( 
@(32?.(DOCO?ZKCIY4[\=WABMN?<]WYH \#8IY4J:H^L 
@5CDSJ-4N3$_;*2-1YE"PG<O]HXX<4H8"B#]&?TJQ8&4 
@][.6/2/W$M'W)\GP/[( <RGH:EWZ4 ?#V0>XW<A_$Q\ 
@=(>IM%^<I:VWK4=X+\/#T9&3>_H$%,\+$X97F1L6J"P 
@VX X^ RY1]OXV$,)"V=HY72>WGHHS:C'9Z7)K:OSTUP 
@;V=\>.7-&Z[??<*"D*<2 4,"A]^3".%1Z'=5(G$5JS0 
@:#IEP$FT,\B7+H3]2%8,9^910%.1'V4+/@^A"$M:/@, 
@R16O'):T_ZJ(4>#4*Y@,,;7;''*(1X)UEL\]Z 37']D 
@^'R&+FO$2%6+4VP;#?NSMDKKU_M"%*Y6+-D2(85&PU8 
@LP>B+;M>"]R);QG+00G6CL&K4\YUN(1OF%O0 PG1UQH 
@N/#1VJ7LLH:V\S73>-OC09"LV2<YZ/EMT6F*6@E-<_L 
@<A!*Y9 U;%@7KEMT>R!DH;8F&/5JO$?JAH^["ZV=SN$ 
@&6W+N0N><O".:@1H937<R-IUTV/J?2,0&Q-DR7V@A6\ 
@*E%U6L8.,BO7=#B2?[@)AU$-=(H;Q W@G3M6R3<9_.X 
@&=*^;JV:N?NC*I]]XZ%(5S+LQ^+19OF8B:<C)VTTPT8 
@PIA3\Z*91LJII'<(?U^P]'8M2VJM7%3OG5V(@_I!GA4 
@=QY874:NW,)X0W4KT!<P: _R23!1GJ1T/&F9<X<U0 @ 
@XT4@L 8S 21$#T+?E3;K?$SQOWG PJ$8IKF%.7_]*SD 
@'D7[AO[<FDN0U>^C_P!YK_@:TZ=81,1K5/G8P3'D9BP 
@A#4DAUH",<3WX?HJ=(D7ZY[.(6:-$]/YT,I[83_QB+< 
@O[ND9/T>+N5XFTA&9.9GY=2\*PM#?]M<>_;LHI(I69  
@.3IBTDO(IJ'':/:^NS'8P=F0QN$1*LBZR7'9HY6'=I@ 
@<FSA@5Y=!KG\UR0G;/3)2-""S>)3P#, U/OV<-;"NJ< 
@,;D<SB!L=O'\Y Y\B!+2CX? ;=/*B!++1(U8!I'B4_X 
@C]=-4<13.\,,'8P\L^,:&$0[_<><4+!23%RU<GR2&]  
@65@X.HQP8"/KOCHBE*:V;D4)I3@I6S7? 8(0-@CQLT< 
@:!2>E3]M0=%D=3<YN/=W6N,/*5*(TP@=Z2_=\QNQTJ( 
@U\7C[,'5!<P@61]C&E2;O[H&"N&1#M?/K2?%]OP6VHX 
@+&\,Z0M3J5/'DZQ0PZ&4>?&?^U7XR:@03T$]B\SWL7  
@25.6-='&@;DD$ '>*:MA@G8F670KN9=-XWW!\*0NE+4 
@(?M_;H-8Y(I)N1CW;3[73*5 US]C66L.H4=4A:A%$V, 
@= [%E&6/R0H?]>R$3E#W*4D$^M6(EEG=E8#PD_LOQ^@ 
@I9"M6:K3R#B9T#GQD7T%<R3U%9 Z4 R^)^U*RQU8AR  
@_G.BF>S,MH+A1?(OG'0S"_=WTG:9^GB/>=-P@M1SH20 
@[>;DIW6SU!$ZL!5G.)]#7*\;&6:YLGT-\AGX\&&Y'&4 
@W'8EGI?W,,\+4H9W@&,MJJGP6FHII\3Q)U+Y)2I3(@4 
@UOMC'D59[Y0Z4&2H"20:8>KT-#B8=,0 6N?+N+TU&$T 
@X*D/5*A9E_):X#^I[8@<U!%0646>$!!^DT#&(86.:!T 
@;$0L&\BYQ%",C"GFU2TU\--I7-5D'A8[:/T^\O<VIG0 
@49'G+=9'K6+\^8/7B4NC8RCH:JZ@#[Z5@P)W-#H J]8 
@.6+PKE>33M:PMJZE^!^0:1&H]ZP)(%2!&T3FG;[7J>T 
@PL3AYWMFY+\%:-G(B]J)0<@:O]J_(!:N@--/OO&T39\ 
@'\P#M!:C J/<H[1O]S[ .@JR-W_71O#I.7$H 5$Q*%P 
@/(\1]5!2VV90X]"_@_P2RKC:[3/<0D@S?(@$OM9[Z@@ 
@'?F S13?X5GH3E2R.D]G\E-T4XR6^".L)M"Y85*CXA< 
@=2&=RZ7[ ^?1AB]4HOZ[8:BU-S=IX.BD-=9=@P8BJ9T 
@DO=C$LC3(G4:@#/T)'W@R5CV6O:LZ+D@D4;,O(YB%(L 
@"P")7*K\G=6HLI@H#=!#T@!#LB+USS0X!^B9 NOTD)T 
@96>O1.U-4G.W./I<N>7Y-%TZ2A], A?J-$K@:KK\=>0 
@J3/L+BP7O2)* 9]T6E _"K5==Y$_.0EHY_K<Z24*R)8 
@=NE&'7.<5GC)T=I9J5T:S+U ]T)4&M,D2<8E1<Z5(\T 
@P.0&Z6QV34U22_BV3?CX252'!#/@FF4\U: 9C6\3UMP 
@MD.#QR8":<K>7CPG9:(\=QU6;W5TWUS.I=;L#Y.X-0P 
@M;V/PXR7-@.WRWC)]&.C_8B8*>IE5# T8/RE!.7#>C0 
@SE2@%YTGT6%2$QTC*C1?-?ZR!"BW_)YVRDV]#,&]<!  
@B#'0<VHMC)68XCM=+@P!=#'XV>5;\B5J*V<B7&T XL0 
@%=PCNH'3QU[H.E35/4UN:93O]O3G-#TV&'H3801YK64 
@,6D;]->%U<A=YIIVB!O4")(M+G]%&YZAX:L0M^E_M/P 
@^M4E<1K3,K0&6&CH4KW8J>JZ9QRD)W][S=MZ]U'+FU, 
@Q4Y]AO4\C$>+0G7>^V/'@LL&$'G5Y)RC)S"A-6_9"40 
@?*5MN+G0<_'"DW'];PHIOD%+#P_SL^11(24 ]/@X%+@ 
@N'Y+)Z!C@'T%(K1V[L0[Z>9+-^74EJZ0Y[)C<B-HCF0 
@1K6\^?KVJR?W9HY5;8;CJL6RW5 !OC)J: >]TEA/^;( 
@:]D]/Y$-#\CYC%X5%:.?B%45!7$#=1P .'>9P6QMER@ 
@JY[^8]VD9DJC(>R8AE.]!M?GC[FFR-G[11W6JT'4R]X 
@/502%P[QB<YS4I?#>M(XQC,O\<Q6V/G63 >JT<9[J(( 
@Z="!S7C[@:Z+H7XJJ4Y. ;KJJ41%9NOM*I\-+A?D:)  
@7JZIAY0N!A%)Z"]!Z,%=L,N\T/.3RP5YW\_V$SJV[:0 
@WF$NT2Z!4<F_?N+KOM0.:CY  ;DYKL=*W.\%YQX:@*( 
@^8N GMTF:74$\ZH =^.=!-P0C)!"MM1LV7Z@G+ IZU  
@SR;[V^<6U!YE13/T:L=.]6'ASG$E!-.HHPV:5-MNIM$ 
@!VC6[,U[M*?!&I6)0SNH$0RM3& ,N/T=9H9#/U=2,BP 
@@*]%=HF:A#ED@B1HFX^4'<]ZN0W ^F?$5@,;F\M(.0\ 
@3\M"4"9K&/=,2C"[/Z%-YS]!%\H0JCMCAVBOQD)G=[P 
@:F>/.?&0HA&TT[!K,/RU-ZUK2P5P[?&-A"8BH?VM@HL 
@4/V"P>[0%,C?3V;@!]U?!,Z#X'[YZX\9%>8^-2:20!4 
@ ;RXN&9S=:3R#FQ O$AIW^4AGIP^+4,&KOSS.FYIL5, 
@7 5-F1H@[WZ.)P0$!/5<GAD--DLA8Y,LYY<!NYW(C($ 
@'E/WY.2EH@NU76DHIQ]EA9,@^SC8VA,&2N@S#>J7WMH 
@OD,E8>TR9J,AQLKNST_<@.G>T!=TE'</Q*#&VT0FS8@ 
@>%9H0G_3*'Y-AQHD15%VD'B?2N#" P&_;"@X?.F*#(H 
@PPS5OPPBC!O$69OT0M"K#RF0?T%IMI-):>;!6/-L)"L 
@+ZB25C*4],>CY:G6$V.UH$D4?%I]QJWN__PJK*N+F&4 
@Q8=KLQCSYA4A(B/ZR(C=<;"5H\ 7!E7JA+C; U%Q0$T 
@SNZ'<YMFHOPTO_#Z4XF/%'6(; Y]@ZT)5V25D>:\ J0 
@)9SZ$:OO\[@*I>7=<;&]P"+1^R%FEY?4HR<O_R.:M*4 
@]PPR2J20HE !'%"UOTK-EYI;G"XEXC_H_.X7LPR%4N( 
@F)TKJ$ NZ57_LC $.Z+7"-/V34/7T^O==OGP 5T*AR@ 
@08X >CXHG'>35-Q]50+&'^=BF3I6G>AA&Q6-VMTBJ18 
@Y:>94@B*AF9C,",@*3BLV_E5F0X<5VX(!<&39IB'G]L 
@&[E#4[RD9ZZ1T7@K05YQ\@5F'4V)6MTF,I6;3LZ>2\H 
@ +;VXR\_#GV?[HE[H/D_DA6B 1G:8E!:YU736,SZ4\( 
@LWGS#\C=\/[HLG9<LD?G(W57TP\C,*(AQ1=\_"QU750 
@15J>&Y"D"L/%UD)@5DBZ:(I@W4[G3H\S*U(MJ2HF>6< 
@FC:3[PVB:&[2&!]%(S8@NW0Z<$7"8UK_::/7^=4&A@H 
@;/BK!:G*7$SX^XQ.=K5^*JUFE^8]#$&[E//8S&A\KN( 
@4HIX8?H"7?"7;BZRL%$>J#<,\*=N2YQPAT6V9^1EK'P 
@G;=? %QS!U=#PS+U>83>5FX,;0?_P%GW)I$!4J$Q%>8 
@^&_$^F'87O^;/^0OR*U'+/V9D%(].(4VELX3'7,SZL8 
@3&%5ERI"&M)+9TF4W<B^Q"1#YIN]0;@G7Y(\O]@8!!< 
@R>F8X\@/^NQ'_BP%(B&B#I_!L<]'BS@*U[.THZE9KQT 
@"G-PW@=Q0&O\%JG(..OP<B"J20>3CUX:;,FOYG.QB8$ 
@CUF_)1BGW;="-%;]D+S:D[+XK.'10(5;JB&)=[0"'], 
@)K&6?]W9 @2I&)-CK9BOK=Z^<M*29B5+^3PY\<$T_TL 
@&7  ?A"8*CJ_MXVJ* LN4\G8:AVT00:RO'E5N.#0SJ  
@FSV(K 0QZ[3.IWE08G.@T\4SU1LF)Z25YM+-5<R>VLH 
@U-D$.](*-8W*7"T::01UD0XBP6/*>R*??$A909D]CKP 
@(\^.^IPY1_72@ ]0'>OPM(X&K&]S($=G(1_O'1,ET"< 
@#I7:MO&X#+L$-KG9T>'J-@_H,7L6=KR_"5)&1CUPX^, 
@_EU3EFIL.TKE5RB= FF&6T4([,GICAKKZ$E-6OV!%GD 
@Y10EFV!0%]D>M(N%;B]SX_S8C.01&ZL1],4'VS2"I1H 
@A0!XY8_<(!C]0KCY"Z_7#<R"[*;(OXZ9IS/)%2SA*3  
@9B266M;*MD5F/CL.!1W,78A-!Q0AK(31Y4<%&_N'^_T 
@7DA/U!JC.F3C]^BZ/;.D[2XL[ -EH< 4=U02LN0"K3< 
@SC=J4*K_K-/7W!$4M2%DP39&)CK$(\G1:K\&;.M&"0( 
@_)C=A!?+LVJ[,G^:C$:]E].%!J&Y\EX#_9RCIWHG\_, 
@/0=4"X3=\$U71/&KX&2=%.D0$M]W[&!A.[F#( 9T0E  
@Y45Z?DDEV&Y9VRN7_C$[K*.NZ.*A(GH]Z8CP1\9'M_@ 
@BN80]2K$YOT,0C%7QXIT)*@\_&H,.S%Y1ZGB'I<OBIP 
@Y ]IGQ6M5S;3)!8C8P.(K3I@6I57[I1R%#A1,V/KJ_0 
@^+#ILPM_VBIX9QAJ=5++: ^0\>;SJ#9**EFA@1^V>F, 
@-H=G J^Z3I6-4TE&^-]3(14QD/[];-O[#8* ==@]7D( 
@0*7).QH8BKP,2_ME>,^GL^L8?3_^8UFSJ7W*507#4?L 
@$8:)2*780R T.S#\!8KX=O2^V+PZH$0(R0Q%]9T65'H 
@]4O7X^C#$S9!SO$=/Q#638_A+4M)29U=@MU\SZ!BNUX 
@%YN_6PI/$R.?T& *-QOJB40'R\?(;8>+!L@32V$' [D 
@IY+0U:W_7Y&!J)2L'=NW#HXS=BO]I"%$4:2@^[)39P, 
@;39%>[8G'X9$3G4-K^,#EM%.7,#Z$24@^;2JVT.$H8  
@5@A39Z@QRH%XF()AU3H2O^%.7?D9?K9?]'XUP#U<!7D 
@'[2>AJF.[^F[84!ZX='<(N*EQ4 \WLRB%\!%QK=EA%L 
@ <:N/)0$P*X[0>PY':'M'<*80P@+H?ID>+/X-SB:6H, 
@9;MGL4";=4!A>4K=- @9"J&(P*KLL [HOH11Y@.3 %4 
@6)L_7ZP>R[*U@>R2^N#/Z'PE(-]OOM<N+TQ)MD9V.), 
@/QP6*P,,>50&F+@N]*2'-F)KS:'GSCULZ>"]SQ_^.8  
@(O*^:BT5W\!#8DO9)K&PG\O1)Y:^(F=3U\^S39_% *@ 
@+PIJ-/;AOE' 7E"U-%XR!.!F%$7R'2WGT8CS"A(/FN0 
@;UNG@8C>/QFA>%!]]6C>VH6%64(=ZDXU"*"/Q&\O 04 
@#@FXMC;MAL2%FI(2+F;W+AYZ*48.?DH.R)91^)2>H9, 
@XD&EVZQ:JZ0X[GY7W_ +Y#LJOWQP9#?O(UXAE=A./04 
@DSZV2;;=S&!?RN,;$\.L&[\.F>Y)]"30Y7"L"NX,3X, 
@O0EY$LTVMJRB8P,=N[U99'W7-X:C7Y!$HR;GIJL/6Q4 
@7+F<*UST*[=>*!TY'8SX.A002)WV2O<!KB"@PHMZO*4 
@/)I]CQ&(!U8DAHU<VKJ>!Q4L)[P@_!0DL490*$+A7#( 
@9K3Q#G@[ JL[V&;BRWRH7+]8W6G]TT7@32+9'?+46V8 
@?*D[="[H3&XL$UTUS0\;QP$=\$CR[)"QH^.(4Q#O?+  
@TQ3Y)(W*2W>_>2H4%B_)&Y0&F;6,P<T7A&(!;$G"ZS( 
@5VZ<I7 U9>KK(5=H'/K58KZVWX5>IBPNW[D]S< 4*9L 
@^"FI]3-81WA\'WC.2J\;N%)2).JKK[LG2$J"/LQ:B/8 
@3$V'@AI/F+_ /G4:2@SLS^31E@)?/-\'\J[K?HO94L\ 
@K+160MR 12J\Y> 0GS<0*]W"9;J52^ERT;Z_ ,LN1LH 
@-\3!50/L,E!  &E%*1/9-VG8WJ @XD97'XO6)Q4/2L4 
@Y3U??6'^UPJIR!:O,\Y(1YP\!I@%:/T(,(MTQ0"B)\< 
@N9<"0"]X"RLHM>JT/"F=KU/U>AF* V K-AC&'^PW]%P 
@4]^4\WL+0[92^"J\BH5[AMLX?[1J_=*8GND ^V(VLFL 
@AQ2/_H^ U<HC S\%<Z-3;WER.RW$.@;4.G>QU.KO:^X 
@:6I>3B/5R%AS+>UWG=P]FSI<'+V@H.,1XQ2Q"W0[@8@ 
@*AH]"A@76:DQ@/ZKP?D-J*XV>X9HYL(RJCXEAKLR=B\ 
@.A.UFUM9](P?]2)K1^T<:EK,(.\ S1*CCU:*RZY@[=L 
@ZZY[T\&6%(3XI);0^$8?:[=#B7SP3Y+Y(=0>*""X=U4 
@A:/JF$ETL>;G[%C%N&"KVP<8[<+K4/=;&<1V!(9<GAP 
@DSD]Z(Z:*'Y%$Q,W7;[P8<ZZ);].IA["F_Y]*%":VD8 
@>?I_7"IO@RFK?:87X!9:;VOV$Z&2CNV]% W"(AR_$9\ 
@=W%-E15Y@Z-J=?YC%J0@GV:O6<^CYC%)'UP\OC+$HD@ 
@Q""K72,.'5)?6,AU/*;E&GQV#<//HZ;[$:64/H4)W%P 
@NP 4352FV"HMM4E+N:<ZNF/8Y T)^Z=/V*V^[%0H2'$ 
@SW5ES-\-W!S"X5]J48<IXY;;H,N9*^H=9#70=&@:,3@ 
@[ W5)BC"D,(>S>U<+G>_L:]M%[LL;NB;?W\Q4++$86( 
@D*(':J7D/V.9L]MOV&O!!O!W$MM*$>+^ZOL9S<TWV8$ 
@=-6,<($>2JFR&\,$:95_D2,7;,"XHQ':G._>1%0;S5T 
@05BDMO<+ \M/A9R V(U)=XV1R$FS)XA_92+>I:?R!#T 
@X^TKT$-_;:K($]G" $6BT^1^I_X@.#_,S)JF-$_YV_  
@=P ^60$5*$DPAQF598PA"2S.9310?RH%&U,#H/I/'@L 
@'4.$FPYO@H,>^XSQ_WMI'D=_?\_6!Y8#O^%8^AA(KP$ 
@R49@Y9S5UFXE.-XNM1EV&]_LQ3Z@%<V#[TMO'ZPW<"H 
@3_K\[]AP[*T@> CP1ZM%=>0_I'UWR8E=*+KSH-56(OX 
@VC&QG"5,1HLT0#VZM38^KI]%5D8:Y*5^+B*[AZ[)%!D 
@K6G:0=\4O>*Y&?%OR&\DQJ4$&D(S'QI?"NX%B;IM=ZD 
@Y?LGSL@@BTT&\PH8B=Z?@Q$R-44^K\C&0/%P$FXR(>0 
@59W]ECP[=6KB2#UQ:7;-8\RWU<$1H3<AVA%WJU+Q97< 
@Y&%\^7;UTX4DLHXXLW#W%%"ZMOU@#VG<D-,98&I6 $, 
@CFT&=L?0!3"<(WNMAKRC6X9V(4C+2?&Q98NW6Q$)_)P 
@G"6:,[S#_ HZ$F*1!%6W)HP<$=<ML*W/8K4?@\J+XIT 
@?&][0L1-?I4RB2L"3J*"9T-N(8,X4:575% &M<Q$K*8 
@),> \"L+I ,.>O7A3B9B[\'K:+#3B68K4/O&9MA]K H 
@-%#SJS\(%M:\._Z:* (+\&R[SF2Z\Q%:-I_^&8^,'08 
@'^AS NZBA#(ZC7]:G Z58:@AH2"W2:NO?/:>GXU[Q"H 
@O)=9P__E2B)F-H$X18K+2$\1=D4&JO:H8D9#TIA[XV0 
@T?27O0%'/BA3+]=U']!Y0U_9L#8-Q./4-M>U>,T #ID 
@-''A6Q$H4  U%_9A4G[=M-,GO!1(S#KA5;8^-[_[CF, 
@#/@FLJXD=^JKSU1=U-IQH<(MZL?+=-VLQ,FV2SCV-QX 
@L13S#;'0VA5;:#)GQC1[\"AT"GT;"55SO"13]?+PD@@ 
@EZB-!**K03S;^VE#V73."<KFLQ2>#\%N0E62WW^F1D4 
@<F;QSJ[$6 =A\4, Q !%Y$3E$U-9*)?^@^S-;CC&794 
@0L5\_'PZ8'^YKC#6BJG]!JYZ"(R*3<;T*<Q_(]J#%(H 
@.T<W<CI0)O&L<6GX/O0-_3VO(BU+FCV#<8P0""04<=\ 
@AB&@,6\@QF/YVCU_8 \PM?;UJQD%_20,KUE0'71P)00 
@"3<H*5TD'YO))V!4H!_#VL+E8-]SO\]EQ"LW2MXHO<< 
@4#JK(+'%GJV</N$UU(;62M 17AY%5'$K@OR;]U27FIX 
@;)=7YZZN[V.1!V!9YM ^W.X#9'H/6U.1H0L]+%\4:IX 
@H=;M# "0)=2\OUJ34R#>MLA"3^-AR\_K]XDQD!49>AP 
@_%/2K(EFB%P<?QSWH<RV6',?E[KB*6E UA?5+U<PFIH 
@&6][D"9=3N7S4H@^QCU4L4F"_!=TZ+UL)HR!@3QR?E, 
@Q4R6WDY^<NT^U3%:B&S6Y6UCO&SG>3-W36KEX&\%<#8 
@+=@Z,E53^305 CP7!$!%"=GX_AD'(!)JF7):3JFP6LX 
@Y]]>X;2+1U7S.-9&-(8OK<^D66>YVO#2P4<&;&3O0OD 
@#IIN!?W8:>@*S'9L!!]CTE^63R:%Z^$JW,!3S*<_@/@ 
@K.@3OKX=)$:.QK5%^R&"Y@JH(5B^G_I%>"0(7)(2+M4 
@6A,-I)I[XD+,AX4N#1IJ9^%^1C&,O"NOEM!K]/3F]BX 
@;T*<B0+O#0R%,$U;DMBK%0 ^T/^)G5A\S:]UCB/X^?P 
@\-1175>O5&"$Z-IV6BZ.D9%V^.V!?L4\V6DH0426IB8 
@07I)7TD 0201-IX/QNO@!ZISMTJH?1G,-]$$0IUDLP0 
@:UCF-U!2$Y>E<95<:+41(#"6IGA/EQX^N<I6_'&,^S( 
@+9/:NIL.I]V#X0@@-"S+L-R Z[9R;D(OCYYD8^M?W"P 
@M;SAPQI- 1?4_1(;%UX #<_$SR+;?F77>80%HEC2//\ 
@#^,:+[(<1[*9Y.<,4UOZ5.8@])YD!C)Q3(G1/MQ!E+L 
@]M #/,0F*KW7O>R?:^*2\%[7-X/ES\WUN6M[MS_.$+@ 
@S0J46+KT7$A1)_@"Y+:.J&%K)0U QB6[;L-"S8I>QB( 
@.@H?78^?WA;PQ^H:=.5W6;\P@@4OHY<X? RI54L-^J$ 
@G9G,TUOCJR0*::P(4O:PP]I_HQW<!%HIZ2-?;OKJ[&, 
@0S5D:G5&M%*>X:TVV$K%Z516+M[#)]A!G$A([$(U'/T 
@@*0C/]VF\TTH6#.2\(Y$'9!<AH'>HZ)6Y:U99_ $!WL 
@YQA7Q,5%JS_#%K>!.VJ6J@EG@P[L8"1G&4HV7UD>TS8 
@,:-)Q."0D_MV,_H?+\2&VT+I%"0SG$O2H>Z'!L))2V  
@I/!C!,6?(>SPS$!_[LSI4EB8@=''UO9MZ!//3AV"=<0 
@8^K(CO>IZSRT]=J$^L0>X<AH!A,P"/@B$@V+I6;;T#D 
@'K#!;8AOJFN^</K&./TN5B?D?X28':L8!<^BR&61EM  
@]BJ0'=1]-N=^Z^G=4/"D:/:[19B.EOLPV56$7Y(#P!H 
@8:MP^"4!=P*QK&R89K;0WT9F@)$GI/!5_=A+VY]C[%$ 
@I5:%N@#%*9FB(KGLM<0AC^U^ OI_D#9<:"JYCVF O(0 
@E FZXC!).WA#T4HYD"+=+58/_I;3_[#]B_:H*Q-&^E, 
@T, O[MVAUE(V!19/M?D^%64YC@@9+D]X6\\%G$98+<8 
@RVT>Q)FX4[ [O;9&[:BPFX#!AL]B$M"R+<P;2?9,LO< 
@,=;K8[!5!O%/_4(;+;&TI2OA(G7_Q0J1,YN1*VBO0!X 
@?H3*N&3&(VAF7//OJ  N0VPG0J2Y&!UU&"%H]QO0^>4 
@XYN6Z>)#U"$7Q.33-FL\Q;%2M6TM:YG5**R^13B%VWX 
@RS8ICUP"G?%)N=-;9R7I#3D:0@$20D6JSN@?!MX2_W< 
@PPQAX#E,_O:+'E?YA[L=41!S;0+YPR4&:*V24R"SX^D 
@@;>&,?!7W9TV5DABC\3GDZ/\: W4L*"C^AZ4@'(684  
@V^S+SS!MS5&&=Y851(B&[EAN\1C' Y][Y?;HP+"$<PH 
@PFP>LRM@GMM[ZXJ+%09"XHT]VCET]% 8B1B=L,:'PJT 
@C!66C\&V)&JGJR"(=&\?'^<:& .I-%0FO P,[IG#"-X 
@\JDXJ_?.@0>#/;2AU-2M6Y/#8XT^2B/IG3EDH%!'/^@ 
@R>NY64M;,-G7>33'UTSH64#PCU<K &X5?]$YG@]$YI\ 
@*K4#OQZPIPC!+I5^C#VV!&ME%6N:-JIP#MT>KM?DO9( 
@B4;(D#G\H_< ZNB0F:6V-(RU_)IY5X\^D&+J\LNP(^T 
@O!!TR0ZQ8JW@C>IO!?1#;KR*_1!@%5V3B"",4^GUK"0 
@!]/,8NC2$D/;M>6!@-4M8"KK&QKWI]02K=3M>6A3=O@ 
@>[IXA/Y;C<@<%_FCN5@HMN]O@X&IX/8TK96>V3V\\84 
@,]QR$H5&FM;C7Q^OF&,/ DZ\F(X:G;9;&L?P<9_'U]( 
@!BPGH*MXB'I^"EW*+39_3:%O\B9S::0\<&Q81#P2U]T 
@)GZ^[%*8JCD?5P83-DN3S[D4@:[9B)LIRI0<+-"%[U0 
@OZG/MGM".$@NI\C66504:P-)G,.LUADH2 HTV90<I9@ 
@6;U(1UZB6S&8*DF3@L[C5EX$M@V\JI7)9N8&](>,OA< 
@Y6O(&K#5B)]O8-_:N_%O*<4+W0D*,W(;+A%*53H4U ( 
@6PKHK8:Q16Q.-_M\R&DN%&OXGC,+,J].,I/&1!QXRR\ 
@S)%+]NY;PA9VO6Q7ZLX&SQBKL71E1-\2)9^X!#2W*C< 
@&<RBI/"P0TR]*-MDZ,BY"5<J;M;( AP#ZA\*Q_G.(F\ 
@ VSC:T?"'_94< HPS@X;I]<34>_)FNPY"QQ_SQ/%/<P 
@3$N4/]VA7=TC)K@?;E'7D_B/\&EC)6,#T+NGE;.4=04 
@ML>FS*G$YE3ZHWC?80.C,'(]\O8&M2O8SOQ.&Y>7'O  
@"> 1(Y>M(2#;14\!X22%9+N=RO_[FYB?GR(_?B.\;,T 
012???I[?S]%0JORGG<+6'0  
022KM'@^+*@_Z?,5U?VD%@0  
`pragma protect end_protected
