// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LUso/Dajm6Eq9xGQoCd+gHO71WqxdxSUElXicasVRATTh8YiteCGzs4Bsk2l/6vb
FDZgIoELrh2fSQlz/qae67oEHsya8iJTiBQ2EN2VIKOkR8HrVF9493zZK3CiPXWv
PZjtnQVUZoATdHchas30WXzgejPQeAgKJ7mHH4jlAI4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19216)
qNVfeqvG62d4+kDxuo21Pz0x5f6XEArDHjX6edI52HhylY8c4yjSB+Tp620LW5PK
Fj4GQ3HIu2owTo09O4k1X6SIEMxuoFoL4khdDZ6nNDjdeXHlxTM8uTucXLorV9/5
BEI/1do0PSPv3UXoNzR3HG2ClsHsyZUFn4csOgMJ4A4B2EknLT/5s4lt7M+UtZeB
XSSJ6ALJazT18mz/dJuZ8YUpb1Tw8Vbpy3L4kldR94RfGDm+xyWdXSe5ggDYAaWy
QMqslC0g62DZt/nSHAV9G1cMnI0fs7Hu94IUrcOUYN4p1vxhLz10zgppnoYC5U3S
0U7u4EdrNTskv2q7tCNy4jmSzvJpebFMCC468ZoGnEPFcqZt6ux2jVsqqmKcr4a/
5iOGnZ9KUGjgC/4zqcUgZsyY77iXlaF8St4MRff2udeUwgikuIUkxcr7V/0TTms7
mAeRVMgIizCOL6bBgyBWk+Bz5Jr44vMhgSb5V95fHU6AONu+/oB+2SxLm4qc6tHg
VF4fwFrkpO9x8zVWhW7rqQEe48z+KCBzqoDzAY/k9N8dkMdx+Jm1ltKJSFQwlF1C
xfuhDKK5to0bQTd1fPyHkkFw/f5l4jN9q5+Br6HK52d+fW9ZddtqX1c/o3NqqMQj
Bs7ynN3jTkddg4uWHBIF9W8fuciyjWLLsXGJV0nF4hXm7RKPkeiSHrX+CcpXTiB8
XOBCyxURSF7zHnJl9GdUBTP0YZlMpJH5wW7RBk/9QSIYYPIOhPbzKch8jjCxGgeS
pnxI7Ck4BfUIL7DMUxgFNlGX3G20DuVK0NTfcb3xFhCq6JPQxIxhBB4SUPnBRmAW
raWW6jo522rUFtXG334JbZaQ8ZCPeEV/kxria/3Ua1dhKRFt12DG+gebwIx6lQ8A
rWWB1UR5MuFdDWuFoKFs2h2fkQVEgxiUhIfJKbH/C9QrlRb3qrZzOnlgOQOy8yZo
2/HUVKBTUL9KEndd48RN/Z3gsMcskDMeMbJt3RDs2uUHrcfUyMqJVtAZzvLfMNEu
wJWUnLEcwnE/emyQ8DJmkvrk3cli67qCDA7CVyQNyfMGFhzGWKa20OTvm+1HtGHQ
S7XnDoucqNNeWO2fDgD/6ZbFz42fpvJf93lBikGJTUSseuEMsQX1rPjRuTWkZx2K
+o+1mpKSHGG+dY/zopgknTo/d9lPQCFVdp9MXzj7ntwnPfTScWCGqlGLbY37O0FP
LGOIdX1do/FJ/YMgxIRi1xueTHUYwSOIBheSZ5iBdfrsV9HE6bvheV6r/m2NiiHa
Ze1aB/9VLvkMTA/a5b4dvU30sapYx7UPqTZKAs86mWzA5mJWEX4h4agbIz7GaKL3
6vYHQ++1N7MuU7uSLPhmOSWlEnNmb2j2YJsS11INOcOzgLyip5OZr017VqixToUW
4unt7nHvmKmzqrkYhCgFvi+cV6yzd193AIorU08ZrAD+tuWZwVdPxgIgyoLGSluG
h6wFplDSBNICOrIsnkw53pFEZ4V4KUMP2tKBUv52+L8ckt0/1l2VBUcoXiMOfcpe
imCksR0lD4MA22h1CaiNeTZiKPalDUZi7uu49znIKNAB2ifHWZYsJdoM5352zGL0
5A7HO9kh4ohUV/pSr5AzkS/eJ7M9GVPaKZN6zinOot2n/ur+5YPXfG1zMQVBkG9B
trhusAHbFKWPLgFzwTSOp0Q537zb75OG1j7fr9iBobp45HRAHdwvDIPnL9m6PyWx
i27o+GlVrw85xQUlVWytSp+JS2R83Br+WbWAYhJQzWRaETvymbdJLGdepRazCp5X
g82tvT0uGXTCl21n+pLBDmzfQ0Ssq3vnSJ5foXzkBUYS7cmA+YgZnoO14HyyBnlu
/xPAHpRIR7nDmoN/mzWwy/UGcQuT/mOK9Tdzukolka84kr7OAO6SuZ5MlNKUsc/X
Q04/Cr6BmXz8GNX9/7yguvV+RPkL9wQBEh+HoNPxtOvzQIjwel6kBXJAdAejiVcN
src7hbPNe0DGd92ZOF2tINaMCMQd96n8x5yBmB5VtVjeTL3O2wtn7lgdnCLNR7g3
vRtTFRNZfHHtbdH5Kao3cvKMZq0dI/AiQ8sLYk8wLKTKmu7reyUUa8r5zg0JtoDT
ZQ7Ek1IYNylo6z4MtkmRWK9XKRd4shK02VmomA8z8wQ0shQrwpqQO9z6UcDea6UY
ZOI1HNwRT1JUgfAp75gjFTFQ7R6PQOc2UJSiaV7Sjrux4jpUEIMfsNruvAhZgqc7
ESz8G+/7s6hVQBmEFihsk86m/eF1fLngrYuds9XLFVi2jHtN50F8/CuFI8c5f+lQ
F4/qrt8V/QVjv0VO4Hry4UqW3ET6XSQVMd9VN3Vq6BFuo9vuXPpTRMWzpJT/CiCf
rMSb1RrKDbuEjXCUPKqUMqCfH2mlD047FRFHRtMNIj1TboLwxZ84ZToo0+9Vh2Vc
oMF3eU0haLb/8MIXOA1eFRWmzcGx3pE4IxZLLDnBqpS0qOMiCfaqeJVnJkgGGhG8
wg4Io4jihWx6AJNLr9gDagO49lRLLWSbgTluWRj+y3knmTf6BFKaFxjI7TNpFR7Z
HVeAouUbv7tuASpxI4fXWe8t2ZYnT+NEE+zXAX/XamEW2GFgsJuI8NX98geNwHJw
YQwu22UTFyNIQAuGVVdmt0JbTC7cE98B7Evie+LI00vX11odYZQD4pFBZdGswjC5
CKOf8rl2i5SdJGKMjhSg4wfBI+n7UJIw8HEEAj6mfB2FshLoHwqud5rcyTtabHZw
Rvu0J0eylCgBmio2igZtKI5TDNRZryb/VpfwCl4cdmZI+kCUfyohFCFBsnDIvMGA
Xsrf1ow0BCspu9q71XpKseFYLMSmL6+SF2qsIpDZL8uBQsDJUofJyT7um9svMnSn
NUnEIbu4nKSDYRunU3yZ8/VrbDZEqJss4MdcwAL2sUYe5N1F2b4Q2J4mLrZMWeN4
3dIggc0OxUve8C2scshbwL/M0PSBxWwFiYjqnAMJhRgQHEZYIvw6HQ5uENFltp9T
UQbh73teEy/kfuF7SOqNFLw1gIgnV0igO0lVZcBVWkOeZb4hlrdF39uSQEo3VKz2
dJB70r4b72Rr7T4/kFVZqTUmKL5bnyWX89UmCM83W9dVCR/hxNbVZ2MxAbV4UwJ7
zJJFbo0m05P9NjsmrAsYYMAyEsgKcX/KJVv72oUokv1g+lWb4FUxs3DKQ9UjtpD9
crCzZXqWlrxx7h/tDFieTxz2+VS++teXT10hSrO/aq+VBwQr1VO8wgiGYo2+MVUu
yvQ/ZygJSptAXn2k6BzwqzXbxgk9gAuaK9JPyS5Q60gX6/+EP+19fzl/I9RDcu71
om2LhAGhfZcHJosLbkwzZLsBSEavpPxcp6VA/bgTxfUjuika+JzSIz9t9UeMLGaF
jaZUfJ6e5na34FMAHHyIZcqeOiitDsr2pbnzuLwUGuCKCTdfh239e+7I0ItB6MG0
Q2GaZcNAhWarnWebl80yHDU8rT78YTlxR6UBqDyRDUNoScjxtCCKW4BGNMYR2NLP
2cNSdPCoLthKuSs0X68wcTVs5+4AlOksXZmrzQjTkvexuu/piZflSXn2Wl5+0QVb
HUV/HYz48xlwc8Fsg//AEhfDmDrdobPQRKY3dQq0iXz6Yt2xl3Ea5ywrAwt99I44
72T/MAmKD3MLoo2eLTM0j4yfmHBUUIv3cCG++EF+jy7HNxYalGQz1tbekyEx9Tbx
dDcNwDYwschZkWmgaQ8FYeVuWdeMf10LTMnoK6iu1kgqRmOXEjygdACg7uq0si/c
eo+XVXGz9FCufe3KBCLRDI0k37zFOQ7oTosKJkfNiU1xtA6uz8hG+7cOj35r4G10
m97xFwrmg8V0CsbtgYUZEARGzwNscV+nfUX0O4m6AtSaJAQz/ghBIawN+6RCi8Kf
vqdie2bsinn1KvnvwF2Tm1fuxaU9oUeaAxON3br9M8lyDqrofeipJ7fq5ULSSh6z
Fyj0cXnVJt6mnEq07pj5AjgIk248dYRVJlwV/E69DIuHgyez/v+QqmNeBEiNem02
Xfg3C+GUPm6uQXxdu3EOYSyNIGmwrNtI6y3Wv0PxnvxH4bWHdQm1fOPE87QiZKXl
hiyOUBhuDJZok6nB0tNT1h9AkHevsaRjinn3hDxShsXGHxLbt0IDDp5KttBrfvxx
SdFVzr8bu7D3LewghbwfEamo/uvCaRRBs+UMXJbx0zDpaueY/IQk4dXuESFdL4TS
qRFqQV6TbremR3VbTAXs9z1V7lQ2LgAXpC4zT68QnZR0gx7BX3pH/WNtU3rgzSQ5
fY0EM/r3g5opYxwpEikyOxdfROap/6Km0KkUWrFzAEvvMJchIIUSqz99XAdonEra
Gatggv2D/cBTHM8hoEbJXtAlNVYReJPWhOg/zjjENRhdOp7n4sy5u+5buAmZOEOB
l5SfSqGRTG1JRqdDZzCe9soBoVkFdjK33hW7MbXV2dzlP5z0O950rYHUYGGAPVNq
pgfvtXVtgQHUqmFvRWMBTIQ9CAQmfLqnr+sc9nhhrBN4R4BgV4WK1ScjkYrVSy2I
793x3YlVr2Vxq/eO69EvBQTykFcSNNYI1/1/EynhPdiSmxpg3HWPSy++TKxddW6M
0j5RMKKzUmgCdFskS7BJ5kXcpqoYQM+MvRE9ocQxT7qIi1iy3b7zNzWr6bfpFGC5
hpjwFLocZj9u1UMsZE1+RDugpKpe9eftmwg59cVVFPWcsvYfFfmdzeOZyqJijg9X
MXOdNzt5l3w9pJzQNRhAFdAH1jE1Sa4QNAQufHUQOsldOZfVJtJXdl7aW3RVfDjV
ipHrTgr4e/oFgeUmyItWAEKF/oEWBsg1E544iiLiHkRX6KvP5KmM/sMjuIJ3vClQ
jkSwCPSqBQGruX868aTujnx97Fobe2meFigt4+W4lpXgPlKUOYpY+R/60veCOGJc
oLPzf3Xmp6o0LxIRQlpaZwF7g3su55AsJlwcP43DMn2aA/Q7gIo0aYvF5O/SkCkk
Yw0jFHV1fKVolobaKb+hbQh0yQG+N+MBHku5IhtLiwbm0B4lzCpedta1sug8fVvE
0aDyzerLOjNNqyhySQuWmFq9uBk4vYlZ0ZYlj5JIE6RBcOi6z0FTIvef2GayaVgw
Hw21sBP46s6oAkR0dbGIneXZ5Awwv/HDbOOsnyoJEbzcYN77Y/CwbhhiAL6bc4HZ
e0iQdtcMqarmwpSQ7EAX2/IeiFw96sDREiLBsM4vIgCwfYUXm0aPi/0JIWHboQm8
QCl2UIN7250Gh/k9UoDfQZIZeTBJIO5/H05n8bHwu968DNNtftMZAsyGKxN99+kT
xJB0C1avPgnk4yTe0rODH+XnG0IG86DtRncUJKj2/jh+RK088xQ1ICmtjSLYUznC
WYE2292UgSiXOz9Dp/06jpiySDGsTcwX/bQhLqPhYYZ+GiTwWd9LDET/mkZxWgpN
iVQX4EgPGxTYwsx3YB5Lg909B+X6A0ZQnjQkHUgc8qX4fPM//SGQFLfIokiPfS4Q
qseXyTGz5URWV1FB0BVH70vCd3bkXR51+a0ff64wddYca+1d7G67SZHAemU62M2e
RA6fBk9HD7Q6V97dgkx9tmrPYJDG4g8pK2NfXACY908YXpkgdrqBJmGJuhnmIPoP
/QVsTTxzxKglMh6Cew3ANF9g8ipQbQphewhJiOeBTd5izwCMlZWB41U/sxIWp919
ybztlw+A66wjUuP7+QaKmJ5SpgWIxdZIDSILqrbqbEwIYBvQOKU74RwG2aYnSpIV
IZ1PPunJYDjWV5Dpct8bqp7gIr8iR2D5Zf2ng3SKbOgIJBETs9F8+FD6CpCt6vSC
HWa5cg4VTYVp8Q5B1ZYXdeXJal2vVKWwZrS+KOdQjSKlYoGSvavMuogBIjTfDqou
C0qZme7aLv8RXfch7fPoPQianNMKRUSow72a5qRXoeqZ1myENjo9CLgOYX1ypV2r
PQMvUG+OJltMroq5vMdmMlhycYmVDFov6ETMgdtZOnnoTVI65woFb4KJqJf0nlnx
oDHxYI6f77pt5vWPolSdDMmMGz1IqOxg+tWjAfp8frOykNpQOC2JfhwVtsYdCZGJ
eOVqGpccMqinXbibTIUsU2QVGdp4G3HfETQX3pBvOs/dp9JC3BcAt72FxEn0ABso
wx2rBU5MbHoNMiJIzocacEkX7jffM2K1hUqb97U0jwDfl7wLRK9xoODvzZTtHeir
3ikYcolou1BSws7woHjnZLHZiyVQdRYkqm9AUwNgrlvepU2aPu7jPrLOnAIPrhLl
yZcq3ow2SNYteY4lE6OYKy/IK9KmrKygVyh7HRtuE2e5v7K5ko9L/SyJYMxLHKKy
90VE7rE/KVqT15pb4miYBzFL6TUjRT1cQzEa0u8SCaEYH0mOqEyCvdZ72s+mFcx+
3QyGsNA7a12bl3x88PKxBktzxsSsJ3ddIbl82UInOICkU7uVy6lRbPlOk2iFw78C
JtApJY+WK3God1FucJF2nhotnt7UQrIfBUc/O7jvFV7zv3/sJkHwbpERVpCpe5m+
88Al75YeEyTr3sAta6lTIfr9hrY29mOYsKFxgRIzq2qgXuq0FRQ5AigxNkdj7wHu
m7ej9WHVjd+cWQN5XvuImMcJboxKJUGsxIDI5BBi/BwfhN4nd4Nkf7YLlNYdMJ74
WCfXKM/VTOrCEOgLIva7qfosq1WRX8b1lkY9AIspPGWBIkRSNfW46AloWaL43dwc
3lbJSjxpPHkvMS9v3fAq0ygCHMohDuUQZsDQU2K4FKyKExrJaUdDBT+UHVNrp+9t
Ca6M04ehgRUeKEcZed8Ab4itjTdF2w+MQCVP6qnf15MmbdPct1aWY/Twq3elniuu
aCvAQjoEe2XgKfIQSTyKkblMt4FPYU3llccIrB7mHf29T4wtysUdnTObKaEDmMTY
T2unhIxTUwegDsmuyb7UIdCO7+UmZSLXl5D8kswCb/yZU4hUucgvMt7025Z2Z8Nu
qPEw4fKPFE97JCkgi1cRdIkHJU7aYpOOEdlTyGxC5+phuTVAUJ/DNQEStHAxokM6
neynfC/eHUgF8JL1p6p0a2dgnlwkuW0/7G2SUivploro5iu/Fpyn8fyjxP2CHphd
kF39JLoTSZ60hD5wjjm/OXSWZAV3kZZ7FkVKezHFJWPsSVP3gUCYmzi5Bkyov3RT
FaLeyaMhjj9n5cqFedmXPhrtmPaFJkA42wvstsochoOv/mvnj/lQxWZ0787/fPVc
nHd/G3O27Omt4bEuPmrsrU3FSC0wd95/ncZPQqMaJQh6sQIUuJkoOjUN0MdTmLV2
x2MPROiq0rKpbYgMSm3vqXL/cQJOod/lPxoPIS2ADwoLsePfDX9TJdMyH5tJxGXS
SSdo76I8vMpVEwWu4I0rsx0qzSwi3nlOmO/SDkUdXRMVgu6r3Dt0NQesc5Tg+4At
fhIhiUKTMWlJALHllo1p7Y8SiWRuYjZ70gIPDF5HuFVflGTaVY1q0PirQXi2HWKt
+nOJiww60aJV/cg8K6A2gadRCfjxMadIaeubok2RUAUpymLXD/gjtvnyXltJmkxn
Dk4gG2hVsrhq6M+UMJmUq4ng7IE7Tqh/VxvczSaQRJrmsdnCSbctmg48fUdG/Ue9
5vFxVQZLFjbVKnLi/ZlRrD+Yq+bTLQF0DlDM9Bqtiu+UDrs2IBIBEZb6Iowz8KbW
ssIDR3HD/GyPOliUyZKf8WXcd9Yx4pDYXqBP4LCSLCJaFLs3QDPHYyPa7DnEAamf
6zjjCHFl7VClpjKHv2wJbUeiGcwadAEFOtaFLw1gxcvKw6lITxggoY1hAp+gQZZq
cPK7W10NO/1EtZDi7rT0E7hR+n4k4oOWcfohF/WdxTlfdGoTxXInAfNaQoQteaJy
6c+AnhWxojeII7tnr1md88zHfrLnkA1qkKmoVLDr9KFcklGGLqTqB14CrOlqqbDe
TyO8THgvWQhiPLcP55OeCWHPUZNk3oz+y/wtNbDAfkGfDKGw7JnT7otdPqJZYXAL
xxxgykmkndDjesTgvGEW5BHHlyEbesvKMoAGXK7toW487ZLbizgvtK1p/nS6Xlas
RrNi86ELH0YWU2dSvs5TBccYQF0sdZ194+n0GEI7fSmt1PRFaoLP2WMG4+Jo0Ddx
JE/+qvFLapc+XHmos0hE4sq6PbljvWxAu4IyIND51+PF+zsczObUAgPwFD1XCZup
HrGLe801l2hiBQ4j9WcAGJeRoORsEEa5AxwP8bpAjIFlnBfITfyvb0WxOPB9ARuD
WxEeyK7wfSVyrVRKH8l4ca8Y6SdGaSGwJtn3qDti+wJgrjSkEd5ufoI1tRFrBpz8
sscVqkNvN2REQ9smluqsL6hZur2SSzuxv2dEKjcagSyACOvUBNWfOtD6AV16cMCM
pJ1oEcWJzQ5BGeiXTR3wF8RvKuM5JRItk9MiZdnn6iFOW9QBI+rRyphjS/B7ii7s
fmiXzVvOXUag9VIrYkpd0RKwvlf/xKWVdn3Vv0QTw8N5y/OJssrp3d66dpatA1S9
coAREYNgl0Zm8LJA5oSlWExrtN+1VlyPzICccP4miPN5RxSLXk75IIc9SWqRkhyX
PvSljFosKLzyG0nkOEE2DXY7w99OOjbrqwjb45RaXNnO18hrzNeDoKVwTaRTa5CS
WXyFcojGLJYN0XcIJGrD1T05F/I003tTziX2W7PShW8zgGo0KJzKVlxz6HEtS7Qb
BQGcCRI0Zbm/HuTftuGG7dzyYgwIIbSoX1fHUa/o7KW3UtIJu6QLyB/6sjNQAo4M
X2WvtBdjqkWcn8XW9KXGJXQd9GhMeoXhkuYEcKZdPiv1NP2C1WYa016C8nuXLILE
oZAUoL6YsiV8trTZzXbfs2hRzHb5hE3yDwGadG3mmCOy0GW3B6YwcYI5ERnKfm5r
Nx9tRdlywtZ4fKDfP/opVH06ygnP8/owpOi45x4sr/7nZYmc2elaqHAatArnOxae
S561e1ZctYn4lAYA1CxkvPNYKkYx/7E9Z9GYJ5IEKmJatjapXdTFqJtp4myBvBQC
hSw8ZsO/ci0GmXfjYCwVZVse3odtYCeEd8tGwMexajT8G9ur7L/n7+08HMVJUZZe
hcRw6bCfceP4Nz354cYh73CSm/yJ6eA0gUWXsl2rZ353vv/4edal+NpWfpsk4ft3
SVxTOZ1Pg5CHf545rjYTZydtYFiCNzPLyKZOgR0HIGgt/7uTtsZ21ER7DI4RX6PY
p0xFdif2aMC7/Fg3kTdGmzWWYMUhutDXxL9ZZ4FNM1vSMg5cHmH51hITdJZMCRvK
UqP9Uau3zhLpzpSpqjCdlr68MHo4js8j7ZygERoPwFntJVFI3itStyGJrei9fnyY
UxTiS89f4rg0bc3/FJ2e3dkngx40TnowEQtXN++JYdd8ulSKsGKIwkwiaKSUPzC+
BwHNYXekPa8OcVn+fD4Wit9Ukjywjb5Icgq/06Il+X9LOj0dOmaevOOlCdT0k1ET
PsnNZ4yH5Sdt//IoKiHH9wFGANk+6nBP7F+n+XRBkQl60XFnd9hESEio736nJZfl
xt3rLAHMXTVm7buZoT+ohwjSruxPyOx46FFefSV6EntuD+qrNi5Bn/FT1ORNvcz2
eUzQcyceBipSm0Zj3uCUciErrjx0tUWW4+iKvM++PzDg7uacgHt1PxAHpPHeGMjg
zEYXOFSknt0dkWO1eO3Is71njz/KsnrHKvpkQDHQ48YaonbieS43XgkLAlZA9fse
jJBLvqOZC7qSq5e1gfEER7X7N7ZxHC0gWwTMsktD6oAuYqe4oAbmqOL1Vg8dsqCh
p0Dhl5tK2Cvw6arFQ0IqjNDn705GloyXkfkY2TS8T8w7S8xFbywODIx6pWWb6ZQ/
IQEAtcBqAJhYrbWYizHEjR3MwFLvmXQlmeKLZJtWiiCZ454NaFAmbHW7SGEoooOi
LS7iNIDwaWWfXMuJS5M0vdiyzbjjKrb3O4c2FmoW6+7J1+Rqg+D4icNnhzkqEeaC
lG9wx+AG60+rlsXeLNusx4fxk1Eb0g9VEDhDbJ7oR+Lj1hYBYvNBvWQHMbnnkF0G
Yt1d6PTSURkXheNMITMie4bjsOitLCfeMzMkyMLjArQdaEBb5OXSSJIX7iNc1F6L
TIC6+KR8yGRHIFxXZvCu0Re8bx6swdmPYLbiYG0kcL5PILFtS4YRq8wFML3z+qEG
5byHYtyMqA3DDp9cSUGpNPa+xn4qSB0AFmgrt7vDBf5mBXAoKTin/RPEfmDJIAO0
EbAOixNIiK2bHsuVzLzwewu5Mm7/dQs8N0B6QjDmaOZDqXQeLe75GxmjyyBhHiYm
ZdnHRGvCWTjqstxzRZmgC+9yJ6g7UX8QtsN2jnGGEHG7UHZB81c+vtii9x+C93SE
J8aBGN62K9N/pk12AYvBHvYdOI3Eb0tzNrYx+n9NlDCnu9NkH7QHrrojkTgMiFVO
U4CUgZONhfjjBNW7pLrw2wiyZ0x2IebMEF6H2se6Cfvsb9cag87LrkiFnqlewOYb
gIToSMIjbT9mIei+dkMY4FpuEPoxOxsUotwXCZhvnwktNEsCHeCFwzLgV2jNntgj
LHwuukQKTKdDOMtRo+JkPRfCNBxbldl4duqRhkSV9bDD7Rm6BkoazuXZM+URDVWC
Miw751lX/07HTgfqyN3GSaYy8+UqXwJgwU6oP3ER2RtJONYfGD5MZd8Rhy/wAIBo
GwLfyg0prR2JACvUf7GK15hpwTEiRIxZXvmjv6Cu199DrWvzc+vFbyLpkGQdicxD
icMz6t62lzg4IqCBTYSrYB78/p1DNKWp1gCM99bR6I9JeGdOyL4gE6XIlgjrTzW9
C5M9tioUAoUVz7BYiSE638LvS52KtqtHozH1V16njuJpHS+o2NE/eDO7REzx2c+T
MtYFM5NV7A0Lm8etx2YuuoQXpMGF17GpoOst3WLfd4K1P1Hi2/Z1zAnzuYJLYgA0
a/58vYLu+mPpK9Ef8/BqhVIxF1raFwbS1hVzfFpar0oPZ1uuYtX5PZ0HgvY2OwEf
t7QG+8q4/6oDx/GfL10mX/FMBIhfe8mvnxmBYUadl2vdTsgobuPLjjVcH0iHFLYS
3/2i0La0vLfRAPswwojSvfiM2sBOPhahRkXQ3eRsV2QtVNPpS7Y2Rd+DmjLJsK+s
ub9zxc4neknRAQKbmTYugV7JePgB6oDYIiu7DP5ZcWeJXJFPXWZEPnUJ5kKZIn67
WvHBrDDh+STcCDFKNuohz73yH7m6DuTS0A7wvXSH9GOFdwrErBmmZYti//UmoaI3
AcTtnTT0/MLGXr+p3673sIhYrAAZh5kFA6UmOZqsRGhUoDu8wHFekiNynUMoUPVa
9MgqXCJPLUyIRlMvEtGRBaWnkqemHYTFWGW8lxT93sufNRrSCZgAf5gUMfGrWyhV
fUwQNGK6ko8BB9MzSpg7ocB+FruH5KdxfVja32x6ALYPleT8DMIzblAmKX/CrueT
XTrr5nxp9KQ4jQYA/80w+NT0cN/Y8otxJJrB0S7/DFdIyxXv59TP2d1M6X3kTQra
T98U+6S/ORxs24OfrocAg6QTnLdlKGLar4FF2YySaZnbu6fYW9qqKbseLTMLBGbH
mJM9IVneRHm2RDpkuw31bkcuEH+PcfCKNZbn3u80TK4TnP8oKARLpTEczZqFK3pP
+usiJtMKq3Mh57RnKh4oA0Rxl8DVvs0WZzA939XIdNRfRSYYz7LPQJymYBra0fFI
GnYOmD+tholqulCbhxZLcf46VU36DMRnGqAEvGcJuTgVqaA5qaRndgmCFSiFQ6Y9
fC1aqWJZK8yY3W1GYQ5up1IiEg2orVbYMpiDEHa2f/Bkj+8ASlPbZt4XRtLLusDq
1H4D89CAG6ScUYWKHq6l1vaAkH1xHyu1GaL4dMMKsSGjYQ9yKpWoHhKGd2+oA6CX
tJ/TbnNBAxdzYsHofpLAkUq3lhML+V5EmwUAdojqhBp1MIlrocSoVnyLW1H8Guvq
ry84Opsc2hiy618ksNklZPyHDkfYK1dab2VwOccmlrQbclAUQQvktK9YFKXIgJlO
DgItdh6GenekLfUWPVoCnzzkiy5h7SJnSoQn/TzOFZi+4rEFrfcgk0M9I0GSIZo8
ZdPBE/dOLIqgqafcjzJE97Qgp3tiRVS+4kw1bQkiKkW4MJX4RjaGyoKPCR+ZCcq9
sEjK5eKgRFUD7zJcFf5iBuwUNRHFoD0c49QyUwSM1Z8T7opEuJayMRTxfSDlVjAh
4f8IOYwhAQmnt4l/2xlfBJaTG8uQ3H5MUq/23FjyZ3NiEGmA2JDyDTEVL5qM9RyN
nGcnnL7Q6EEWLhdrXxIY78Bo1ggkv2z6zgavLGrEn/t3YBaJz7U05F3/MJBit2u+
Ytu0XFMjipfNk/vV9kg++rRCzLrQ0d/LC5fYjP+AvsLKm5PhTWzApLNE9QqUR3KL
gUfHC2zDKZIe3pdMAA8a9DQDBIFvvoy0Hz4c93dyEDZbTOAvLjuhOdyUzbWRZS71
YzAflBZ63wpphXh9d2VGk36uRk9xzmYo48wyKuhpAgfn4WPKtj7dzZR2B/jdduLE
HYcycGEtzKqItuCvoaKuPX0Q/mqV6JLWFNthEIs31cT0tVVHNN3BaoCWhorbK4XA
fDQ52q08gaehsyojYXFjc5mtN6dqzxk9oQGKtHmTTF+nvHY3N5yRQJeO5dGcdXO2
jKmGenN9SjZwXfZ+GcBe9xfZ+w0wZC5i/gIjTU+mDZu0mwvZ30f7HBqYXShzSB+y
x+fO03A8SwviJDbWapRdmsrWdC2c2u5Su4+S1m3dEERKw/EOeXsfaygE4psO9mAC
RblCU5suTBZqQur3fdio3HGry3s4qZFqUz5I7vIEnlbXyrOa/v+FFcQ4oLL5Gmgs
qeooaxFTnvaT7j6rYNnzcdGQ3l8qh1whmF+RbkWV26SlBk8Mi6bwz+8NDz32BTHO
uNcXZmuXmsHW1OSkMwUN9S04KKf6gBARnr9JpjX7JsSDxiBWe5o4ZelzWqW78smN
HwhA82FR4IQLt1T7fF9e+Cq9N13tvJ5pLVQM+ImVoXDoy5P1vaEv92UQvGfjG7yB
oYXwp7c6P5Onsa4bqRS8qxeFLsf8ds+0+ouTvrIhXCSPLx70cGGN54+XqJwNQvIA
4a3SDt1zRYE8jGH//gckL9Ix54l0MoJssDirzAp1y/+MF0to7GQ36mQPJ5GWuCXr
OiWr6d9UwMvGiv6lsTOlUuxiOYZt2nN69wgdZzh3ghxyb6FZgoRrT9Fb+UKHH6Br
d/5GJBNfzj0zAdvGisBSYZReBepQf2IqH333BouC5iW+okMVRuOFRJNdwjtgIE1S
GCSNxEcrOKnMGkWn86SFxOdEUvGTQ5JCQtjbJuRqIq7RbJxW6bNTQOyxgMd2yOsZ
QE337SyBCoVARTZ1VGGgDyntEXKa3/BH9vlx2SwJSnqtz8TfYBDgH0+sYkhT5IFU
eIhPctPaNVxHnh1EFCuchWekbmy8+6MHQr9EcTZ6RiH3rnoc/01dypQZPaQhjTHr
hlakE6tiSpGi27sF/fvhYrNdB0iOm3+drnQ+3E7nvMTapjAdXiFd0BKWV0kTUCmB
fpI5AHlhgQzhoAOJe1V5jlgBbUl9ojqMdljJjOQNwFKlqIZg0RQ4Buz080iE6PdF
1Co0FLtvMg4BMjRz/Bcev9sE9s6A2m55QGeXwaomAvFUKVctdS9fN782u8qU92Q7
RzcfZ+NixmE1Jmq/0NgGo+11l9MaFfBtsZxTRaOfPCOnapjIzG2vNoAICqDs2XQB
OwBcER2lgXYMpy8t/Ao8PKsYTOem91RLcoqRSLxorHZsVQJtZh591bml2Cwk698f
XZF2rA7zfXVqO0wKYN3btbD3Jab78UYEK6I3SazOC6x0jFeyXeDhoiWG97dUDrOd
r9bHWKfLt33zX7xjRis2VLYtvzbkgRhS0iThyGfdDJDONKTuAY4NCAwS9xQRppI/
t/SdNfjcSJ1CLrFuMfG03ldgMccop28NYI7NG09KmhVocL4ChthTfQl1Jfb4zek/
Idk1XoBEX8oOnIybBuxjlQWte7/FFEePPICswB609lnAPzURLgg/TbrbsTDHHMz9
QADQk71xzJwbCQ4FdDrEnC/geBtGvmP2t2rZo3RLHM04kNY/bkPVqXBuY4EGGeyV
LEXV2PuGXx2azn2Cy1eSwP95QIP4gsiHF3pk/zZU4lf8w69E6Aj6FnzCMgeErqMm
6DF6KDhxL8cwiRalz5pti5Jv3oFYsEW5Cy+Rzlff6cp2Bls2meoEhunf0w33uwub
Yyjmbl2BPgkMMVHtNqPy0depZVmaaJSISyrMf5XorEyxqGdCF2EFJjQKk26Pj4Ln
tPR66ws/VBzBW8f6SaixfundwTfi67ZoUA0HNduPRXMqwn6Xn32qrvA3Dl8+qB27
quZuj5/oxJP7BkxJ1MxBNLZM9vKaoGwg++DHmEXr5hc5pAEho3OunxBDqCeIJTQq
UjIsydT+9AxEzQa+B4WEMex65dkqTXVjgzSOudSw2DAbfgYlzKY9snWA/d4QwCMu
Ldg4JS22Gf0pSg+5l6kA9PLhFCZgpylZOPe/m2Oy+pv33LwOt8fk60xZk8XtPHLw
1qWrJORZG0VCBIfSFz5umsGitqUlBxUY1EgDP/Wg5xjcQH3SUe7FHwZoXSNWNgOT
xn/u7LkK0BOop7uOBTrSf3Zu3c21snvEK2rStbwlvX9Ao7jJK4TAOmW3d4v0mdir
ZJWzGljSqWNWdgbZ+o1nEtSNYBR+fGjwqXdU0lSEmyfjPEVBoGWIL6QTTJaigI8a
VLaZA/Qt09eQnTlp+qJdYxUewzFa1nIndWATcHXr+hYmgHrkrgR5pjJL2BYtDqDj
jdfuIJEI+H5CGYygFgLxaO4DY7SFJ6gCyUXTva7MfuPVCLRWW/hlMQh7NavdYRGl
nPXxxzg20U/tu+mVmKAePj15LQ/7lrmu3neZy4kqDuoh2b7fOm2qvYq1gGs+y2g7
wFb8MJJn67deDt23vQ8NekQ+fo3lAXIDDUYAc0sgdoBupMNcGa4ul2ge32joYDdu
TboG8QU+VkjOenaXiNmKq4VrCpDuyIUqwTFAgzZ1Oi6XQ44erc5ssk4Q9ZXfkMO+
JVbdCxrHSfo3vlJH+JGHy77blNK3BGjdyazwqlAw/RQIrS+GKxthLZUiE/iGBdl3
YlFqKx4+SleZUnjxykBtY8Kc1xzvjyZbcjR0bb3PBnyNMlL3LH8vIYMrbeCRKUGh
49IeLz7x+MzFsEpJvsPRwX3kXmzb248/oNrd2S93i6hneMEkz1xU76uPNKAeixd2
+EnZadkrRtXD2YweQqhV7Cax90PchgJKdg/xw30nT8ZmlP1p1Q9AL3XcKJGlsBgi
+SORnSGtt2+okkpIaRQ8OKFOOMVZ5gaRE/yOB+qw5m54W+jdeXTBR08rrZfKedtM
2HH29+XkhyQAPBf+wyxCnmIq7qk2unWjEwyKX3O0kHP1pLuek+QnKUlR9zsrPALy
7Z3w8bIWzl1ELzzXcTFtdLUlV5YDaaBtpCQQHKlsoqZAxI771qxZLfZBrXcShahD
6g9NiXF7HbSN/ygfYOBXSJFAZwfPEuROnyd7lKpkRvDuEo/MweMxIqNOuiMjLwVD
vGN1XvHhiCyuGxTR7vBqOIfQcoBTnTdc2hpWH1G/pTRnrRUFe8AVkdAdHVRYsH6V
zbIiTOgxLBfSRIum3yfcSIzzl6Pz8YCT4jeurzKWHKJbtqUDf8VbjySPjG1cAhUS
fO3fWKGR3+R+LQwfO4wjSO9bFyS2GRMltrLoDT3vzaVQ27X79VfPAzLWbS2f7O3u
ij2VhKrdUp4KHv7iZe8Mfc2Bx3nRrSQa4P5ZjOVf1gV/kgZ2trn9M7QDB+UBhVZA
MNC/ljTJIwzpR3mU7DvMHDSvOPhRSAwOoVr9ZM9uaNAYx25iYXFrVGTh6+GN+ekv
wJvPmo3hJrFhRsNDB7+qPKFY8AezyGf9420QQuklfQq4yf52JeHtReNwffTRUFDb
FI+IFtXiIsp0YLUUPyNEIesl5wJLbqlXNBMKkjOvHFl+PBospbcrTM3zoSfl9tXP
/Bqwds+unSmsbEA2p2xDt8JtOdBEH/qgXBdWItPa838ydgCcISSXLkmJp8Ua2CRC
6z2jtbjeT8L1M90GbHIOI+9WDh54eCpgUoKVAZzfZl6nvteBq1PX10rAeue6vk0G
i66acwfFWZmkHMZYTfbFjxJZLrJqnyLFE8e9RpRki1u8U1otF6Qzb/ZmigysyMiu
gIZ/zGz53hs/D81vc9BhV5iqSzbyDSLvrsjTf8ziOWC/JSQWXf3btmKTcpLstNgl
TCC+x85ww0A7GR6DI1N2K2igkqZ10lA8+0zpyNkG2umkfrFYfvPcQTCRMKDKb1m2
Cj8nw547x66SU/t/lz7pL9FNLVAk/22sNH/+gZ2vbGlzC+6vQW36gzR2qvUM3AYy
8x41GMnVZyN2nGER8colHhTBnPuAqH5fqg6kqBVhqMLzX1XW7UoPBeTQIYfeCM9l
D/8oEbhtlOIfL+8BS0yI1FfY1oQxuzoZ6Z3wV9Bqs1iSxx1w0VcbWXdiY/gLuF5u
Ol0fIHXGmfB5Svk6iPToOT+2r2XDjYNXYJAIHYIJUpXhxNMsts2aNakS6OQF8wkK
xPyN992AmrazXs/6DaO+IWQ+vrZ7yiI5cpVl7PGlDyXj9AF243q4k+i06j7ro8Fu
JGAKuKU7FsUPmuHBlkuzO7KIDf5uHwoZhFcryRoY332KGV0qiFl7kHYYX4ZynsiF
6fGje1fQzLNqYxD4EKizCzHuZZ//sI7HR3XJCr0ZCkmMtIqjNCEfEB3nnmfkmfpJ
US8jqdQGLv7YOg9BQSVhuSYF8nz2a9CtkAIYbjOqb+tm8Dqmw3oyccLD8H8WS1ri
ZUhgzBYqFPnUlYlbUiKbA4xwJ7XWIoYRwD+rWkSJtdXk95bzkpkGnxhNUx2NWLxR
ixdXkXzB8b6p+/3G0DFA/zcY0LCy5fl+J+puehEvVbuCigTjsP0508wNn6hIYtfz
38gt6xoLJXMsZTPL9WWKjhneWv4YNObwFxtafBSBzXQt2RsyEoDs4ZDNqCF7od2O
G3c0Frw4ml0aaClSVXgSq0XsRq7SpvoG8NNSwYeVgpr9MtexgNBZElZPlLikfelQ
/KUVmQHmTTjPa4t/pOmVEc6Hrbf6QdcPUqi8AdIJeu/N585PmFqaIuHFfkhWKs00
q1Lcw1n+HjDIEqmt15xbqwfIlp8gUc1VS1QR8a+q3nMgZnbWsCQr/zeNIT8PrmD8
ykamx4kfhc8UMX8A3C4MnNofqlaHjHm/DgYhAdQkW+u2nJKDAnKqFTLmZvNuVA/D
3JI6/ZUuYzrdaGWZr4REJGJ2UpE9mZ9irCaoC5S9MvTG/aYxIJKxvJd1+zOsqcwt
Q0tg6H/vUs96vjaCCtlXMNqMRd6A752/5FzMbwwl5qwb2T/HpbW8AjowEJ+6zAeF
8+ukZu0QXGvvn141mlaieYk9Kdc8JEMUZNAq1aQZHA57SeSeDsc45lz2TxCAfP6u
zkt+mb8g0FIKWLBTXbQ6Vlqjih3ymFJdYNRvXyeCC4R0aIGegg1MoAG9l5rbbUtH
NLksWaRg1zhdGknCOcJM+BljHoswBYjRcTzGY8RSXSiLAdhoDS6VaDYxZNaj/qnA
IExJz7y/AnrAx5Bby6+QFfCyrytvRAN1gYynb/G/cGvQrAWT1o6EfWjmxEnFR/GS
cGACD4eBvvhcd43anyNpks3ns42p3nI+kfJ3lLNeybLQE2CpyWYY/Dqqz8aHKw0D
M4+S2QHXe2bzBJI640xue3WOmo7VeCa0bIM18BdzJVRLJH5lDKneEvlM0nYlYU3L
Gj6HtrZIbh4yev76mCNEC1nWvAULbYZM8RGa8sRDnMcRkA9Mc14NjK6CUfqNm8vO
qp9+Smqs2h1fqJ8aiVaN/XT17iZs/4iaKtvlRIeHwZ4OsiM5lJeDLPG3+2qcS0pc
I0skXUKlg0Q9XajtZikgah3bJnhOcppF05LFX3ZDB657Px/gbQ+n3mmpplrra5Q9
Qi4Rg5aSMa3OAwZqjlBvVG19CD+zIjZkp3jMXDKkxzYFQxlXBwFkeCRz+xi4oZJA
LDQENRO6oX5c44E3hJUJOCD7gyrKX0l0WPxu6T8MwBeZqjxl1UxBs1ERs26yE5TN
NkXHLoTeJ9egdYdJgSjwL0bjrxIJXaHCa4ZMxVnaFwWBZRDJHWyYy1yBq8wOMbAi
n2sJNtSP5S5hbc8Gy3m+H7W3mot+3D4UvZeDVRS4gwypfNFac0YyU0fK+h/R2cma
APshnrjG8dcXQMj78V2RohwdFl76uQMXVmYahq5XljjiBTE4nUjxGe9XY49+Fohc
sT0RpFmDf/psvJfir8KOREET3oXFX4XdfeYxZZUav9IIrJO2jfWcb0RoYwDUbFLI
tVjOX7r5JIoVBvy4nI+TNKX1CtRdGX6UuV7/Fn7qJ1HFea3sQnxkelLZEch22UPq
QGtkQEuDaMVUmR6iZNyKoMtuNfIH/L45olm3LMscmPf1CJr7XoC7SHoNgnvdCbs/
/Ti7+I952ACq+T14QdXVdp38lLJJa6l+xKnEfLXSrpCUA6W9E/oDIQnvxvxbTLWC
boPr4h9abUALk6YRmcKupUIg2b9kZIBvPaPdjXyrh04sUhLF9pRgGZk95YjAxfIA
iftrJe/BzfQ9oFsYTMcPfCt9lXlr2jNtNrbqj+6/L208cybkNaS91W5p2JUjwJag
2krozBEaS4FCc9NjdEQLDHMtry6eg2uf/4gfYsL7RS2v9FFaePPIY6l8j25f27LK
FfYDwC2d77becR8ilYNvBxUG35JoeUlthbPSW+LK11/U2pXrOq6wWNEKPfN8YCzI
UyKy74rZvhpppmrDoA8KNityZGkvZbpeHvqKDinewyjg/xte2SBT5NaVd5bALGiP
/ufkmI1NK5e98/Lq5tahtslFkUg/p2CgGN7UBOdCMCHdSZJ9AjjAlPe2R4aZwyCA
NdNBvrGIJy/satfxm+njhxakjlD+M/M/Hhdp2reKNKzdSnQjVkvrtKnC9E8J/i39
66zrA0ZzrlczltSCXHpowwUmeCmnVjrCPmohUDbxsZYF9gtAqMR27HgUaZW0xrrf
ZM6vzYWwIIJMMSTqnjwL55Na2reI0MUrPCkgKBNshHZI/VuNjg9VF43rzBIGau0W
t55kP1Q6DYa0GxTmptFPmQd06s72KUh56yy19m5mcHNonSs/LzgUT50OcFbWAdP6
Y0DFsqNuUcd1iK4l/u8MbHkt/IkuGPdgEfV8AqB2AWgpyp/fuHM7+1EizXaYw8mA
xWjjDNb/44gAy7mLSGyV23DEFgbXUkjYOQ42iloDstlFOLwdSMJijiTHAQo9XZGq
nagt4K85cO50bFNlIJvAaXUCKnBfKLPdhv1ZSCtZUXL/diR5e1TyV/3nut/iSH3F
h91JdBNvbASNfTCfyAF1B5fquJu1Dtcni1E7+tOBVEDQnVhsqmoK9JZJbkVWFatJ
dOYlReFINXZk2VGEt8nVSA48Mqx5fZ2uzk7TF75p9Xd5ioFqRJxlr9pperBEHLxI
/2pO8TV03wIZ592+A2Gwry228aI6a/1jSDBSpZ5agXSOYPBukhSZ9+saUHsHMMd9
FBwgV8QNVHJQ0C7nKI02jR8P8RGDnGrVYzyU2BBHESBtvHBZgnWErEqO6GjoDj9N
n6xaqebhd+zYFgs35vCiKDKddXtiRF4Wt+NetjK4xV4MUi6nTR/3KJ7DwOAG7SwC
S237bstnqeL3HPIg2G8bTkeKRuNpu77FfsLIhCW6GdSSgX07HdU762CQGeZjJ9m5
ClXQoNXA2FD+mgMYn2BBldKxUzFZ2LoHwXZpLwerL0u22ihN6xxi5WjQg497lEtg
1t8rydfwjBtvDFDpcsVwkoOT8mbwcmOqfMfbZ5SQKAttD823UtyvmTsKdS6KL168
xgqez7MVlMDyvmgU409EVXEg19/aXu8hzCbjqEOAiahZfVQ0T+Tx3N/uMDO7uBeY
2C8gq6PFC3165olVz3TkKkqyeR3tvWHmzgdh3Dtpr0R3WdsASvctkJSCVLr7uGik
x/kB22PHDs/5FlpbYfs6S/JiIRIXPD3DaQkHDgOeXfzQdZ8cnbsyJ7qyO1l8TK9k
6G3CxDnrnWp61oPQ7NJr25tJJtf+1K7rnStBvOS/QimJiQRfz3E52CR8IHvHEH9T
C7kEz6C7JiIaiYn7dnxRu+Pf6fycmm2tiVS2+oCVW+m0Y6MffHjoFWhOQcqRbAe3
JRrNIjFaOZ6VcYP+N2CmS0RrFfIJVdsznb5PAxAXp0lF1YZu+ZhxQ241HHjHy17r
IRTtAgBhltUPWpIEPeXYTARYzx+dlk/wvGLR5Jqd3w7YrD2OqPdlM+yiO8rCWOfF
0B/7nfG+1TZ8m0HbSPJ2+qfeLfEBEcIw5XxUMsgkFJ9E7DLtPdpdTi1CCYliO1Ab
7DHHjslXAtkMMgPSDLvJxDJIerwxNCmdnfxOwpcxlFSYYTbS1934UMmFhbxGMUcc
Rk/VNAs96iLAQ2X8Tr9a3LibwxAFpZ7zrGKi6epYJz+xGoP1V1YMARrc0h6sy3GH
hvR6QEmZmnZ67oVgslcQ4eDYYXLdbhrzI7IweYvYTBPL+CY0H8bgGzfQCbe/y/WP
3Oz+9c/ie8J4Zq8Hh2bwBDAYyv7bmrdmFUi/b/4pb80YlfoskwAEsmmO5zY8nuP0
XVH5XJ/F2nRqeAeVWI17Z6MJtLF+wmkwZiGYfxpiq24wWLsJLB8MN+64dGrTKWlz
4Cf7MZSNMyHpdv2aMW+9aYNKYQLc1IPmWtE+UyuOgcBKeitHqoliDch9Wt7XAQEA
bZzdUH9qySGuzqLMeAGLDx96HDxs5bAFyGkTY8NRVaP4gfgj7lgE7E1q0hK16RAF
LNAw3Xlbmgh4rlrWmUCH2hvy1S4FFg1w5bmYWHIVbWDakSwkKAClD5bBx8TseP6G
0nPPNNNK8aFhVfwJOq2ef2pmya4Gw6cjEz9hRvyFVAKNKH58R14HkSwenTiSKWjz
NFK/bzpwdtKYCkNml0yiQX/GLCkhsXDbTPqihobXWWTBpNjZZ5Kj3cYG7skMDgzy
I2dsG8XEsb55mz0/qFJ1KUwsduYy/oSgZCR5fxsb4g7wo+7Vx0J5lkUGqhb12c+D
2t/W9SmSlbrpe3UpDfzmXqPAcz3rboTRsKmlVUbIfdjjQo/6/57goEkSkvDYqTmu
wuNvO5jAo8qaaIWgIIbqYuV6oaCOXFCa9J4EIwDeh2sPWRaIIhxld0Vf06un+8gL
Q0Waf4fYiWvO2qrAYFGWfAy0JzM6ehnemJ9XGoB0WF2rToLhNPtj4cBlm3BExJY4
J3Dpd/udKkC7zrbZQ/5OuXHCRAFtU6onrxJXJjRo9XpLiiU0xlTpJGfiGmxzPjAT
sQ2k2bJj9cKehxrgwg+i4+LlM3C08lA7BTPd122vxsHt2V2rk57TDvBNo9FVBbXQ
zIRXWfqTHTgCSWElvdjFGYPdzYaCb7tU0w8xyUA4Qm8NoQJTBe23TdFKnnzCVVwj
mTAwdZdXnW0lGIoxYV7vZU8fk3KvgQ2kdKZN26bLcVmlEYVgD/C/vFu5QmtEpj7p
fUWpTkixwyrYXN03I15zGPiek8QD2HzKEMTHl8xR6Q6P3EMm+/lOIiiSeQxPaqF/
3Ns9EtXBSFqD3ZLZD6RgXpH9AVJGKTSQVlyj4VK9ZlmXz3ZKKZ18VJei6d46ZEiu
RjO37+tunFR8ifypfdbM/4GFCR3AkUknvRysZeF4B/E+7SGApTLMDrwlQViqyJif
dsEOph7/FSqUeWHn4fd3eN2k7m+sUFQF5j6Hv+gJ/4VZiANrdFNBxMoYewS4OKnE
Xdb9JYbp/coybYWZ37W7q0qybxLxzAT0zoJSRB3SiSJ2K+/aaVD2yGcTfccYWAvW
Oi2e4/b3LfOStHOSUo6fBuApkOykqxYmdSUNG7gvVWyGq/D5LGH01piBkUR43j1U
iqkkhyxz1UwithLZaRsYCvpiVwv7raK2Q/y1/MwnROS3lMg2/RhbFP9YuR/GGpoI
oNBo86MihZ4Ay7LYPw84Co3xLEaqw4yoHHmbB+E93GECLbBGtdQQVRVNHL4mu8QB
K01dV7tGXEnrH+WlVQW9MXOHc/jK6qKADGXhTnQSJbXr3v0HMtjkgOBrmC0X5VUb
O0aPrdjgWjNvqwCROsDJXD+xCZaanrL8M1E43cRj8o0rHfgmH3U5nkem3Gbnz/DZ
eAThwcpNS140JHLuqlcUsskj5lw92T/338mCEFPymoAyB/MazW8g3JT5qRYuD5a8
l+x6q9podKsOrka1RabnM9F+LsG3AdxtESTF6L4Y0i0YDAgctjPzjGvTD/w7+/q+
/SUfEGHtZzeq3fRz9X9LjxNvCLlBat8Stqg8LnYcY50OYr62FWX66IxQUk4hLWju
ayuZJ3a4CEM1Z39CsNp8Al86WZ2E54fcWB0cD4Sw187rpMRMm/ilMzeljWQ51JOX
8slRGSpowl+8LF5M73JkgW4aE7PEWbzOIuyr9q2xaN+09zs4uLxMPGOif2kePHvJ
2TNvQcjZnxr4zZjJrbhKxdcmQIYxGgF94E74RSlsgDigVTcQMs8uYFE82QE7MCkQ
nsIRdl1psnT3wDm7vzFuTIZMXcSEYizokIdGJhAJ5r4Eeqa6GehzLaMsF9trVKd5
kFZ8td05HdSBDykhaJQ91wjW7g5ONbdribpS8+tixhFSGgv0m+JNgx5gUYd7dNI1
NiIqt7OnAigeOMd/4zKJH59ElPAdW/3qHcYFv65BkhsiKdfEuI4VX39uFZN6us9g
QuNjPWi1T5J9i9X8jZXBjHvo7kbPJy1Lljwoq79IZIVqEf+3eMnxJkMQUBdTdtJM
Xz7WfD9Q6jMtaYJrKoOVRczMo9ywbNIG3SYrrpj5IwYTjssGFfMtmSrKMl4gUbsI
+ptTAzvOVdp3tY9Pwu1EUU2TKZNrmWkTrkwZSDpkH+vrSClLUcjKugWDiGC2L69L
knX0I7QURjVpdi2d0lWCZps2sGyJgdS+kg0N1i+vlfKFUXz4n2ri1KXKYyMBfGeI
3VeZ5DgdECFrJkuVpBQqR1Bgv/AcRy5jif9NtaUtB5qv+Hj0FyXlrW8/TkzQp8dg
gM4wnGHs3SghUR2bnOlfbcSKWhQnhRoDuvvyJ/qNPIe5f1LdQc1o+251ywy9arwZ
fzmc0nDjJlqRNFJkg+qxosq5fX9J197ZJejmvfO7ef4T4CSpIrkNlP4JCQXsyQ9Q
ZXlw3zZy3NE1GS2xjXrCMAv8o+MCuDOVhOFeO5z5Dx+wqY0RXtrClKCAm8nEvTya
j/S/XNkmB4YSGZ7m2C/YC3QnCdF/kbPOSAfh84c0jetAbq4tPJKARrnZB9LSg+mH
o+rUvET+mS1qcYmAOMQ/EB48BtGeF8bySCqShRGmze218FYVBxzkj3aA7XoCkymP
J2Wmmtk5rJqM49swMZ6jESATS7uuZDU15Vjly4i5jpF5bKpP8MZHCKp92qaQNxUO
yJTYo+0WwR/VG6aMzYXH/RGNjYyZKEPyfbGq3y+Z5hnjy6fpXri2hL1+5Af+hhPY
oAQNTZbzlbah5Xx7gSykcD28l8Aol3oSOJm6SL18g/+FKdI4kAuAbUUtDhzn9gSO
1mHMhalfi2FD1jV93uMC/NH+C8Ja8wI5IiZHCq2I0W7AC9XNkuxPBSzi36gh71Z2
US0rpZ5BQNs9tfQBYw5y2na1oDrLMcqBbf7T/K1kiMLeqdEkOxm+QyFmbkyR/2DL
EUFU24dV8FcvIOI3a/2JLFLubmpSmHOSugVCYUF05UxieaufKy7fg8dJeEPpU9Ul
BxW/CxhZzUmaDzMbQDkx50Naats/2bqqDF8p4qX2C/qGv+RZhV7SvZit+yed5AvM
LTxdS6dfbLeztQlXLYJpBtWc/uk8p570Njq5jZXiJlrWUYLuhk52CJ0KT5Bj7K4D
1dxuFL64FJpfGSKEXtKzIP1+NxJlLr2FOxROYa0zruZFkUCIGP7tBB5wQ5UXMYkc
6RoJxR6y48TOKPxpGwob/kgc9CiEhYOVqlYrvOVbffWrjCo2q0kY3Un40z0w0FxM
4YE+nSFyhVzdes69upxRX+yNtI4pKKWCPnKoQhVFtNqOBc8ptgdqDcqoxwPsm1CI
MRfYLyuLsDbZpcxTDCJJvU3NeYC3elK5FPqvThiy2fvY9Bjnl/31DAHx6du4B+ey
YDiwkKbjoGIhMZJ8F5AoR+049OJLekpW0qWxw3wq7+3XQbodv+fOnvknWgESO4gK
HHgL6hjtmbBDc3wAaa76GyfOmaFkbmUpVxlnFK8AdptQgiyl2jf1Am13MhOo2iwp
z8p9JdEwVLUYIdN/PM5O6g/iP971tvCRtiir8Ta2zB5dTSvT0vJLpr/+nSxWYYk/
wMaN9XQKCfJ6qJPCmeyE3y425CR+VpoByqdQhYw49hBmcORJ+5csByIUxNyHoSKn
dhhCMOE5BgQHjJEZe48ev1Q1GPoknAeplK1aseB+or3ilhgxwvVONTmtbQVJcps/
SoPF6089eQp8ZEjvt0n6cq1CiLeMZf7p5zpWBvqv54M2g1i1io6tuJmAyGaPYMtD
AZFey7Qe7FJ62I0lm/f+YkPyuDVDgFoeLsQLZQz7yqE7HYQTnYFyy5JU1lMFZAB3
1Xkkkck1ftKkLXvoQYZ4hgKoHKJUrWQBcjCOQPXLV0LbNRaX2kIMYqAni4RZdZtK
k/RjzFUpiRU8eNEX49wo146vuQivQ28fFgEs2leSHK63lNu6GC0Mk7MCs79WiHa5
I/j5XfLW40tHEdW7PTTW67+Pm3P1+54EhP9LMYUQOurHTqKNC911yKQhUAeX59I7
g81xlOGOLTapk49xcX002gNmNIS08u7GgAsa5ic5xV15muKAldb2KaznDrWMyXi9
scX4P4ru+/oIZQfClnwMDARK6wQPD0wD7zBRRSP5YycznAIujC5Xm1RLFVMCTAWk
reWLKHin0cvWsb34p0/viDOSrBcCwNO2Je5Z4U2Jvg9eK7NxONcpLO9OKPBk6UEe
ElbzOZ8Vi11WjqwSWWyK6QF/WQP0ojpM8Eoy97So6KF8M9r/9VIf3+8QkX6TjY8g
T331gvzus8DJwd9ywAgxLRl1TwA6hJvzhl2Md/3IlbWdumqMm7XiJ1eDyTEfmRy8
PZLUSMJz36jVLicWsaroS9wZE+KvYyNYMeajxYjNpAQq/Dn9ObX1YhJI/xYm1B+e
GvvuZ/ypYtH3iy1X2LlE+a+8K5kbEs0L2N50njQ65V+LBQcRXkyqTtTKvHe5wCBo
vYeOn6+Oc1zNFABpgHzl3/Uec8l+hqAFmWkXUFU4UMSisfZGkZkqGz2/0xXykgEs
Sor3/frPEZYDf1TomBkuxcYQHkwDbcP7fC26S6ID6X0JpU44y9xT8iA0YPX4yj4n
LA8ol+y9ad67nzPUPjjkps/6y0q96WugEJX/Qu0H7d3HhWCpUQQnJi5/PE2LJ8Te
fhe2J6DWXFqGjDYUnVpS7qhoTAjia5RGwVxlvgZZZQ+aXRMcDPHA0qziY4eGQoph
lqzHuyjbkRYkPXlvrY0p7A==
`pragma protect end_protected
