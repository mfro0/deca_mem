// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KNNtDlichurHrvDUdQEo4yYxZONlw77+ZJNmQkSu2jJggVjYnUCdr7bJ/MX/+9CJ
3rm03mexlQAnf9srTDTrmd/oNga1ncnMacg4sNhS1KcXh61EC2ZT3dostEuZa11Q
Vz9WTtLysVZoRUjvX13Wk5dy4zJEFNR1/OxykzwDiJfm4+E5ikyBhQ==
//pragma protect end_key_block
//pragma protect digest_block
VlXbxRlhAVavEOO0j+cxjHnQnTw=
//pragma protect end_digest_block
//pragma protect data_block
FZr9t72oTJ3e+m/NHx285Eqs9BoRBIrajMfI+8hCElFjvCC3MaclvT4WZDZSpxis
TYDYSu8dXleoko6v8bwyYI/tEDi8QMtz8ewgLZI4ru+iQtVFGVtQEeA88Hki6NwN
4qwGJhRzpMZpKnCSGfHg60yLNspxxXzETZ5Fm5v0iIv2cAzSaxFXaQnNPS8S3kqt
DQZsZ/pY0mBCV2Ugd86FCLhV8/M+wPVmQhv4pC1NGaeu7UFpG3+jjxOxkmBPJFMx
kxIxOlJPAwr8QIcWitrrcvM+bt7++k1JLqiETGco4jZGoCf1yuOomkNYX4sUykAG
+ecInL1pdJXQuQMrKYbvwTL/9z7PvgAGy4QouoDqwv0MyPYpIo9vo9y40SOaedv+
z8FO29msRuybNdd3dufdTuigWtf1EEqBn0OOnEQtAHgxQqJD9RT42PjrzS9X9cuv
wyVvPRoEr7wS5XNqt4N5Bj6diDJM200sFgKBjmyXfGdXWEc0UTbUoNoWQTu/IORH
8RnA2J+XRk5owpIV9w16Wo0DGgkdflvdviOh0YdMTY0y0dRdsmbfWbEctmDfVQUp
skHg4T1b8DdtMrszO3xKaa6QJPNs2tQ9nBNZeP8owAjm0uUDLUuNxcMjsVzK1ljT
kR3k5rEx7Evdj1RruBFVCyselQJWvxY69c38QKmGFTsUE4SRNKrhDpLhCW9M7CaF
gRyXsQvLml38S7XL8cE2DBRyBMB7GPkdgELo7XPVZE/gDb3Ug5M7PLZzavbBPKcS
zF/SF2Uhr8WpN03nkE2LqPd3BFmhWvLiSrzGk46VFlolyxi7isHG6Zh9yGfWkV0b
gavu5G3bpQo1MREkVKCN8CnDWaSMg2uFZNizzQBwRfr59VJL5KZ0DIAwqHAxS7jB
lwRjL+or0bdsnznuJ+2zNpgFw0dg2hxlX+wRz1kIX+SPdLTLUCR5IxC5Vb0HJ6Xn
Ktgnb/ZE5TwSutOwa7rHam2epsZPtV/PCxKtJEVPP5E1uD8cl0DBG9kATmhT5u9w
7lPu8nKSQZWF8bOq/1KEXo2hYc6njEllPm+OxGZ3NVlbJH1EyajTRhvAPLxzaVUS
Rs5NPIz3VBiUzMzE4pJ+F63UxuL/SR8mcB3nke1ejOkLfPF1dh4V8jRKKBznnfRf
oqqzMJHxVq4NFaw+THB4wJnnZRJU7fMDwi/jM3zNAROAf00vbCqtCogOgn6aLpnx
Vn1vg5KfgEXNQy46Y0VJopiP5s0e5ZICSdrkMGXssIRy2SQBscBtXP5yRhlRB3Qu
cvOa+cCvT8LO6ZJiQX/+QgxRuqghhoAm5YEZhHas069XBFe0DE2TOzfb61mCRceV
R6pHZBdJRoQqV7uxW4G7HYJ3UkOMAB/CT8zB4SOGgPBoZMFTg9C2PtITg4e6++ge
GOx3IXulS6kyS5g9vLkkX8BCQNvUML2D5ueA8ojdLALNNlOockKr7B/alRQsU/F/
3/B0RbGw6norcRBe3WctXqQJPf8VwjBboLQWHKhGZey+W/NBRu9zR3lufQykyZhE
0R61tbGLAl9RQAWSogXz0yKCBmnSRPS0o3iFi5r+8PnkZL3Z/EzFFv5JET7MKyxi
fHFZk/PtFCFsNf0/LyEIVWKHmGUVKPCdYckAUS3jY9fB3oOOLy+3nKWFRYGbd2mA
vqOXYLWq7SpaU+BgAc0cOQwbsjL63bYn5l8Blvpch+0LlmJTuvNE8WNAWnOhCJA2
s8nUslLEIBoSBjjIsKlLDJ2eFTXaFB0SUUq9vhEKl5PDOeX6JMqngjpBO1pAFwDq
5zz0TqlklCRVt3qJX+yTiT40tYLIh2J70+74Wud/PzqJOikTSknozdQ/4dfuEm0U
YbY0nMZH+MKxhSAVYw7hAEsvvQ3u3e5MVPlmegKixk/ugKNmy8VlY3HweyuQBqco
ciIEwlPrAPSjaBQt+cqAUcrKE94haRWKPYKpeAQOeU2NWNCwz4liF2tbOXdKXnBQ
NzTIpHmn/xSO9Zxkq9ufzMsftccyoPuRXRr+nFsCPLoDqOFqeGa6AJDC+delkzrQ
u4oP+tCO67Sc29P0jOFQKTGbMMUI0t+QSCVMUsMDrU1w/ogCDFxvnq8rT6lxPaTN
704uctVeqqMXIvAJG4F6xCk0Y+s2jXN7+1YeC/8ldhqHYZYl10226Gw8Zw22X0hx
Cw4a5cv75x60nf6PI2OURIFtgc0Xc4Fo+Y2q0S7V3dmbLbpUwE2FL/fDFYW00YIu
poBq4jtprx7eT9dWO43geI0uT1aKcXZuoLjg+G2oBCCZsIHWlg2f6w7g+JU1el9E
WvfMCdzRD+x909n7pCEOdLkxAeip10iRd4T9tNK9aEk8e1p19wnZUkuXLkTHDAFd
8py8UaZSFVcA73Obc/3BWpbzb++QRThg2saRgwi7bQ5k6XCz6+Vt1Asm5rTAxl3G
2CfaO8uV6saa+JjFt+hj3DzWoEK8jTGKHvqL0XVS9dFWUEL40k58sgfsy2mzN4yZ
3j0kLVaqB2HaOvoTsTy8FKsmtQ3UbO2N7t+vPQ7F0SZKbnuPK8MxRuYdClYQmad6
/0rP6xd+6+8/a9nrsB+CpSXFa0irDjCrMp4se9Je2Zn6G48Vo6uZhu2uUczQ3Etv
sbCReSM5uNi6xgvUki7tSyFXkgnCmrwOI6KuCiuzHf5TpHndfDOQcY3sL/y/4sc3
U1yrrk+fCp+tOpL805IUXpjQGClIgMR4LbGLsX7otEyqssxDzYQchmtzOkOhZ2Bf
9ifAJZdnYEmbura179+982UjIcayySpMU7aup0H55cNda/RcBiVlWyfbeL5ZnmTP
5aYDaLokkh2gzck5/9/qzwSeFUsX5FR+Kh9olhDiMhmsjAgzEFFd9dh5ujLeuLVP
deASDE8JQuqs1zJE+Zb4ahWWO2WsKBq8elvCELLb4n1qkwUOJYxLDtaroAiPbEDE
LZHnmP1d6GDHVfqR2w7VZBQ7dzFrz6xpVWgO49hrqtdHwSDldicZFIKLTGt0i3+J
ONsEIqEx3Y/gWPzulmDlhdMgGyGQjcJ68dN0JcBZ3K4OVGe1U8SPTaVTkMyCaBa5
FC6jLQfYcWOqoNjq2BljgwmFAofO+6BnFzssp2LITafOU6jCqoe/LCq31sgR9+K8
kAitxnMLbnu3+g7BdVxIouXValvnnSKAXpy3gTxykuCoPo1BD8pmX10JfxkwW8yk
NEVEKUBM5QW9V5olf0yErv8SPUu2da0X5PBGLqMugwDTMr47pnrG4q97lnHtx9JK
M3CiE3HU0KmhZK+dz/zRFN2U65jeEikeQ5cwlAjBCNirU8kF+6Thgp+hJj2Q43cC
9wC6eblWBcbm9FrkHfECG8EooudQwLZWzrVU4LhVp8D/eA4fccIpZTUJud+ca3cR
Vez370wDJT5ImFEqobHVngghklv+O3xNB4hjT+XCXjHJSkETvKyxQJN0uMy5pii6
ppbR4jWYICD59wDDQbQwhcv18kh14zf3EOrS2YhTBtjC0jJF+yeBzgr6FZB4NmpJ
6kDWGFAQqhGKJY//wjGJ6oU2yhFVbxToOrZIV6nMIpGwFZR3U5ejf8R5TqAwHEEs
V92Ljg8gARkbvYgacPNUKBej1GW7JNSaTBJB3yvkKcesHDEo5etathJoIGhJdwB6
Eg4AHwJRz7vWinJf/QKN5HJ/zgPzQAJRz8ra3DIsfOTwH+5xglpuJoqecvcPClCF
nETLSszfFi3RLCWXQGAjtRvcbK7RSUbODP/y9n437lnp/vfw1GmGQXfxbVOrWwei
Uh+0JgFkvAPK6mlMDoz9vIK/iGzrl03cLNAjYTXdAC1UUbmOR2hrWMaDLUdtxuq0
6aCt5lNVthiT2BgBGQ3RbKOX3gDmivsfTTjm5oyKF0GN6ZMBTD63cR1xfKLKgHAp
D2w6z2CkW4wmFORrTlGlI0WGY7lR8UuR6LAwcqByDhxD+F2YPMjrizUFXPtBb7yI
LpX145mVDX06SB+Xs/4xmFMBa2vkmfvMAxDnHeikcKuQBTXKkIC8JcW81HQgdzjM
JyJynzn9yRZQNP6S/Gp5oEeD63s9mkn0eFF0nVz1ewZS2Y7dF8qgLKdmBmUEPMCT
AoyrFzNvHuGHZDPCWlWg9oY+4zLJQW4G8kwGTZa6/xcKnOSe22KYHltcBszVZgLa
s+4imlonHSzzWY6sU2USkyE/ncmewXCr64mje3Ge/ARhtWtZuNj7OmHk6wwTfRwk
ZC7/f00BQnGzn7iiUPNLuGND9XSeLEXxWjxOigFUYFPbu3ZPZEPG8tAreVzSCBQE
NjHz04qHg2VOhu65atAtZ+K3iWj8uTKaaHpw5rNnWmOePChKQ/exyBFhO4hREs94
vZjVF4CE20qn6EBKJj1fSk16qPKAlzksWs+WDaxt45VDRpjkIyt93f6BYMKK+wGc
o8q8AdhWBYxaPRj6wQYCPmrcK6MQwEa1X1WCSx4MmECt4fOPxfjEQSCI3iNHMouv
etUsxESBIKBlhdWMzNP2mo8R0M2ODuPJYuxdL1OFj46Bgc+0jdDt+818hsyY7GIK
aSuRILfQujbtOadeZPDoSfCgSbcIlBGc1ysA4wxiI13fukz3ljAWGami7KML+XzV
5eqBuxO001KrXASPbSVP3u5Zz/y8CGJF41eX6sEJaU43YkFeT4xh4SLqOUklbhAc
d6vqFbiQDV1ETtVkWszQ/qxuwxxBHahbO6HNqGOK4lKcAu5awneBwsPHaetIltrg
Q+2KUPLdMoxcUf8eS9pI6MfGx8SeJpY/TvW2Kd81Xo0pZMotRxSxTxBCeFAHrB6c
4OKA6t4mDLTieQlAv4Xmnp+qvkqN2r4170FzgF1eXzgrIISKaSuxntPP+ZbrZ3Hq
y7xGFGIVGS/xxINZPDLp0yCN4QOOXUvYsfJpmhkSKBGAHYTqA9CtVhnK694NPUFG
914VobxG8Qcnb8oo1iWb2hFoKq2GKZQWf+psSD2vmOna80YeAbTBoHb8FePry7db
jebVR8vXKND/PGwqcKnkZ0z5lWwBE5t+IFhlhdRZpxg6OCNsZEtDCGbELv4bTdgQ
+gkfYiHpOQb6dN2Ws2r9mbhYvH9WoEQi9t/z3A5mHcz2bPnv/Dgcyxyzqto9O3Ur
lYt5c4NRU8n4gREmRJcFr13lwbBp/y9GXqEKP8MT5dX3myg6BVE7MxYyHWKLFn25
p1PamEAja2vzAbmf8YI0T+S5TpLzhBHryQrhSIKIugLdkWqtNHHkHVVve0Bah7T4
TuUMiSvuRfJJT2eIJHzDQglPPkdDgDwyirvjM7Bc5W9g0qJMLIvbs2WpNWMYonc1
7rbHCBQbydwDyc1UE3rm29WS3nnU/JPACYOOWjdjwelKTctzsPRleqCok3qnfXEj
6Mb6Y08LnM1budzdZIvqev5+yIrTe9/g+Mh1KOy4dKibxJaoWYIvy9IUD5B9GWJk
kMsYlHsD3ShPq6lXZKABmyb4VmEEUYfI3YuD1yyI73u5S+pBl+ioErJ/oz5k2exq
HiN3bkfRJsO/2qjQ791Waoj4GIorBS8YE5pYFuzvzkkTuqW1GKJZWeySBQRRiAk6
/6iuxyvgm4yt4uWz7R+9MjhW3LleN2SNL3MCy36qaiMNqGmdATe9MdsfMO7O+VAw
6sTETplWnA7MySvb5mk2Kgo7ZhfJOkEF8w6Khga6F32gB2MELzoLjFFAESWmMIc2
3b7eVGyTeVPmNBPixqknDWgJOAFNBfkxEgHl1Rkw+kTVEk8LL2IfItD4vn7acgD9
uhMGZpkRE6QDwthRqHsmgCTVEYQ7ypoHA8G/7GdQMDPztPp9pYUoeQulp61gPlww
tG+RKlJAekEYm89Tb4S4hOG90wOcygql7V/FGXH2n6CpnfbIf+LbIKmRuiW4wWPU
Bo9IOsZ7ZbAnz73a23JyiTOnhBmx+QSuQSn+CNF4epomWrdJfNKrAH/e9c7k4Xc4
kGK96D728wj9qWc0MZbo9SeeH8uZJwcszEAt4lg7hGGsz+ANbK1L1+4Q4wUkRfzc
dWtThVkp/hTE3KgJdwI2gNAhG+a1frYk/+CcQOnsxLWbkJsyr+3Sl4Z8Ku9i+1py
HIjeLBG/OsYDinK0wTjy4TogeGjXGETJU4HGpbXPFkzfgc6Ro0YVrTrOAAS7AIIX
1vqqbnARvY1IfL1MltRGsT/WvzLl6l4VW3X+aDyc/riMgjm6BWC170KHC2BIJKCB
bd0BoeJpYhgvdOV6V9qeIZ0RgBEFd73IefO4eCXSoodmR3URkdiNRTkPsKUFU60Y
T1n2L9F1PETGpdd6s6KvaTjnnK32F14B7hvGJLY7oy9acLHPyWknnF59YgFGmbjT
X5cBANZAewPUrd8U7UMczlhFMLlt1JIals1TjC2xfauWLoJaAwU+4R/oujmvPVZb
n0irnSgX1p9WEwO+LCHLD5e6bag7e7UlE2D1QMHWmVIctO7chkwR6E6li5GrqCgm
I52S6ZmTzmfYzRyJdFZDZ41kjjsRDuw/Mj0mlGJV9OiSKLDijgPRRBFmXswGuzAm
eVR1msWrtsPQsQM7ZfbvXttp+Eq+CbGjdFRxsBGNY+rdkmZ84WY1lrX2fkddZ1OI
7w5jZdvZ6J0GxLMRuJmYV2hvfMlu0TVgHl0eDHnUM1WlrlO5tUJF3zjwb3X2jDb8
BUPVVS67s2szFk0k6oP1cyz7j7Wqt0aTvT1RqYigxKRkt59fhgRrJfEqAarFyBpi
eTEstUNq6fYjriTATH9647mS7pvsx8pOOUOVHXKzW5h0st5ScGAXZkvUV5zroxXV
ApdgAtgZk8aG86Q0t/fO/8OT7jxsB5kdMoKMgElDdtDzTxOPTi7ArtzTyUCvzSs+
pteAQeRrQ7/WRfle+On8KMRcsPcLr+Ad3yfmSPg8Cg8X1kgfUy3Eh+QYLYkmU9w7
kEVouJ2yeqXODDka+sh8+WiaDPf/++xlp1eThhoTEv2HrJqQNwWyk35hbo9+GRB4
w1VzDlGEWfgwMQKPuXzSp803NoQjly+3Jip+AlaTFmN2eTI/LfVXnwbtnsdcQemI
CYhopQqSRUY+gYYpHPNvHAaL0nSq8fb4grzEjSWWjkCNvFS2ozlDHyjj2s3suqHw
Fun3MV/XE/TpkVcxFwdlAzpeeHJRNm0T8/6+dk9IjCS3NKawM8fmDZkP4L694Lx3
YuieAMq8rAcVodC2edr4rJKvoax6XCAIPlCVfNynz7oW8lC5A2RoKX3KttaXnQxR
6TZtNdTEXxrD0mok+66Hg5GIC0Ixl0lPALENA6eNOUuXddtgH4Ik2fvpwZVmwms9
pXkx0ehqf44jtYB/bwTLGs3PgvfTJxX49CljFaF6ZdtBIDnqLFdktBXMslLo44x7
6rCHpDNRVRoH+GcKeIfue6Tp25GcW3FBW8hw0Qy6TXAG3ukPmJD7DIAkunkGhDFe
lIQBE4N70xJYVxqBOuSgru8cM3as6jU5OQ1F3rV4B6OOIaspg5qjTuUdAdLdsxGt
ohv6mBlawcuDRXCZ0GJmjA+2Svig4CIG2Yk7jzRPliLwySHSChOEJSSwX6Y8kx6K
5O7k4RdK/GXCX97p6wL5LH/TFa2w8iXBD2PG8QM68b2E1cswncROZdY0Qv6OuCdW
CP1ZOy9O76oDN+65agOrOEMTxOSgNdZkqlVMUD1Qjg8TYJpg6nM6qvnmAJoEo58C
tLnDe0oEHMWZyJspsJefw1wntIDllsiVCeL0H1p2LJe4y2vSbyQK+M9t9FZ+0ibr
Ca5XLN/WJ6gobTRzh5Qt8xSAoqf+eUiz9YbY/bLZDxT8nGhiefAhISrf2iXC/gS5
Y/otrc52huKRtpvhF/deXSz+4YqIptLuKgTUjmboSIaGXzjmALBxl2aU7fTLY9O3
zDR48nwUrwSl0jpyx9Ff/j9rvheqKswRVHrAvWqZMA8MdncGfrioQPlLNS4r5Qwf
5xuM6+/yrAfOplseKvQ8GT4WxoDKaOA2yXzUt2mVTDUL2IGaP7OyYfaZdBML8Sjl
XUYMP3kcKgzbDH8AeQD+nPqeCFFD9lD20ZQlcqmTwusoq5WN6C/GYgu5WWMrRv3J
CQ61/mu/NnA87ePtfnS+J1aA4ntc1EIbAockLmVRlK16DWXm1K2lbi8pkVm5Cb4y
SivIf4cXztv8vMfD9/U6ovQY6YHcZb2lr+O7kXivaaL25mfxLcDjNQkj7Rj/iYS5
lYYc9GvTO+DeUu6vy+egRZxjmYPWBPd8uuejQY5UseY476J4y/0+5hodvg+l3xho
dnBKFvNYqRP0DaWiZUM6wNgqgrFnEJ/lhGgLiC+eLCRq24Ra9N4OpPNxrePslIAA
fuBULYa7CgmfVL9WZTsbDhzqh111lullpYglfSXkV/ceuVbVF2X9M2lnw2mDphXO
+E8YDFaPEPXNKmQ010VHY8g5t1h0ZtZcd+rwpqO0WKnpYOxiydKb73imDbLFmODD
dM9Mt9k/2gQnBDeqqrJjnrBgVyrkNlN3a2kCyG7aGwnuFHNcYo1vDqmWP2DsobVu
2st//5sJ7IEt8nDVhjwoNYjuiGDySH6TUmjiTjKsHj/ysWEl2UIOnD9aa7UTgty+
YS12ocHB0GCiRY4PprxUI/Y8CnRU2LvfIVIru6mp5Uuukbp6pzwtFUtPjhIb4kS1
11hR+bdqAQQxzXYF2AyHLYgz2SG6OSOh9f4xj1aLsZ8yTJR81oT9v0nvg1MXNU+u
DSSBko89Caw8O43OqF33Q9OLjMdWaYqu9uwaHseZunktRKlLw4HPTdblJT0bTFDt
EogEdhXqgfuDqeAc64nJFOu2JikOwAP1B85PFR1aZSPDT2+QTcqCxYkI1qtIuFtw
+bysltUTMZIhyfze2oYFccpoQlJSJ4fqaBtNCNWo7VjvSD8VBIIz95h38c/Efgdd
I9n0W6y7mDJU15do+oojVP1gn+v2CP5+UWHDfIEDcicTM6KhW+zsz9+mTpfNBu20
tQ5PajPEtpq+OuzCFuTwEsm1jsHp4xRyo8SphLQof+BfIoxpQRHSYB/flp5uUNbq
aQA1PFRpVlja1MsZs8lp+C5ZgBSfpzMqecTP3ImGorvAX7hz0jEYzW0H73J3A/do
//9qP2M98UHpK0i3Tr+cI8dshDOePCJhhIg42MlACBkLTn+RC4obc+Am72lGbs8o
iCrubCvV11SZxlqwA8ymNbpXyi5uPAavVsxLmzH/bLE+sWatkSB+hfqbe5a0w8LK
JAex6jVqMGU4BjBDCfogfCh6csdBexJWT+q9pUWScBknksvUD3/iBI/bmjj8j5Bu
N+UiPQw7hVrDbsg2F0t9Cltd+Eld5PGi80+bmwawRnKxpny3URa6PKjxOlWi5+e1
4L6S7OLEz87lZfmDJYLDl3HwS0sZNe9vZFdTq/CW2zp0RCfefPoqLyszCGpqf6zD
6SvhJ01JDu03PQZRuORapqUcyc4k9d+bgYAZgkMB9RAkmrolMI3pxu4y5cetrfdm
64DYfOdYmj1felt3eGLZRkZ+qRSdxT0bsI9uVuBWVjWqi6Q1U/Ngkx8hswTOG+Tk
7c6l5h/mair2aYzpM8PAJ4KbN8vAwMG/VMsJhcA4zJC1qJd6S8hJIa7tz2TBzuzK
L/GKEkXpy3PXv8v1VGGrICgmASfMzSKBddHKQdOlYHA0aa0rehG9PDBD/4HjRbmr
2QFM443ijP3IuOV/iuAC9BFaqmOsfEL0cZ0nhVMp9vgi39D/U14s2ONv4K77WfhM
Q45xAVQjVXkUDx0+TaX652wGqo5ayWvviz95BG3jLBS5XxESr/uj62Uod+9DAbrg
EVRvEbMfNqPXLvbpOpa0xJoJq59r+zEbfUShscIoc+sp/TWY2r9f0r9WFZwXr8u+
mYcmwiGeQVBkgpSs2zrD4A6WpuqLi+1tX7QC2jsJhZUo+Eme+H7lI668eqJQG5Zb
Te6370pZqU5qGlvBfnRQ/5uQLcy0JXxZ6MK3d5pyWT6aMfcyjNWiEjAsK9ksox02
vNKrHbQqAeBHmczvbXGWb3QXwICBRWsM8/c6ar+4iN8W2dNYHoy9JFpUC/Z0CQj+
yjVMRqhryY/pBOPOanDT3cKPaenYQoh+fGXiTye0/OqJdiPTxgWNiBqASFw9AqAv
CJewbe8kHVMqc1jAX7D3wRTqfG11dLLusDEV7EgFQlcmz508kRs4TymXiPvQJqL4
H2Pt+ye6D/QxUnXoUfMZS6kQLUEls/2q0qgSyWufaeA7/kVdNNfgME21leM52G/k
ldkTyzaoAxMQpZbtJziNgXfwY1AD2+FxdPEYBrcNZ2Neq94Clb4XX7uDzj9cJh58
i318VrEFyCzl8hYmr8g2GavfM9EQH/pqo249qCR7+K7NYrk1NKMxDqLNFJvYMQsc
XEeHiXPhhjBmZfVF/ZtUDd22MLW5xNKXuye8guSmc9zFh3FT2iYAKg+nWorNsdQ4
OgjVb8kp4K5bVWTczY/dq9fGUNV7hmCd57ZXnsANyD3YXD6bzj4QT0dQJFRN9WuH
zQRXR+F/b802Vf/sNoRVOcfmdw6KQFCzaG69ehXsxqvh5ggj8YXFa1xKSVWk5YCl
8kPIT0mL9s9fuTe4AYStZmJcYuTfLVelkSWy/yZVCrE+7TscrZHNxgYFlHnyNP4V
+wnLZaf54rrNOOlotqIAAUWpiCwCzz3dw7bhUZWiSfBY5oMGQ+GAOjdrNv2NRw5y
w531Pw/drN9mjfnVk2RfzwOZ9wteyyz2S7T0izdiShMXyLRJpu4pibzOJN0VBumO
c22SqONGzv4QIDTgAJt189jRVJJ2xa/ONlkmvF8ulcpTEk/KtRuPpBUdHyrU4oxd
HTG6ue6lV45fsKiq/SZXgozaj3Slx5+dwA99vG4GVOBiVVbBUIeUgjLvVgSK8uvW
MTzCiTGn3HZ+1Lp2IpcJ02nBrTzx+0GPT3GyRxElNAJxyWhzoXiyDE8S9rkvYDzi
WgLLn9skCiEH91JY++viisKlMyb9uxh42ubz8+GZlSmwSHKzj+DRfcm0jeSw9HC8
nFrWfVrUnpvUh4OXiJkQUNWvPisaXy2IFlswEZAL2nLDC9V43lFlbFzMcQPXKYSZ
ioJfy+xxTJ/1+7P66hrR9WcnJIyjnJQk6gdKrB3xdvmn9rruVEcpNuz00KRkcOfa
EnHjxTREtYmIRDwQo9QE6m4V0WaQGoDFPniPAIPn9/dek0QV6YT+pjP20h7jw3rQ
wqjszsq6IClf2yYB54zk5ZoI7ijQqgtRcTgTl/BLvHmbC4Y74a7kcTwydmY3Csh2
KvWO6vDfsIA1DM8T+Md+eSjWsG2eXSOc3xT4q04qIfEqlag66o+lYn6PVVHNzhSk
fhOUm2KakSI2W+NPEpNmN6OrQ3wOYd6mSZ64H4GMpLurhDAdZFhslW76y/K/D5e2
364U4ezsWfo8g+mdyDm1xAnq86N7hxKZ4tbVBNrfLaUzgnOxr1pk09VhzDa9Wqaa
zc9uskNSzPdUYxPWqJWxCqtI2qAzhY/VWFB0FvokKVDmgiXjdr6ysa5uOyhuk9F0
r5QBdrDwVhUnHYDqNnjf8IFQn+tmlPV/GIrJJcxaw/AWjivn3RJ37epXsRVA+zVs
1aePyqpifanuCOgt/FBMT5rqP+Px/Flaaixto0epVZXToKTCzmNbRombTCtOTVk4
VXnp+qJ14mbIh+PX2HeJVQvj8AB2jZEY0XHF7ucnE5Ll9qL2cpHpmXBSxduCRHF9
yF5WlhGptfeKSLAxXpJRAH+DOoLlwMFdIW931veBlyKrr50H2K8ICxG7DQ/HUYwc
QW5IqrUdtqx4dY9PvplunrMqC00w7M4JjldwnGFFjXfCAFDjJTA/Hc/trh5ugJ1y
zlZyO6ALi2LFjzAIP6SlpxzBdEwtoqdKEqJmZ69b7v7c3WuASIgMsEIHCNXIZTgc
YbYjVQHnMVP8CoCeMzTxL+a+Orqi0n3P4CuZKhomDXCLjziCifwqi517T9Bk/PEw
lrE0AvNv5yY4SraE1S45uXoUCVavtuRL74qFGJL1LyxvflDYtGXf7J7ZNF3oIM8R
1rpIidbcHYoazBdjeQwX19mqCbRJO4wT/DEYcn1inQnnxA47WBh5a7zV9ci/Gleb
XhF2MPgpuHBwUyReCSikkNj8NeTNOwk3DwHttv+99weQsLXP+KHGw+eCQPwf3DG6
vlmFilQyEli8J827H4Bo1rR7isMYyWURMH4bXSsak75vx1+qcSdfUMtkl6VsQ7MG
dTtqnA785zbsGqCeznIFRbca0ScJkM6WIrQYT4H+wXGef2JU5KvlFPhvn7wnN6x+
Xji3Lf8Xrl7NHWHkKKta7Hah6OpSproibOJ+GWioAq1sfYqe7r6k+mJj0/34TdT7
VPWB5my0ajd71cy1lvqlPrTdhaLwIb5wnPXfvjmAGMf4vbjUjRO7ph1yNc78dsS7
grgfMGmYyuLjdaGTlmgBlfwM7Upcy0TgGP5b9K3p5UUgIPbmz4z91XZpfF6GiGK9
QDGfMYdWJjgK9Vw/kX4NaIXVP/5TBPalOHBySjD7Ywowsd5CGbbwGGcTs1oQgqWK
Am3J900ROBI9O89a8UXN9tcAf/FKo+BBpFgd7fJu05UEYPZ2jZABvJf+7eF6xlG6
M5VV4C/j8Wf2GRXi2FT9OgCRUsz6DRw3A3LZ1YhZj/MnREt8roJFwSMz5yKmXPX9
jAN64dbQ2LP0l6qextmZi/Nwn+UzrysYDOaxX6QkfSktkP9AvRsSXJ+crpdMn90y
+B8T/9Tdz0XVb3m9aiHy1xnly51bUOIS7VAoM+GfgSTCutBIqHIhCk63xPpJpeso
Pgo1U1uPBeSrR6zI/zCQQ4rPAxpnylnVkIRXGTUWOa1WcSK0WL/fiThFRsxtHImO
W7VTJ+2+K6gn8MjunPNc6cQxUChOf5fKQOf40JBwHRWB7bXHZgtWiRXY9Mx+SZKy
iXhpr0hPOAn3h0fH1gPU6Y9Hi7hF6/VBvbVUX5d+uUJM/J1jDyDeuQ7sC0FvBHMg
/+OGwCvp36gtFN1lTi8gqI0bMaUHdnWNpPPwxCut8HbeweAAMrDHsDxQAD77YPRM
bfpL/vUHQf7nnJUflG5AROrNtOR/Otu/siPaESGEMbyoo/yHCG3ygikkQcZ8W8gz
WIc0syTe2ruSUSjHEP4w+h5aKXJ0lFiZeMN6ygWOK/NxWCy2F1eJBl3+lepf2lt5
VD2SIxCCkLIBeODpPUMXdI2d6En2dfpJhZliX6oE8oRoh84IqRgAkMg9nnImJiNx
19SvlulTVyipezIdeG0Rckx7U5TIaHw/qp2fWOdEE1YhYqjaGB6pojGvxrHlOUo+
ahrsgql/Vy/NBKb/XxRzuhJLPBFqk+q9Rs4eeSZ1Oyeb7e/hB711tyK9w3EA84Go
L0fMjLjQsLxb+qtlOdE95HAvJgpzh/NMrAanP5zsqAHRL11ZfH50JtXDgrigSR6j
mhTs5uDDzc8EPk93E3Rfx9QfYfxvpGbyTrIqoYc1ObSK74SBrHzTQjZOG208k4pR
gHi7ic+tubWZGUSkzVDl62qDqWAktPFDaK+DeUdu7PUEtKmrlNafmhTlmYj6x3eL
WxGaYHiCsiGbKT3/xLKOLZfgQyaTYRFKscvfW2Rm9t3wRdEZy+2PatS0jUF04f6+
DnDrXmggjmz4Z3Q9Gr4twyKfc/xggQf4+7qMYnmgX3lmNqqCQpEmOE2jPc4cDZMP
0avGic4pqpbyRmLxwXtZiCPo7k4qMKBKRAF+b+5t7zHQFpkIlLCxK39+AmePUgWU
FBllmBpENUITpJLayi4flVhTt5aeIeWURhwCOSQeegLITYXUXeTv5Wtkh8ZauWea
Npgc8iEAMV1MkDh038H7apOgcc96jouN4nGSqtzLqu1rMZBo7HCXDWejr4LBwNHn
w7VZz2cCTxF9ousLy7stdCNKFwke9mWLy4Iz/QP5/Bszm0e0i1+xEbg8Z4bl9gva
/B5OtzWrPVwfcIsggYW+FgQxYCU8lXGZM3kCuGgDnO87JYwbfzh9aBJ2y0wyF+2p
kP1Y0xaX2hoReBWO9xNdm9MIwOhoL5FpMs2otfKrRO5MnAzNaNm/TmeQnPyhKf4N
dKErLcvM5WK4sBtzBtXwecVyDBZ+0MERJtk8PZFCuEnec3KKJc+PtTtzkjr9ebkw
EWjJeeU/HEet9FAnnrRT0Pa/YSTLvPCzvIMUL5bzu5zCm3xyuAe85trU+jlMh73j
MgbE5Ektfh3zMjzsEWCbMKtIeCjt7IP95MNA1PGwEvip7VQKhaSTxm2sFbGUsvyP
tddmcH3n/x1/woR7CZ97ao5vvISJPrlj2e9bVAk9OMFnqT0Q8fcy17/lsPqVlhWy
yL9CR2OfJQVrBQBHNsu6ZpPTDCBXGIb090kSFPixKM+o0mG4hlKMfxMHA+43XNvz
NMwKqewssCCBJNhLrBIP9/pYR3NtQ0CwKxsLDdmrX8i0qkjnoXlz1mN4q7nrdnTc
7ciaDaNaEe1lxzMtdFRr/yj3oPjBYV9ih5ZnKMfy1/EU+QDoWcQthAzaLY2NT4Ax
FW4Or/sRLdrk49yXU2GI79AxApAzPvocI0ir2Ct2MFvzfuplZNvIcXW9bRkL+zU4
epJUewj4YaSHtyo5jeDDFJxOxa/xD7HJjkwh+Yb4lrs8/ZqIjZGdLd5ctZsmX4nP
06TixhbUqffEzFg+bAg2A5ZwtZ678XpdvrewkuOWOCuLNispCwjp+SHhdz9RQEX9
Dh6oeo7194KzdR+HHLDcmErdAtASwlHSAOT7BuqHQKh6KjYKF+TsT7eW5Yp5c8nZ
gxG3dxxs8CMQJhUew4oaFV6gKcUSSr0Cs/zXIuMX7mfPTtPDLRsd1gPWaaHkjyyR
mAYeQSwEFfTZJmXSrFnnJdFWN5t8rCE0JbjMyWJ8E5zjcihQcBFnaEcFMbJU8vp5
0/fzw7j1auFZpNsTIoqWHrDl/rNAUyBt1byt+zhxxy8hYjxWDc+VgrnP+QgMx0NB
9VugNPfV1vaRRZ2vuK8Kd8CHpJ18XzHUwSeB46L6BPr8YQME3RQFtVRDCg4s4Hxf
fAFfa0qkvQYDdP7yMCux61WGHPXCtQ/RAdiW6ODMt7uLVWtcFe5YwxaqHlo5GWAQ
0oJ/9uMLxJhdrSJwe5lqn6B6P2+I3skXmLkKJOBESAtg3jebzcjcghZSuElaSdK1
6MhLXAloFKzm8Uze6MeM2CzWkDHq/OZfP5aPa0rKhw0xZyOiyQPYmIA9NUZTmeXC
T07Vicga2AEZAybPSAG707lmYkDIhb5eXKkWpscNh9wZHbVYIiImd3mv8NOsRZh7
qyP9SULt5lg9p1NsCHmWD5PbJPw6Qxgv/NcgOPp7nYVH/+dDEAy1t6HjGvuMBRlq
lkMoU2Lir8rV9cOpSvof9Rm2GUmja2NYTZX4pmh5mWxsv+nmdcKE1xVVDDXGvm3W
7oohfaQxlB7mQzmtdBPk6iyKRHTkSOui6VQRsFTAamlhVbn1sAoMDyWKiGQEryH4
H5OU4LZpe8f4KKjMqBk9+ZJYQwXXwqZkdmIrtkrO0vxWe0QEV9Y6vMwPfuZRMcJh
FQYB/187HRcjgoCKF5+k3IIyvVHI47j4pHJj276ivsPhEnl88vEiPnBtuSt88VHb
WAs/3qvn9nJnOXuPu1slluAuthHl0OwBh0XSgZ6mYbVfZwnpmXp9oR7YhvRLJdPl
ahm5vwMguatXAweTp3FGYDZS0hQWxhIeDoX2IZLhoq7zQaQcVpM3wJpEXk4POb0m
6LyidLVGfeYizyQCJD2XuhhBJQfQw5XfahhW2wm+XsRnVzxxhroj7UdydeN08jgj
ft0XUzL6OpIQZqq90sCNs3c8g//MSicaDZsgENncC7jcn2W6iHoh3jiQiVWDxAVU
KoX0w4RMhkFCDn3xMBVpI89N00dHJhJg2lwYNa3XaMznjRCO9d4UqryDp1Dwyg5q
Pyh29YmSn/RoR9ZsDaqTia7CLbbugPzZq3batSDEgP8gCcCgE3pqpIhHkbN6zVBw
tFO6YYqRNqgOGj9RmoLpBBGaVSLHm1EJM0VbtkSuHi7MObZpgOvIXT9sm3G/lesG
tap361qU+FCEy83hJpg72dMvXkYzx5poSsigqnIMm81qC8hzaKVhIPwY1i/UUujL
Xij1KegId8r2m0BaoUBk3sKdlOa6rZU/CaWO7QKOliknsYVDErJIURYYhKWc4am5
3C+FgcAW/kLLOgJGs/J2u8Ce/wLQAmd9p0oq2UUNClWUYibxCDnXzkFga+7xUibF
UW6cH/3MqR+luJb9b+jYhpR69cGWleOTgecTkeY7SbSwr/q7PHOUo5t+FnhNBsYK
FHPUDWO4gb2mFYTy2L6a5svUAxBO5/R0CihAq91h1FyUrTVH7g8y+SMx5unt4mWQ
78SHfSBNjkPWWIXpecOion0X+UqT5XXaMRetDDfEnfAPjnR3uWYE/awRiyW39p7f
7BHXnCZfiWucivRuQi1Q0BQ3DaOyrCxBI9xUddgwqYQEWYmSq7MjoFXCoptK6zZP
0sejmpI4eUl9NLvN24/P3JjjRXjpS/M6BhrXl89jxhIaHh2ku+6N9VPs4qBh6YdP
z8S7dXcon9JfBWukkDVXEZlcYonzPSiwjm4T1C2rBIs2Z4QxwbGmo50GfyHPLYuG
qMn5biwV3Eor6DviQS6QOiC/aBo8jVDJf44juget6t8rMl2Ekxw8MsJOmz2pyue7
Hj1PFZvk+ifkDirvmSvhFXFhzz0ccuyD7gNsLSThY0zH/SxbsYjSpMaIbhyQgszI
ye7Mj+p19DjfM9D5js3W4Hy1o8SIvHM7iKU2CQQGep+635VlKtkZQBhiua6LNzXa
OTxIsxJ/MqoDgQafo11OXbcL2WqFHumSNT+f4JQvRQEiKF9KjcQ1AQzPPTSDgFnj
hCRaQ85ke9R0Es9liNBP70PF8ZzTG7mK6hqbVulTIuzjhwUiypjO6QS+0yd8X5bi
yBo2zAQgzY+0LsVJVUF/U9fwVz9VzH8rSjHD6jOiMr7I+axU+IzFrrIub4RCBR7i
A0HNJruP1H+EK71ni2rZFTMSsQGmUlUI8fx9DiJmaNyrWCio/env0YQY0PrlUqOX
pJNArDsOL0ha82fiA29jl6Ug+enTGx9cKh97orCs0+wpYZWwwKQFxB9OQA1yi4z2
Wv3ovVhQFM6xLN0KDLNANyN/CNfputOldZKTALulo4R+VOBEMURuPFS5QsTEqQxh
J6nH3LuQ8H+fZEH2IGFsA3hV5NadepRs/AotsOb5UdPDe/MW4I6JHa6fW26OWlWT
2PMCxXIlrH2JfsDjNyrGgRTYTK8sdtimbRRXjnwmGpAAm7ywoLSkSE9RZ3Aqyo6w
GaSw2LPP6Ite0YFqWeuTO3JD/vLB+nI5ACfEgefZx3o63Ekj5ZASUNXFjHnKypvq
PnYXmn2mjrbjC0Pi3nJI3FFTTBnK565wdLrZgthhIxq169Y6Zighq4HscpJvwlqj
rMyMISe6DHb6nQdd49c4QytMCuake2MDG62easdWbo0EYvTEFpXMC31mA5vOcaLK
DiI41J99lmiuYRhjhCI/9aCXJmt/oVFiNKhVCo4YMUF+XqxbIjcg0t3N3Dbd6m3t
L35FdvB5rr7bZ5EtULwGMCdwLjcIr1XwWzdRaNvb+BbwCw9pnTEPPSN0soVPXbHJ
lZHhPAJGcW4yRubSR7hw0NMHw6enID20Hu5xm6EAmEy6hKpJm/uE7iLjx2RGRK3N
nW3SSqpq9XTHysRqnjiP3Y6WKRqJz4L4quiY+uTApEMNZ/bldhy9oRfXkmgvl5h1
G3Pv2hdUfkrcpzl8OW/ENOX4LIPA11EsAFSnZmwdxQdPOSfW2Q/wlYwbsbxKmBLz
U1jy/NMR+uiig7EVH/h8bJQdJHrfw+tB154xX72eFMbx//cds/1QXdlLLG3yl2of
iBtvyMCD/sjiWSQKujf3KtOupKWkMWo+RNtLT76u/NiXcW3RTMNyCyF5ncU8/n45
pDvz2ePZS1tlibCQDcJw455Qbq+AccszR+ep3EnW3p49OrTZCTUEz0idjhwBkb8I
uK2aID6OzSu6wSuR6A2DR8rAp1+9hIXHl9fJZPULkB6l0hLH9VwSUgxf8D9kzsOA
Db5VmxGesicJwPgSRsR6CtlJbrzABcsM/jXca0VyjaX1yZJ50JCsHDLigTRgQ654
/KiVbdbTE/TNgYXapkIKOgNZ1enKJnYgCwO+DtKInHbGbKQHUWqV7aPGv5r/6nqJ

//pragma protect end_data_block
//pragma protect digest_block
5dGosfRCCP2utBOIWFSPnJbUDdM=
//pragma protect end_digest_block
//pragma protect end_protected
