// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
V5ZZu7ubMqaclW9UfS3xqDE1lTPQsTxUXlNnkkv2Rqk0NPDrZpRGYGREkW1F0X2J3ipKmRHx3n8W
pz+sK9w8X8v4co3uqd4lSSe0zHKdjmRTgHXRhQ3MKN325sYPULfKYvP/DjHe6vjB/YzhsNqc8kXu
uZMbWZBHggl6+9ehXqm+tv7dhKikIKVAOouIixYsmtlHhu11U1tvxqtMw3dtbdAUBIUlGpAXDHtq
kYi0Xbw+ikHxr28FfPIFcbj+GRdq/wZoPk53rARfRV7T5iByP3ZJGi1ut3ddE/OIqyBHGamyftLL
2DM0dB9AmczJ76YqonvB12sQaQ4GO2BiZM54LQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17376)
p8NHmonx635B3RDd+X8P2MOFcG3iKp9RCooyi9PYHw/27h4E4Fpyw52fIaNNBz5sdypBYsF2n2WV
gVCqq9j5HiCx2VDGUeuy2BN0S4E+0/uSe/YF0lw5SEP+vJcObMbddUiCI9cgqhZeftXzdgqtlssD
+dywaGf0xonLdrTZM0wp99Fr5GMRlX3eK733CRJwYrm8KZ6Q34qVmA/95Kjry7LVQb/XSRgD+JkE
0ZrF0ZF6Nz/i1skp6r7iEBDaKns/yisyZEi7SB0H4zXexG+U2hrMzNNf4fbUymRFrwwtQRFc7iDB
RYI97pSPzREVQZVhYkT36PBI3gn3E7KQ07WAFEFXoHgYdfy2SqOo+lf4Ro1gkh3FqphvBy5E6FDw
1DpXsuN+D4D4458D+ToCxBQsu7bOP8xuS1PL24cMzU9o+v8r/0yf/olgAtwjXQrdIgMoryW7wW+I
ohbRrbNHlFfCtykiuiflmED6TyCcVtVoqabS1DcfOLyw5cCEaht5CPXdB5JoFSB8iRbe/UflZ2xv
OjYgpGf+wN07SLa91kdevvH5ZRPs+8Hi3dqsjAELxQQlNZ7sy0/A1spaFbmANPwv98BJEVG+9sO5
DmklEiAcsOsRn9nEVPTd/xxTobHNpO5ZY2CrD6kriG3ZyikeoUxb/mYvVSb1W6Ea7ZTR1VF4QoNy
2qivjFtoyzcgZ5oXWr9U3m62we4khMhU74qJtxQj4l0kCC6ZwmzjDzJ2ZqhkJVTY3u46lQQ1YYjD
99rKSuDJkEamEOP61dIr9b9LhUYMnSmr67SefG7OiU4IQnqCHZ3RlFdWMF6QcQQZv6OLI6SWSx1J
9eG2AuF9tmZZgVqwO8yCrDLUKS9BGzviHkGXJ3xruJu/D+hdVEF+448bX1IF5egF8D+aAi3uWdOu
Y7vsMq2as5sbZRX8LKEkus04BMemTgS3A34wOeJoKncPfMaMm+xN08t0bsPzIzCdcyUX+v24Zqi5
ZzOSGX5Uz6lGfSEs+WK2YvzNnctX7qQhn5YN4af3ABeTsheytVpdV7yDqZlKsoC+SenLMs2zVEAT
4TGabkwjTEl1n6MoO8plFh011c51PgVZNsri4DJTUwOe+6dvAJ1x6BVZ3Pmpc90F6ijd2lgCbLVv
OciVh2CzZCJJum81+wa0gIRm7Bj0xHWRZeetQUyYaqffsCXP4REOUp0bLCeD3B5A2/yYefuSJsLw
pl/yfX30ubR2MsfTN3C5jkCvjirb4I7aGc5CnhGNrDQ2dHQj3AVrDqSSOPoy15WacPOT0MkcZ+/G
SzBwFE10SmD+Uxal4F9tEJlmcJ0bewsTwc5pkL5lAmggyKigSUdi2pa3UGKpQiuq3kq3OUDbcLeG
BywpoVi57wHCsRfxVQHmMO6CEj3xIGNz7jw2Lp6ERrPDrTPZUM7LYebLHn41tvTfL8kDi+KifRJH
mnhngBuvLlHGsoBU1AywBXXKr7ulPhB3rNBkLc4zdcAj2m4cHTMY3DIejj513BW6MENiE3O4GX/G
PIrqzpaT/EqNt1bsoVnOYLIhVl/QECx6vwaOhzgFPnbn4EpLt3Yte9EqwL0Klwp6d9Oz4X7xXH4x
A6QeMZUXB1uorlOycEx7gpVnKs1BTTeSD43bHa2xaocMuma6JW/y1GcaGgWjY6BoZ8DRWUt8QCJC
Q81IWcP1A7PpA4ukJ4+38hnAzmpVxHU9t/3E4XI49syTU2gEEowyVK2XjzvwBSICmS+AwXOMEz1x
x0xypm6rZRo/ashY8zX8d3BT+q+/CCWdXpKlFNoMsOwdwYI+3dHCIMx03T1r9mb92GMzrZwsEsMt
PcfpS3ar1xtvjNMH+EUvRT6Y0IqlOpuT56DcBH5hAdRyVFeXzvB3tuWO4eeavLBFmnkOV5XU60te
Y9SDszssjyhIqJ81WjyAiB6m3LCwKu1x6plMT9cmU7bVHorPWti0JrzWg1CZjRwHb3t1J243bODN
+GRlwNQCrONN47jC97rp4v2bpwxVbBoMpeDhZXpca7UXsALddIpAHrYTTQ+2L2VueEnmejeBBgK8
DLdl42UwTWcHAv0FvQI5A1lWRfvRdgBbeTdJX/jnvDY3Y2UhdGQZ2CJoNPpneTlO9dKb3Dw0lQTz
lrNV+aa7uS4StLb08SNhCCSbO8erKq3JEFUnG14IZILy3dlpfqTOc11ErffB3fHUWPpeoWkATClf
uWynRg4E6V39KF8DPmQ3MiKlneyxdqqhelGLe6r7fcQg41+Sswj2UPob/Hs0pflhT9Rv3qBF+lAh
TPILeLNfKnc+ctS4L1iBUc8iAFiXDBc6PoTjT349TjwwtQCOIwW9/C2PRjftpfIMuEcgzF1B+93o
MjQhDYgGsuDFdHeV1k731ARgAgotQybmNmW2Id1O20eF23TKqYx49l2AIMxZwcgMlkInhxJ4muAD
1+vLc0I5ln3XPKV70KwkJxYK8bzV6FWYLO8BsfrmAqaog/EHLwXccNzHYl7Ah/wpK0z6cLVBE+HX
6CKs82qOSd6XsviWmkAq4nBFG1tB5kmWjWfaHGMTbq/NV6E+lLbxaRXKf6Q5zrTlBTDp9j/cUXOi
tBAtaEz2HzjCsqtuxpQOPm5rk52eIcP4UjROtdVkx8KXHVmsqD9n24nfnjbR6ND0kJPjBJOrSRHH
eBI1zTPjpxfRe+p+1r/eVgpXCERfmbvgxEAFcErkot1b7DVdR5enKEyCN6xS5ofLOrzh2d2XydIM
6vqjVx08I9lyx0iKneqS1ZrQEODZQ+y7RN/RSgIueq5CYxoNQLVHp274CJyVgXJsEoZoKkwKfoDr
yTifoItPXipbu070X4avqwHD48u7Ld6A99aWrzEH7tKvh235HX/Y43u89EneHpqF8+5gW15JMUOx
wD991cHBKFcTQkKXwkRANT0CBl4Pvt/SOKMQLwxcXw1+3VIt5AvfHdolZrigKm3xma6+f+WFVoOZ
fkDlvnKG3lAxiKFRvwhWrTYBZZSR+PKa57x56B0QGzjz3SjlxLSBaEGKEHxtbgtnFyCTqK0qZ+B/
sCkzNnVXk2Rc0bDUKiXz2BRZ+gzELUsIt9WuTQBBjlfKf+At25tDQBZD+8RP5PiLewn4A2e3OEmD
yvppSXjvAjbqPxG8H6w+47MaWMwMdn/CYYEWOMWbhG3dZCnkxXGkz35CwihecUR9Cve5gZpm8INP
hCLl7P3JeEHyO/A4+TgP1OMkVLV1yRG2B8jDQQSzYKSl03l88b2ByC3GAES6pbBgn/rZ/z25JwVA
ksb39bLA0HSc08qtshiyekDXXbeHeRJX5P79Z1szDqKcuKbs+lHvXhbey4DW6yeF4SL+UjMRGajx
LPTv9cmOvXHpWMTuDQPqtfaZAkBmy295gsY1t9294eLByAj3TjnPFIKDDgg9ozP4OuU3HL8b2F99
S6X2r8f34nvlGHaW6vuamJQUpGKWi8Ka+g9qwsf3Yo1IlhESCEMpwHCNDpXyJXYrV4pR4uLB3ctx
UBkQSwi09UkoNM0GwEmzlNer8GawhcGXomfr1/4XpHMk6MwJhPOemjsa/wZ4PSHZcuXswlFvD34N
dFjjD4T13XeyoWv1PrxMBbcReSlXq9iqPV8MIVi5vg+m6Px3mW+eYkbExzURhbQyJ7L4bbtbeIeN
B8NCM7AzaSRNw2ux/PfPuSajhsER/mV4op98vuT3vAq68d3PEWO1ZZDw+rLdh3cwaZIFXF6KDPO8
ovi2mYJWq6kihIOoPpUbhU3ouBZiZaUHIq7AT/9r/7zkN0SACbnAmiYCPfyrJL2k5YglXpooPhOC
jVoaNTmk5m1bwtyWVaPVAxmJiM8MA6agJMxounzLPSGAtTHo0K7RaDSFKK47VM942oFqO9UDlw0d
MjyKvTtEMH0UUxxTJ7dDCB28FwhSbtS5pfVV7cq2rVl70RxP0Y9n8KOos1rbW7bLXWHaIzwdombI
ipEXZiN4Ny2bu8WSbfRi5fG58GPXmb7vCniVII/TyPhmRaoemITJTH3i94AV4IEdtj9/BVzSxdd8
+T5GPUFhzT2u6ZqSjwpRslzObB/Ryn7cID4UQNanAfVm756+odPUqXKlLp1QNRQZFadjA0h2pX7m
KHzVYdcCNWDFIvuXyBPKH6lWZadbdvd1uNLe8G6Ah95wV0c924CerXx7cWfchbDCEuKK5BOZA/NF
OSTr13XMuilVXkPDO4X3YAcR9eX7oxpxQkilR6zWWnKFp9pV8UVrfX8R0wiv1AZnT7xxWL3BsKvl
YvZdZLeSyoqA1fBcZHreuL20pljBa9qORGNC2IuBC+l/ZBKPQLmTMlvD2Nq1/j667luvz0p+98De
1IGE9fziKBj7BQxwsVmkSUjdrLTj56BsNLuqKLpBtIFRsL12LQrAL9dVAgXHaN4VvfLqn+YjEzc3
GPpWUpcBn4MZqHRIR11/Ewn1Dfqx2EsUWulzFG/875YdUjcKRhVC5M4DbAWid9oZertiR/mwDbPj
0IXw8w3gF139HgW/dJfeN7zaJV4V0G86pH+EvV6rxeODRCJoig4hZRJdVSHqHKY1MJfu5CEE6zdL
UFdBaZvXpzSvEd8SL/KU7KocRZwUMarvB5PHxuJpcDocIxp2J37BAClTzSN7a9o/UmegXk6Y6ouq
BrlQzgwSzXcPwHmVHSqb3VuayAIE2KUomzduVUFnJ9Vy1dE90VOeMR4rOnehqdKTM9IlRD3dzigf
twzEeGIDaI149hstTwzM1uJgLs5W33+AUD1b3GAAoziMmSJ7R9A9PHXWZee3kVymp9dBfpN07v12
VR2BlIxWUZbX6g8qgNXW0t/wmVQliMKnmn/KGxaE0eL5aG1xwCthsP60v/6OVJc1CuRevPeTOwOL
IAfTfEa3g8WLjw67Z1Ss7MBMX+2NCq70Fv6/iQyt7/fWN6Ec0pJxpQdvvJCOIzn3/mR7sscp4bGf
IP3MzSQEN5ezF6Y98U/TFp7cJyZSOb2KZTGKHq/UVm/8/pJbZD11NF539BstZIA+jCr+o4XJICiF
S/+L7c1YMHpVpk3xg6yp9pqKUSPVNwkykPnlItbx5DIdORbnv02nvabmkk6c34k/T5b/2mgPMcBN
IaM5wji0Rf6T7TD0ZnY/c9LkLY3hwxdDYL7SqKUHbh6xkqDbB6QhChuD6sa7lyxdGNEiYAiTon1A
EhjjsOUwHqCx3Sae/hoj6EtHxln0y8MOkyibLDpOCBUAAdBKsbia34+FDzDSuoSHnhOuATRBXKM3
7/nIou3ZjgkK6q+tpNG5+vhMg+EB3Ep+k7JId50zGIYOL4+epfPMv/MM5GtW8N2WuQmMjHBtajT0
mDw6SUVFBnYsq+brjkxtJc+K6I+kS1N88dbshy4aOsCAS6GdXxzttgqW2uUprbPDvbNwNzAcdjhz
lQugl9n6fF9odkttgyBFaJLYLzDE1wKiOXi7U5I1nmc/anEGtL/i78I84C0/c60U6TbtdIaIcjNt
ROQju8HvSeqkLdKzCn5jVEw7aexO5KlrPeeVmEN5ABJIHd3Y1EB/CYrh08qexLdbGRm5kR2SlibM
7W2mBG5fC4kutMYhM6KW2UZon5DeAFCZHMh4xAQi1TnJhdeSCtsK6PNxlx2O1eUhH2bjEtiV0fKW
pL7ggCaxGFXOd0Pu2ZKFjm0iJ5AUhoYwE4kkGjC7Jhlf6R/7tsCYHZBSIubJB/mz4Qb3vDaxIYfM
sbp3TuMVwkBOWCMcZtjtQqODQY7izXOfvaEfswzFadt1BxKXPuFEIh+wqAI41YJa7Jq6qHfX/3NJ
vLH1JumoVxNonAZYceKWYRM92a6xWnRJWOwJqGfr6Ra0ONaT9vSLmPpeCA1HVjpwymiQWLhFI8JY
SN0XxJMLtKVSydKo/rOQ5H1/fiNDmbQTrcopTEN6yyVkr8RUuAgKS+FXxkrT0P9mMlE32lMYlz7q
Yw12rn7ix1Y4Xx4V90JLqDR/KZPQFAaB26DLQrBW9C4VonwxNonLdl2Y36lxPdSOfBPmeOzVYIA8
66ESJzmbflfrTRraOrojjci7i+J4luDXqWxNzsiF2dbolke5YmAlOjpW8mI2EGlT7mj0XTOLnbXS
4edk+9x/C0YJwWECBi+A6AaVTmuWMKUNpTca1eaKoK46WWgcjzmEhhvQvvb5peTSuGHVia1wi1wM
yiUQggfN6syovdiJZvncBWDT6+u5lzuNlrMdfy3c16RQXrllsMz1FyL25Sn34OZWXoDNOsz407me
egV40Pf9YTVpfngFDX+FDonGyBZKX+ZMxWB9B5HRaJXnrOIBQ5SIzy02RHDFXLDnHRF99GIQS85l
sk5QcP5tLXDfTzq84R+3Zmsuaxywwtjaqd65vSHmYw9UYOHI2bDSEEvlnyokd/CNq9g8qMf9sKMK
vsUQJi4Ls6jSZcp/xIkr2o8PZQjcJUtYqvrfBeqAtm1W7Lqs47kFCwCH7Xmw3y4kISjOx97Pjru9
MufhzZk/VkycN6dvzdqZejCfG2hkaBzr7a98VGqOaL52au+RtRAvq946XbHNIwIMtPOI786dltmH
2XX5dG5RUVIHhUYDo/fH1C+taJ9EkEmZOMxBf4i0V/jTvns6BKbM+dkL4WbslUJ4bqQzrWSoMYlV
jfI2uf6mCSOkpAoC9ceIXCFaNp22lPheOU7J60RFm6ZIVM+hxmj0kWyEGkWQ3yec0RPh1kmlYPL4
0lMcXQOe0M3+nY0OmXwhWyDlt56Y/gmTaXW11/NflZibLJ/X2j6FpYfz4MDaZuDyt9Jwf/bl/YfR
B0W+/iW3ut50WUiWE8Bv3DklqFgpTmpmBOrDtUIxDB6nwpP+WevFpwQVsTWy+CpXB3kMU29ywpLM
+aCYFfOES51wfEwl33FTu5eOgOG/WgdolY68MoGdpvrA+rbnQEzHgs9Hw1H5JaM67D213H3god1X
u+LlwaH9/auiVq3rzHZuR28CxdHHMYMpiE8H6ZpatQo5w8UN3dJdAyatXFV4mmlfPckOCVkHprn8
8M5AT4olpgjjTSIFNgtLwr06Hve69Jl8D0hknF6aemlRyoP18+iQAfyUGhyZmXINGjVvy4aO7bt3
nszf6NFTzl2j6yONS73fuocz/bpiTfebwVqMFdNRhCwESwQGEVCXVysx1+wVEC19SY3ZlYCYGAYL
P0idVz8BPHKdEAlVwUCHwNPwbRyi6gifeek32RIj0JwCdMc6Idj5PldUshBCJ0S98MXr1ePszhOe
wnzVTnS8+ZQ7qZoTlig/yE9dVvfDwkriGRHFIQAaqW0hk4EFxk1Jyurp1hNJn2pslpAuUZEC1Fv9
Lri6M0vurGgaNbkSS7Ku5yjUDkEcTJO1VLVNWUd/HAkpanNK5EIbuG8bnh5sUQ8UEEB1e7H5mFQQ
u/j9ssUcyuOXd2sys6uRnY0LUfSj0gsbZNbsykr7pP/Ujd/tbLyZXXM1Zov+IpYP8JCgexhuDD2c
VZqk+bfei3KrvqwcdKQ6dwoUsLXDO5HscMIANED86O6MDyf0iNXM+Me0fMlZp4x/v/I1HAsDF6s5
ISeTIm27ksVS+OCLoMCASjG9HPdLs7cWwtWQ3lxFFq1zY6G/UsnDD82St433Qfs7Y6HyHqn9KbF5
E/ZGNqFaEpLgd+zOLpW8dggQtAb/OO+tklGxTX8qjV8EqU83cuOp8qvYezih3v4yJVSddsenMXch
KLX9Y05oX1qY/ZHoO1JKKCAxBGNDQRSMKE9G3UtJpmyqmqKAHo03oIerlq7PdTbepCRZKUY/zKTz
BUD7otmB6hy+2Tuh1Ka/bmfXb/cj8l6mZ5mcqvupj+kacqRmZy/NpkBqRXJiOvaOHjoVheoWOABf
Ud16XRz2Wb7+iWaXtHCegGi7Nikhr5Mr/gCicDNF/WEidh59OGb9YwS4Mz60aVjWAKROEOVFjI8b
43nu7oYOKcUb2lcByRZBRrCcFbPa0k1mxpTK3vEBdND/KobqCAp/CO7Uq4yCX8hGwttSsX/IAepM
j3x0pZ+0XluNmsu/bB7LZywY8VNEriKzL8oySnZ0cN1AT03R/8TJAoX2WPDGpuyTZbzTMh8Ka8PL
CwfspXE1N8mE0B3Ubf0j8iP0dJ5CYFNVki+5FRzGroaji3wu3z9snP2uBRjoH+0vU3Z34+NBOuOz
826EPUjFSyd2Logs91M7CZUh4B8ER/ok6G6gLWpVE7XTsT+DnAdP3XxgRxEI5hKqucFAS8OlcHqD
VqjPJ3BKZZlG6GfC6bqU/+xOnC7ukWOdaEQdJNwcgXydfAvf4Fx1JJN+tL9/whyzZVnBhgE6pUaz
B6OaiNKObz4ePtOnX1qEsYfTWi93/GGY/upl2twR9kGALQ/UoRV14hNqQecum72TJG+y9UVpd1cN
2X7e8S4fyZ3Vzf1wjY8rskS3onMrhp8GWp3VtF0Jm4p3cWXbTzWWPRYm2+UmWv0sCsojD4rzkPTP
R1xJssqwv2gdpeQ9q5wqsUBB+zPaMZIR036xrxk+ZN4pO1d9JzS/7JnHWTr4RDIP/9Hw65FgIBH2
NDLzvJoHPwOOBDYyAUBTfz40CLZNyJ2afHxqRx1qtl6QfHOXVIIFbNGBWH1G5ARCe+NhVgdH2pYR
9lREUnQ9+jj/gRYblj2FeXP0tK2McX2lbPPbNF/1LMsrKpYF8H0/ckuBnbeRFUGnb1ufkMX5Al/P
MxVndpVzYiGh38r9YTR3HzDf1cVz77lFnhl4rzjsSmX/ifb9Jtezpliog8smkS2ImXeXlncduHIA
GrKhBNBGPL4BszieDTqjPi/keJN4oR9BMZKH0gFbTFjQJTKPDi3rfAtcEazvEwNx6+3YrtU7/avZ
0PrRHIoG2XBHhtp8iylNOC9eyWUZuLwbGjgKlEBR8Nw/eMe0exGL9SnIKZT2AzUyWVHhKdt/Zy03
S84W6EYGSkxYHpze1qONHrNFpxDSgLBi5n89pIzNPdtTajvBCylfMWLuZaQPIGOKUgQRrkVhpISl
C1k5PG3vWC4I73IVCqGm4nMA5aVPrC0YJ6wXr9C0+ne2+ZIM7D5swGnsV1A2fnAI/4PXDClTvBvB
85Ta9iig4Q4uIMnZ8orKZSv+bR7/hjZ3fj9ehabh/Jos71aVpeJBQIzvqVsqdfyvWk1zJV0Qi/eg
mdJmaQ3YbpVrqCPXs0J+xSQOPchsW2s0XPIz60dxv5pikk55AwuPTpLTAOzR+8E3YMkgOZqpolmf
uzwOZ/OUy0/rWiB3don7/oiiKn2FVQ/I5/54h/xgAI2RSG0g/9u7J9BP98gn2kCrrB1x+67nxOSr
24aF2V2ASByY4jT8ygnCSBVp3DAzqs0Ss0WFawmovLIE1QL/edbcsIgNUT8wDh3R/9JAs9Lrn6z3
u13lrxuIi6UMbiLiEci6+srkk3TuqVMJV9j9w4lrFm2EhAZtCUG3B9tOvS/0V+THcUEclvm1qzyj
vsejjSdS1ZvMRI6+sB/0bWbIyWGsPsacX8KQHZCsCgFxJGjxxRik2Pp+PJfcsTMBXKud0YB+FwB4
hXiLkMeLLNK+QEQsxKoJW1KEYQMPNTGDfZlXUr5b1v6H3AXES3nz3GXc8esjD7qjyoujAs/DLc3S
p4dU7x6AnBVmEh8UP8boIq9SnFAQ9BL8Hk5xfn8X8Y31k7FXGQReom5IoillHIFoe2KnTQCyVmIp
KM7ICN9KQlux2KkuiCjhQVdPKaeEA/amZXHvVe2Mn4Hw0xgDowoBr/HU9kyf/jbYVBzbdt+ZKqhR
VhE3nPxTTtozoVkxgLhgH78/PdqcrQDU8trbjPJ5k/JmKVX98jOZUnXMWSqF/fuVXSHaUKFhCeCv
oXq58UyM4b/DlZgKVgdtMrSnf8Y7sNbPKnmTxknTd9y6l8Mtie2L41GR9QhrszLUUokp6bQ2F7Mo
XByU2M9uAXR4HhSu+Asnzuo79kvAA+n/DCxQtS9uCxp+vZ1SV6ERvo7DWqpTE5+P2qRFk13Xgzvv
m4U36oWvy82Xac3APCD4P0JFsmftZj01JU8UMpNj6QOb53O6rlAWVSCwAEbwBct/Tg8CzJdENSbM
cv7indz47DOhVoKBVsRw1kj0OhtEzOYP6R4s7RadDrh1T3yl3HQHn3LzLxKIqoOT3HiFiUANwqEQ
Jhbss0vWBWwS5RCC1usdbU1PeamGqBeXJF67khyAvUQLqYfmSgbnVoqK73Udf6egwraX7tbsBsNH
cvFXOcT969Q0Y7ooSTI51RvxTYFPDrufhOX5r9y0TDWROIClFRcpZM6R5bRZ0dP/ss1zHd89L5hx
aDXZ/oP5SeoZgr8ml+d0KGF4jYmgIjz8Pfj6bcAwd45MQpzZ4+JrtS51e1/35e6qckiOOOjujqhz
yeJnRTTYf9yuQ7RO3VeQobrCq6Gyl9CKKg6eVFzLPaJU+IQjxNWXpycWed+M8aS51OrgNWEWiBGz
OFcg/k1Mng9gVtmEPaHBpIf+aPPk8vARUcX+wIElayMF0nuTYb+ZoqhQ8hNKzxl1PydlEIzpUKuN
Gj6NX8J/q2lpg8f6xyEOFPGn9Cu5z+2kGyP0boWHvhEIvFn1B0Oh5lDsIxp1OrHSlobwdSoBKVWq
+WPGVXd2YzhXx0XTD87lqQXRmE7aDsuj3ggOeVUBc53fEVXiN+yzqlctAQxCfJoLHhk/IqctfR+C
UFeXX7vlKP4GaZpHIVtyf8JmtkxP4dmORB2xa2vTaJc9g8WKw49763ff6p2pg8QGili4OyQzuRF9
nqYozKYws3c7A1z57fbc/OuS24QM/er06pahvO2NhX37ZqKV8eVEiudKG8pruQd3p4LZertxXuIL
91cYtpQ+JCiTWdH3ev41r9QIgrHJDyBDAxGl2yX/g0ozzXTy9IKFqt0vn+6u7Rb4Ylbm9iDB1Tzs
U534YdhcnUdUBy04HFwhIE0XgNoKrW3IcnDenatbKedzGawK4kGO7DPuoK3vKvapc75NDJGjodma
pjqMriduC7GGJOBBE1bNhek6GLT3M0Nf36j3L6q5ZdMfysWaxNUGYiW045V5tqmvYIP5366BxVVS
Kc4j/jQ0sQnV3iQEQER90wk9KPiX9WEMlNEA0aoE12VhDs8UbQrx6QgzDx6UMNnpHM5IdgkePf4Z
gCf7cvGQnsB4+xNG3CH4IikEJpaG4lwfoKupHmU7BWDJR1ITeA37VHJzkuFuaBgCuNNyYNlFseBv
WrpFLmcF7C5mr886QLII7y4NAmwQfdNstWdxuEPw+GGbgqOEilDVFYbjEVpzYW18RRuvhOgPNmTK
YplWDr2hA3Jm1EBuFFo4XQsdXAL7A9sqOlGibHQq9ZeoZ+fbqNgv3IyiRYozKcsj7Q52kTLFez+y
jyxjaJMHOakPXvOG8OeTD6Q41VHlpt6BtH+ObcFzhh0Zlb3nq49Kp7u5nJ+HifjJ8b/g93ij/OCs
w7jsi/qwze46R9utAwyOTeR+WzYtEj0FVePdyWLGTP9q8NLa8H2XDsKd83a4hIhhUXO94tIw9M1b
f5KKtosNEXAHUeCJ6i5tGIzQO8r0f6R/H51wdiiKLXOG5+07gxf3f7oYgZk5/rv4aWEwt0vcElyS
EGQ/g+6sp7/NtKOgKE65rNKFUg4CdEx/2RZl1Mxo/bmd2UOH7Q1ve9HxomBp3EBEPPFfqelwNFRh
vHRdlY0Ta4Eg4T8z/CMQdawyrjjAmy9S/760eeL4Qun8h9hCWMwhB7YwEu9RTpfUkKYTtID2rllj
24pliO9W2Pe3/XQnaPuRsCsZ8s0Zf/ZlxAavt4vvR87hYJ5QTeY9pkFXllU2+PTzGSNATV2VUhT9
NJ+gXZw+8aEJJHEQbBokffuHeO2i0oP5mFITg3RlAY2/uIwJuCe0NlCRfrIznaosCSErue3LklnS
JQ9/Ba6LbQLIOlzx8mxGgxl0DLAn/mYJuUipiN9l/75jIogxpXrNWzXm0dW6okZm9TV7COTTbH+/
eJ68WoyG3LcoyNZr5aWRydQbRVNppp7+ivIkcbcQJbas/eE30wVge5iJgjxfU+wKwRqxlW7jF9ob
rDT69CFucLTskgV6wCCCMfYfC+r5JuqrxMo+Y4U0DguFgBOnFp3dCGsWAJhThZ0ZIaaolHPJWkrD
pzhb2eHnKR4l30S2XXdZPPtL9eGVrRIF45TKabTSEfSv3OcQi8+JP2dA5vQEqkcTwnRPc7hvQdy5
f7iLQAhvul8xGPtjAC0kCH3nAXQyV4hkmVOh7bj3Pj47nyMPV3oMBBsZp32kwvWqJDJhOPM8cOUm
akMW+KnW9muj8+k2cPMW7zKVstImH7fmMkC24gLV0/Qgh8pXL+/L2mIwptg03Y0spLtYYlKeY+hT
18x3BSWAczipv5IwHEeyrozDPyw9852eigxmjUpHxFDPz+zEFD2QeAMyu5hJkvc3Yp9o5Nx6MNX4
Q7w+BSHJ/uDjd6PvKeOVp0+mhwb3pUZp3uHiIjzGlcciF31coxUorquofqdKfHNAq8t5eK3/cUtq
5+SzH7qDyWqn35Ra8sQlKeuIF3yDer4ODr12vfYCK9pSL+pcke7woQv7rYS+X/rqX+/1jaisIMvh
DFQ1kMevK3CLPKVotu5ipVe0SXqIADebbw6JEwSfOiLr5gwUb9z7uuW3drOItnlp11J7NlA/YR4G
tBDrYdDUm3s0WpEO30R28FdgRm4Y/g5KyeU5C4OVOKdz7cqso2lEC8w/RciWHpcjTmy8qS8zGLQo
QBZQtI8aEyYYRGrs20lG2kqn6Da8iiNOqfMXHzaArOFuM64bpXKvFDBfaaJBqmXkQSp8vp/FkkZ4
G4yP1TfX0jnz2ds4LjuDSkXxBA1lPbEIsLnmoFr1OWQJphCiC3WrNW6QWRanAZU/rQeXMP4laL+o
JY44jIP0kRZgc1PHxgi9ESQRp5h4dnn5QiQ6Uuq8xYE4r16sZSQIhUvqR46b2SloFiaCWdVSW0Ge
ZuEerCQURqhzFbntpaiuIn3D0IsbQxqlJ4vG/9h2TM9GqLyMCpLUf0zN95cncqdd9Hz01tOgv8Fi
9ZxyjpYKgqMe6r0Pn1wmnl1Awi4xnGJvsRl7wcVH0Xzo+QdGw0bTxiv0zpx4Ug1QGNkK2HNJbxSF
K/AW+0UkLyz20coRK8dyZJsCQBIWCLJeYZ9ecWNWohMK1IJ7NYCbFePu9FR3KQpCe0PDNtQUVbgo
0wdFv1Ib/niAAwVGsRWnMRVAilg0nr2DJ3DE6DAhrQwrYRI2gsD7O0q4jKe+iXg9kchQEQMAy3Z1
gU9+sI23VKMCVlvQAIoPbOkYOiYqrQzwtNdPYn20WAFyJm+ySyBWkkYwCa7C5qZbqvfz+EzTZg31
2ViGDmEW8p1eQta1gFNsdkvPsXR5MzjWoQiLdHWWKnBM6OBLM7lNF1GjtOradS7QSSQXJTR25Gqg
yrVJf9m7DJ3P9zrU/WtVpuc92k+dX36b7qZQKlniOQyUg1XuE2QARvD1y5VdMJ30iSi7i+lR++re
xZdpaoRpH1Xqp8ZQ/I3WYskB9bXFnYDdFbhCsX6cdkZ4Qz3V+GwPr4keX2dNuAQN6NEmVEt9lcBp
D7C7jjrlnB07UcINW3Im6ifC6jCOtsJR+/lWxFLhEVKDOmQSIm8pNCahpktusGlwD7x2kGIdX9jE
MWF6SjrIOGQxy690atQLJJWy73tfIwb62fchUCjO0Lo4z4DScHTSnGuNiGbSasFQQ5lKbTO8qJ38
mpyZq6K6SEV5vAScEC119dYFkHvKOYNDuio13HpenR4/3j69lSJdwoIBbX0nWolcrZRUFzMwZNQv
9gRqVyWb3zbSfKA0oc6vxGdbp6vTUecNR/E64eObHneGXBy3JwaRyxQS99TjLm4sWjB/eroOe5iX
slTLU7L5vrRzeyqNB6oRMkzA+3WiiCgszzlEKwesq9GZ+s8Zg7K4MOd0D2rc9St0nUFphJhbSJPL
kPei/1h7/bw5R0/t/hGrRWI145XseqrBWHKCDGWf1w0tYWYz6V+5KRkKOZoHeLQc+gzY6M+n//fo
4gycTvObdzDux2Lp1E7lW7a8AGFPhoS9SEOzsWexrdLjXjD7mZ9FNi6tDDtOZ3L7lVGw1nKsvrNd
NhkMmcrMEdw9Xal6S+IKYnybKnBWQko9oeVC5HcpygCgoZDwu+1mmW4klukYnzJijveEddtvVXag
Qrobo7b3FKvoX9bCsmBTMUWTJ/xqjIY1OGecgCav5A7/07ft+Fj+5ZksPvTqA9qzRp5IlCrU7yPx
dARHCu9tNcq+mhMaVSQxsJrWcXHUJEU5kc42+HrJlurtbroAFyxocQ3iF2wcgAzFz+ulQLecPbKa
bHDP3y5+oJ+pcETKFjUsVDWmXx1zWfKw4LTffVeubQ11mDACqzEJRpLiNKk8EwoCs5IkKF1ozl7F
v/QfjJvLN5FgJEfUAOm8WTFxKsQyo3KXT7898Vp3ypImjAi5RvmezdRriYP6HfK+hUsjhySyh586
n5WELCD5CEtSSaaZB3g4PI+KsS5gavc2PbhtuykPHSCrDYUszBxZQ6TX27Vh8DK0ZrRL+zIb1T/x
ONACba9/uDduxbgVA7sqnhyoAfeukT2jaYKSvWmbfuaXVuVIk8YG77Qq/vIW5WgF4T+m8vNKxFMT
uLDVgOYVkgaPrtmb1Gk3XThQZ8kepsAQ4Ep26Ix2K5xvVNMRr156yIZdoLya/yX+WycP4EltQGS+
07GqkB5hO5YmfrczwlQ3yTmnSM9q7/F9nFkx8eF8aqYW2IgMvYoGOAynCmSk4QIJk8nAgALn5rSL
y5bXaVVorcLdM9jj9QMu4WP3bzTsw1wzBMzss5ytWzT2f8BYyzrv4a+phn7aiQz/FJZeYYtsJk4Y
6goxk4vyKYd7Uw46owLNoFh2a3FSB0D3TzEg8lKq9WnYz+7CKnK40Eb4Hxhshf1UIvCs213nRKvi
hcSH2/44nBz1slF71ScTm6XmvvdxJXUwOtQ8/A/G0QttMa/jhYQnMvHN0kRn+idsZ1emxjUahJIl
NBzgHVcuOCJy/OzhJ2OWAgYByGPalGnqFwPHrhkX/1ARu7C6IHlKsoe0oYfEtdjDh0iU3hwjCXuI
LYyOe8CU0TKTq8JIcMlAk3T5t4275Ua5PkugJgrGxzCCuIq2DlNg8SCybsDuf3VVO+XzoJtO7rqX
Ech1qPfDZ4Z83NyBP2HaxNyewgEGZK5tfV1cU77NIIWV5Evrp4gIvdpe56iXEMCrwaYtjfKVo1Ed
E1EMOH+VIcnjHHsvlh4pbteyX0o0AidcZyB8CN5ATVPSQ5z7uO0neSO7nSwGRUFnMPmGaYpJ57I1
QJAzL1NrVCwQfFqJYzUv0wpq+eq7D4njY+wcL+iWSyLN4yLmxbcrT5USiilbzbByrE0bC2OZLdug
/9faMqfGkKiQzpd0bs5JhDMCQonbebQh9eN9ILjXALKsAuh4egZAYowFmZWe9l2e5ichtLHEz4OQ
Vn7AsEaygR8DvTV+gTyGzVbVIto7GAnzvDbchGjgRzVi5YnkBtdycFCuJktBooUlfKLfTIdMD7gP
XabVsaWYFlrXmUzdlTC6pKmZpateXQLKTgJgKTSLj2/Zwf6d1Hy2BauIVVGFS6dAtkns0U5Cg50f
kEmPXfkrbBNz5w6KMu7BSsOYBaNAa34sGDcbNWQRag/T8a+E+uEVWJCZpmv2DZLSBlygqLYyTapF
JgkHeO5drUjTrc1xw0MhtR9cDlNxEFzECJF8SRkTSghd8AVPGR/C4YFp5bF6MdGLSzOxtec7pSAf
JAc6jayXjGHHdoClNyrZbvKe4adtCo4sjTcq4T9TEVDOnVr51j+vmNHKZmiu5UKfSWVpEM9TMEyX
iGj+0R3+NZS8zlgVCtIHXD1KBOkYRjuFZL+EUZhcDWJH48+TyLfTqrTVXR4V2umcr+xmh7Fpupf1
H7ZLYFYdSnMRsF+q6Uh+g44Qu1VXSqtgJUf5Se8DgHyW473GvFHxfdptlJro0uV1sQJy5rvQS0zN
/6QLC8amM/M+YV/VGy2ihEak5Km9KEwuawnQg7UhMz8BnCwpVo1o6NOpi0Nd++G2ayp+Wx+hXh+6
+vI9h0FexmuS4MJnNFb5N75cob7NSnLD2ujsVVNNBXP6Xddf3AV8t9x56GqmfMhmkpFkihNhmPpT
Bo9R0oNX/mQ3ITQ4AP/x5++zSRuDO5x3FLW1zTvRx4ZKvpzXzZAm2XX3HSpc6MDSs5/4XwVqY74E
pxKgOD10F4IRp54Iz6IYwhwILPYpZBLA8bv684QJ4BsQxDMvOxDezoRPFU1WqgHGMdiGAWCRYsOa
xFC8UQTgjep/m1+lZP72s5XI/b6bEuVdx2ODQM7NP6GZyE5WSLQH9csjfNp4DflkVj6B/id4tRdO
JVUdJ+4RSASIeEJWT80DNzVrCiNpJgWEpJpy8tRR61VBIPl1GeZAQFAmBp3Y4o486gG8qckdl3do
mK2SDOA9ei0P/8P3wnpk2U2UsSyZXDQ070/FHUy0Jns5Gzo+D382Zd0XcgtH3BRNP8+kmtbB7n2z
d+KbDlw6bivbZxQq9G94rR7anXup4ba38DDPIGAcKMGVoLUT1Bpj4LzgD5+rclXp4VslU97TwIbO
+Jsh06oqxhYzG72AiFO063VT7/jIaVR2zHLShRo0R1/q2jYhSzUGlC0poWDaUjFZxcAAU88uBdQq
UqZD5ZJgoaDHK0nlD6uucZc7Mo5+e/DFPnxYvaTyUmy9N0fVa75VVjVh971aaqVOGVpKT+RzD/kG
OIc0UdPL+v0GSSZd5DjDyGO3y+KSl/EIAV/UUaRTgDgO66T6DNDdQqvdWKG+5nB72A+g6HblXcwg
ICo9Ifz2y1nDSk36Frl/z2aNYbNGU4nY1PTsM/CCpID1/1qB6Hro2MiEOBLAjzpCjCyg3cJiE0AZ
TjQ12imMre9vgADb6oKwJXp/5Z5k0E6U7e1lgN2VwmqwYdQ6GeS82G682s7p/0Cvy7zgNETTvDdU
aule2BiPUquhMmoa2R8OdgMgHw5sDEBOsBFQQOdo2lUEkvgiAuwQLNm3VC//xFORwErCwVKHezLm
6q3arLc/s/PkpHEIYTm8el8S77R0NxuHoojJX0h5wXMywVeGoik8RTz2qETC5AjqxD1P34Hmz38m
4RCI99McKTOc0fWbPa7lp79wu1wWt51tS1jDSH7jvrB0YlxnKagoDhzLVoDNvF9UvKaJ0HQ7O+Xb
5fTT5MJReXtUoomNRtZrj6ZLSUp/f3wB2PgG4lcV2iIgT4PkolXrcikRif6aMPemBtLAMORNbpN/
ZID0z8wK8ET8FidqRM2hg7p45sP8mqsb1XEMLv87wnhzwLbJKId0kahy/bepmPwIQfJGWTrukLXG
6q+tmLYFQdasXDZkAbhpYSCPpDHu4VF2Zfgi1J2YoLiT7ORgOlZGmLuiW8FkCtIldNC4S6uv5qMZ
lBFCTBDNAFtWJfnxlo+6+YPKGuZGBsOVTud+rHRYlKsWfduF/PlXUQnDWVYEJRoig/Bcd/oR7McY
xc5XQMB2wrX1DVjwDtCsfZJ/D/RkM6OInNMt33Z0XBh2WYk9Jccw2LXV+SzNVuHO5nirKzyaU/nm
PfE+wlVbWYPNLTsxPfkbtq17srOLZZJOAStzKIDK0QqbHtw/SnHfZPbSR+cFHU8uT3RlbmVKJUHA
deHiyxcawZEaO9uVbuq8s4Ne3k9MBRwiCkslCbG0NzI1SbH0kd7UKeJ85iFfm8JHt+eDJSMa2N3A
bi57JhitwodhFGZxUw6eBjtlK4DnAZFbERW+igVjGcoYAM/yCMXRRIr9aIItAHLr98doJG7Fmnu9
ggW48AZgtAIlTcCfpUm+px3CGcEtjGnW8yY5pG3muU8mAqsuPrSdvidydY/UTIZIwNQLK3AD/4G3
VTZbxSdC4YWprEgCdkbHslHJ/KIxbbjbmZ4PtdKYcJbFLxUNwb0vWLgUBhkPUOGreM6ZD1uYNk+Z
KndRJfLGCj4fx0kPtS2Jh050Xnlmss+6PSSQirt5BW0HFR1co9Wz4bu4zLy4g9nqJx0RLLZNJhnN
uqItbSCTbcHCvf+eT/2Ny6GejG5CBnmtc9WMDC1BinwNPspUtvMMqtuFlvlsc03NsKZnwx4cjW4A
o33HG1f3bRfOWIbJpHOYSE+VRpGxEVko2mk9cfD5Fz2DBbZFLZjUeVLK9p9MHwRoBbAe8MWYiF08
ejtZ+NOcfkEkWPQPHnsRj+rz34c0hAzIvet4Jk7pe9ZQFSVaNkYYRJ8lSM+cCJk1guU3Ef/7N/01
R/BcKLQUgzS7YbomK4gsF6IQeyMrBDgBZhX95xRVUZxqHWLb31QTZCFDsHMQnFjk6FOp9+z83It0
BXGiwbbADPT1tPmKIBOxjOqYmsH04tb0HPzd5mOJhTdXQP6NuEb7f498Z5aDaUFrA3wYRugZ6XN4
HhxAdmY1fcBo6s3QlmRc+uiMXowtWQiL/bqlWcqfsW0nuNzz698XHyCsXU89ipWM5sWCDmV+Pl1C
yBYMshNC0FQb8bzgCHzYpKcxi5GcJd0OhBFIsudKwF+CWnHLFeyycaX9xmXH2915mVndzz8snVoE
Ib8dWrnJVs+GXVoN8ir9D93CNHLqR4Ao8JEiMy1lqznIpXUVvGr2V0lAw+jy22lzFEAJbwoQT2Di
8M7XCijg0xy8vVdsIhAN0EkBh60sE2V5TkhH4PejNFk+MF4/tilhN5zusKVPfMd91qb6jpMOs9Od
zT6yni2Z45eqjh3J7Wv/OAD46SPdzowhHc/vhs4+Wa5g2FJRLs+4uNQPtsIDQEFTcIDUCqTKL+ph
YKrEFBksx3FHVg6RDF8iH6P0iOHIDLjBrWBxfRRZEjZPxEUdoYD20jviRhz0oF1jeqfHlu6x58hM
Yna1WbnxFW9VawaJ8aJdq+4py3pLwBQV8cuqwp08zHvzdvOeYLWAbZSdwUE4gUqd8IJmoww7MINe
PZbS9GSbqplxNQUkJ2vI71hNGj7q3wdDEGZePNMBlCQJ5iOcnQgDfS4VLbZNdDFXvVJqftmlIH9T
STIAyGrDppaInpFxJI7xbvUTr1v0gpsI+lIDQz/WMilo325mxwl3QEJwf9Ro9l+aHzqIOfxE5vJz
40VA3WooZvYpCltfEA6k2ocDloIcvfcDjAMX3ndD8/o8dzAoBN+UWdnJqain5My2LnmdtHxTcdPQ
XpDtJhDOyqCSNUH3Zg5k/mCmgiRbF2oteLSaHbfhiPO+ubwjh4ifTe1v3RUYTxwE2hQVMc5JaEo0
kAw+8M6efTJN9ZlPKvXM9PMZ+NT+6nwypNZ0aoasoVSmcML8zwRX6ejAv0OP2w7v0PMMvC3A109f
IA9FW+Qh0O7GHXO+1om5JWJoLG7E7sxHf3VWVs3O7/hvFOSiMhMKAmPdyWWoqA46LpCMYfc/WasE
21Z2UAdN8qxV9nyxbY1FuSGhiV37ezv1chF8fnoJPGr/A72TvgqvcWabJwQltG8UUSo8qCW9MuSR
XpYiALt5x2gX6rc1vCzQCJJxW8N8WabZsWXTKmIb2sw8v7aeXC02AVqZK0x8ptLRi0NGsYhwwJzn
GRvv9odcI+BRcV+aCaCf1++fNSxZNco0MJ5rtHRL7dmvxr6xuaFaX1D/AKvh+/A14K105/MwRvQW
ZQ45fNxcEzqDjnrXb+cFgcctdxleJCewI1hKJeM1XcnfOz7UJyHhDUXW30tv+la/v9c0Gyop9yPE
3l8PBjhpKpmFYSjqL9Bnzr1XZe8+CoDNqbyhFWPeM2GAPPSf8UCzrm9pDQyKYFcfE04SJyy9aoAm
dFnzIfv9f8t96cIpTmba2ApWeJzBJdS108XEBXVMaBMcWUqywP9vSUXm1l4gV4f03TCwSXg3+ySx
UkMHd6S3ak1ZNAmi3b/qpj98C1VeB6vvdEmBLbRtvE2piSqVOz4z6JQx1hmJSLluh6JtkMk+jfnr
2hX3uu+98Sfi9O9llmwunsH3LQeVI+G1mYaO5Kp0Ism9TrjIPrwpxRsXzTXLk3Xwj07XvkkgRMh2
RMRUoG3h6gneYxT7vJEv2NUrXQJKdOtPm+wPb3bJxGQektUDm+FMQkH0Ddjfilv1sgbK1f5kGMjo
WrMwf3wFXLak3Y85xQyoSeGNA130or+UK20ZmMZ5WKXEYb0ssCyeGo/+0gynAI9+TBkNv81UOhCn
Ea+jcaZ7pDX7UK6T9BT2kkNSKseNTmu/TR9SP4XbpKbP2+HfqNI562zlzoknOjBDV8/uFFZ8izSf
qQa1L/drlVSdRL0BXMUC9QAbxHtj8SYMgBA2rX0vtE4R9fKgEBFY02IyYLWmoHVRX2+XXKDgyx21
zqlf9mbEJrVO11WFpZgUmI2MRYDnX2mXZL1QLYh0/G160WO0kdM4nFsahUegMAy6naXDcphS3HcR
xlY1lE9x8yUnszdSZqusYMFKbwaKhSAdIoWRP0SXyOsxo3mFM1nsKVRK77fMtWYCTR0i3XFk3yf8
e4IkLxbLmTV6cADLvIa3cE444i7Hwk9hP0YueyQ39CWn87iRSTSmEqHFApD1BmNILsGwOpBRiEYx
KCqOgclSH9ltY3nmSxcCjbdRANGWBi7qulhogozuhs0N/N3yrO9e/NK47eHSwIAFJTQp1WRg5D7i
7CEm7dw99ngnweQP+j7VFJALP0/ziYCUb1BWM1E+ByFH3dCxJOavbSxDswK88QwKqSAT0xrE8M0/
zuCGPyV8oi593GC1pprkO0bmgvvu0Nu/2SRtR4chaXnhAX7IqorhbWtkxdA9hQ2rhuiAWMa+PsR5
AlCGOd9Fovv1NfT8RVA+FdzvLCVOKbHObgj/A01L8PineTQZyi+1eObFU0EZuvXTzYda9ppjsjCx
86vw0+3iXzfqDpXK39VJTvYts5899ajdNi+02q0tpV500o1WWgOnKljgu8LG0Gwkn+LKGmIp50/K
raOol4DfX0/EPcjcC1NKeb7TeK4dZCpauMylOO6XV6xo5ZijTA3/SsndND1bMe0bFR0mXqs1M8mo
FkuifqGxc7yFdxC6EqxwL2cT+8xcMwShhERV8Eqy7R4qtUljBh/7qPk6p3BjtKHDGuDa1s8YgeRj
2rVEnlDPAsnhweiRaJNs7FfvEu0y4OvumjaI1p9nEXTH9M0rESpnZB8HfJDwLc0vBieQQY7lcpDT
NplsYYwdYNxzIPspBxQ4CV42a8dylLS0DdNyd49jKtalSqpk1V1EQh89N2VNF8DizzePhy8QBf0Q
LEoEwz2Woku9NJVM59xlUr+pqdkrLNL0I/ghtnAvhSrVEpzM0JxAN73qHQE13J1LriQasJeZ0t4S
rxoHQCo4jHAHitwKCsZPJhdpRlSaAaFjRzbFysKpDK/K3fIfyPuehvgsH4Ke9NeF/dyaj3EtkBBT
A3Nt+pKK83Sx2c9Cls97C+QMYHjsXNXkI1zWj4mKqRykoYMwMPNiRpnuKOvug0e6qIMQBlJkFhAH
zkEdm56XpnZggmqE7e9Rt6JtHvpfuJxFgzqEPt1yjM2CxPpTAX7GmaAM2IaLtqX5JaCvNU7q2amt
xGnQAhWkFRlha36Tm5RfvRbf0bpa0bz4K5l5/0+k1gbo6nyidJQwpO/7G/A/B2MiRc5r/ERVI9kF
ILvrBmwAmzsw36TcPCoT0hkwUea46Meur/+jhlLCS9pF+eplRZPeMFwg4DDJGzOjuNSW+dlIPFZF
F2uaoRdFupfzDUkFPThqSe5xmPug+yTcIskTj2JzUMn15WRKRuXUxA2nA4eqcBst4K20QfaJFZ33
wWbnE1EPeeL6fju8A3zsqEZLCdvHlV6LY6sANQOXFUSrDiiSsNWOaWt6Bmap8nZasi2Cfn7xXMuy
mWXb5aJ2yTEGH4OwmfSzU5ebpdkmYIaLJKCyFcAAEeni0ljioqm2wRnmGyduSNBSRfF3KUFyPUYT
vfpt5MNph0A9dIqNWCxZITODpURmZlCX3BFMvOEMbnsEvqjFjrvC1TwRDd6kH1EMZwOnN8/XX9uP
MyTkwB3fJ8vgv+6vxYagmM8T8b1BmtxAkNcvATnFgyPgJDwKlwFD0ZJQ8YhJZ1jrNBFDbT1JxB/y
j8THA+avIke/FKR+QAV4y+rI3VDAkwLXkByTBhvtl0+oRy+8NbNk1YWnsy3oH8ZOIVDEmrUOT78W
tCoHtij0XNVwbsPge7OxpZ3MsxEclODiwup0qJFinLyYajYu5EzqtlTBlmZBCSyXOrYt/XsKv+XX
c/U+VHG8Kc4qr0bnb3aPH9ljPixY0ltErIXcIzLWWJBay8472YHlUKcL+fWchYmKx6W4IYYx+SfA
ARhFaoBbx/5TORr8oFONknjalAKjpug+tgVmaY1JBtbDtdMnWzsvUuYhIyC8wKFD9buaiyZ5BV2m
ZPqkdEbum+OFhA88MClap4VOZrC73azvLEmcMiaO+dazf0XyM+jtGLnjLVymFQ0MYgEv3PLEWyU3
bbTYa3Re+wdriH9L2DkYutgav7U/QbMwRPWnFRI0bdR1do3DWke86kCZ5eduAHgEIjyeP2IbaJmN
BCo/cFkErvfnIFDh1UBZ7uHsKfr2y90tTVb/w3kK6rV2HN1vsoHogKAj0QS7OmgRZ6l5VGFy2toB
l0zBF2oz56OekfFUAxUTEO9P2NYGxpQov9VTqD1RuLvk45GL8wYyaLnJtk6/tOkm2c2ZNEVNwsG7
zKegTO7/Yp3L7ErwKCDjBEDFi363XdSMJsm/QYiJx/5VmqEUnJjQsRwyqf8O9ivEVmbN/Cup/pyG
CCTvT2WY4ha2GYxtIrRHB65mJN9HwM1kkL97mW/Fso6V5Zu5wgafDLQuZyDfkoFj2c+fpY6b2mPS
kuAydUzk4Dh4jllBA+toyBBTHcJRIhHAAZrAapRZ+Csp3tAuqMaJXP8ZauUaK9bGELFfQPQmindz
CmCz2ag9PlZwgpnE4TvSfoqu4sK43s9Twb2sFhYMJ3kXQBUOAL+UhTbAHTI55DNy46ZgSeq8cc9L
06KjbzbYW9BzUjS/J8hFF+65cFQiMkHms9KBe6QNfOi1Oe29c4vHaqbL4EhcWR9uzUoLu9dIU20i
iSegMvNMa7AGCkqVMvJvjN1hForCLGZBKnqILMQU26HTt7xcfhTiBuORQTWGpsvyg8vG/vKjq2pX
1OOaBWeKzCQn0AKKGdot6rK/sHtWfMlz+jBH/SOqwyBuyUz+8WPLOQBEWDYzfMbg
`pragma protect end_protected
