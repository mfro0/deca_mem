// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c+GJxUWqPNezB8yVxmmD+ConZS+ioLUu2eVAYHItV8Xzvrhjm4AHk8L+UjoEIa+S
z2AhrRqRIPVVFSIZGDdzYMExO7VB5wMQG77W67GcAAadjIepbCc6F5N7dQTV8NU+
5yjAUesZCWpTOW/iOteYDHFDkbVdQHyakmjgy7laZjA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 56688)
rSLdk/aJX7Lvvy4R7z68acZ59e/LQ8CatqaRxVHIIeDs8WyD3V4Ye6TldDlPW73O
DuK9yksPO2MVeRmIH9JlDukDw8Iwk1Ri1G/UmVXg0aj+GRmp5FIZTUsp8wCeYrO9
xBgPx9P3D7lyfIEP9EGPQdtyQdp+aEV7WjZchOF7J+Bq63CxLSPf/9NXJAEpRMQQ
rKRrBk5dffxtWQsEm2vzpZs0y8MCfhjKRpcERPg/sJNZGSVIFXjfFZiYpvyFpnFV
eBb1nbXce0o3HjYT3S1LzW7NzaDzUT8GM68V0JJ6CKJr35y4ZepYk69wZrVYbKC6
WUhoyaeH1vjJLAV2Ss9AiLGbnVbEdRsUhTlTGyQwt3WBhUP6kLNMiUJhNnsRvXFp
MgbgPJ587pdRnJYdT7x/enGkdpJbmvNEwKTnohjPnzt5nJ0hxBVimz3wFGeheKH1
0iiKa1xV2H3bnMmRxJ1ldO7jbszlSP0SgTugH7VX7OaBO7o0KA2nVSNohpec5fhG
dp0JcIT0G+nRTsz4QeLG7j3BJlWHDAHJTunLt5ZiDpwb52S5RoQ31f+u/F5bZpnD
jMDJErizPDc96WJPlJLQiTQzUx4phTXY4Lrwkw3zdFqGxMcuSWPO/u8FvLJCPMSq
/2g5g3j6vkCDEysvnf/fLRXqQoQtrRTKIL/zWdrXy2FeOnLSBvNA6D5g/84aGlOF
VEX+YcVubxSF6rauQoXcJNb+IBlVT4SDdHk3Jjb4uVhq6rYJqI6FFkZLhNVZYvWa
4rNIh+DKxTZGaen0QVDuh4V0ZpmhE9WQAcYbtCir6DYAzxJ4q83PH7bEt+qt+K72
5+oDFijLEAZj25d8qn/EJTVUWLbXzZaGUzkU7aMl+di343eQ/XGZU5SbLkvNgQok
WShmPCtIOkLhqn/yK6Tdd9qmLEhRcsY3dVUcZaByP0eTCjU6DqhPPLrQOn5UqQac
8uHhXdjT9zKE6nOQJ8rK0FvPSEAnpKn+IJPbqQfzK836eAMAAOSZATg53WcB/ZJB
DlFJe93QB1vrTs1yNlrJAiGIZpcSW3xBnE4o942ozD/3b3rPAwdiijTEEGJyra/X
h2bQStT02XjodZ1UbbnF2qBJbek+EF4XzLTxSqEdjzZMBIplRbPIVf2fWIf2p0rD
S69YR/2QvEVNTOUdaWUrXFri7JoVc/qOE0slDshpOB2eOrhtdSYkhFU1Bfb49WHv
MOxlmhSmBHOvSjst2BEzOnMVAC6Ys8yaqN525VU0BpdwxJXc+9kcZtYYIE/XLY/n
7WdnEj4lObG//obSXv62IzO4qq0jHXjc4mScdInGsdLkX8D1ATBFRgIg9tDzaZm7
Yx3EDCw4da6cEt+7J86hoia3+aYqd+D1oTdUlFWXkNQX1Twkkt4hCKAQ7QnmgJxH
9DWknA8xr+wVjdREvWg34lzfiX9vtJZN/ijfL0i5p6sEnEbShh9HarOuXLPeRlav
v3kT05yomjpUjx29paxR1oaPp8jQi2qFc/EeD5Zwhsi5aSrYIwKtyEfY369PSSgd
+wY0auXoCNENnwcfUgWMDvloPtciNftSr+Wor3agP+IkzLNjNsf1AqYw8/xv45QJ
HE2ZQnPhdJMTECfqtvZgURZAwb8skCB0xdG8WkIHgt77nyLUldMPjVRi8MRRARJ0
H0lnq2Jb5CB/7LYbl7UtgITlKj/08rO0j7fv0VI2CZG3/YnCZMAtZC0eMgPw3HfD
M1quSYMAp+mX3uRtgxB3oeZyPfc7zkTQdU6NGxZMi40dL7GlejDUSlRIcCGEAG5G
2JePsisbxuTPkdeSSWV15b4Z2UnGaHTJDCiuc7Bxr3RI6k5TzMT8VD0kMIIXChts
EwLIaIJDyehIwvJcvWzTRLNyZDNdnlYP4pbjI46XRKZvUhf9G+f14aCd2TAU9Ox7
vpH4R2Hc+Vd4z3b2T6TUJc+UHitZOTwWTC2YMUDXMv9OuHSwPbq58xXbv0r85+PU
wcUZUFxKcz39WHKxc9GQfVewT7RjYlZ78mUC2l1xKblXYl6uI874cj+YvUsmrH97
+Q1oVUIqz6bZD4cSRgNhGaxpoPZkrwn8jFLOviDo3xlMcvqGI8DoE4rpsTOynh92
PBX4MkpM3fLl/dJfY8AY3J+LGg3Hc7aYCAjHbqfvFEnyb5GDpgk7HBtJI0CETRNh
m3Lf0I1HhNUfzt1IFifVxAeUY1xmQ6C4AZScweL7FBRkmgoAux8sUZgMcf76RyiG
V9nIUBtDZJkZ9zUIoEneH7Qli7kjMNfV0yLrWi/GG8xRTEJby8o15GO+5vfBYntN
2sguAsfS3qr9Ems3erfgzD/e75GR6f+k0kea4/FlYEQ3gajH1fd8kx21QqZX3/Du
sELDL8Qr2lhNlYAOZcl6Gybi+9Yow4PXgdiWbDbHKEVI/28M+waxXshLoreuvKaY
NKeZAn3cR7CLcgbZ6faM74wM6RGIsNmZwRZNd17glELiNQ6H/gkjdhSdSLRI/2i0
YbM45Ugk9z61wyCCNgrQ1cgVjg4gH1cY+tGW8CBIy+O3vldeKOLAmaLFuCCw0ILX
fDo0L98A9e3GwJybt2EvTCbJ1EKzOYoeYFoOzk8UVUCUtILm+V2lBe5ChyEdBk3f
JuqcD/hyTyV/LsC49yzOdmATf71gMkBuL6cqeBXh97KgUbjBJr9ulDcZdkM7s1+1
yfTCDFiUn1tnZC23aa5Ba+9LfmhfGrFRYKPrIh3+a/EkI2B+Rn71NAhrg89MJSLY
MqmwJwH7NSlcw3z9QRjk6cQZjOFvA8n/eZq/d1bMj5laJXenvSLGYXd3DedU231r
8fAohdPM8hQwHqTLlMv3ZUC9pyOXskGmjWoTqyjSWSFkd1AQVN9EHrbS1xtLaR65
3Pwn5HeMDQ+BmFDDGERhPUvIegRFYy8E6naXpaSqIn4fJrY8Nuc9unim6DGHmzjd
RNHBptoxw3/My9Im5radvAHc15DzOhKyX1zhzVsuVkD8o99m51YTgFVOaDML3dhk
lua6SAffwocTUeF2CXEXRnEXC4hFPVZi6Q5gfyHjan5c4o+yoyM6fTPQGTqNKyRM
SgZvlBdjjcl9NFZf9YYgJQT9GR1841ftsWgswYBJAhs01hkbX9dLJlDUcC38Akx8
gS/tC4TZxnDPirPRj+6PewBfVMlAAtj1dua7pOQjFltO+dms1f6Gpky3Qz41uBHn
RJRo9reOr/SKZ3gcnmkT4PXRxr4KqH1caQ/iuomJ/2aIRX6D3qdidGXT0WH0yYHA
TOpXHffejm8j+oFg7NaaHlw2rCeHTZRuXR17f8x+NSG9B2j6t3cbOEkoMDEN00Qt
CU8ReShMrhmoQhj4ppQ/JyTlkdarwifaSdJJuU3yeDhmcCPX31EI+8PjfgRTpLTR
yfha3kf7SgeWlpn8ZRJS/mnFkqUd3XVQ82qb/QCpAUeUo/JTXRSBqLNEthn7eMNs
IAUsn1um+WFuyBRn0K+5lpQDtTQ39n4N0WGQZ6iNN6Mp1gBOAMyhs8faLMWpN//s
/kGqfyUy+6Lj79HtuRRw0ixgLxPjAH7DEGR3BjxLHYKWMsXKAl1cbk+VgzKsnGdq
pSMp+0k3ncUdY9EEXp050zYQ6cEl46rksuMYvgUvBkE8UNKrpH2/uuodDA1gRZnQ
/HmS9u1AZFZwLNkNxVXyaLDI0RvM8HVZIWFx6Br1Txt151U2lZw4AfH07RFRMc9s
7CCLw6N5EIFZfCJiHvnbBXONwSxE4bsPNUnK6+oui5QrgjoSeY3FVUhbfpGwGGdf
aLmiDKqFWul+Stzem/pShk/20h9CYSQJRXYTdXNm20TWJ2Xf+cNIQ0tE9klEZfkv
lCT++49lKld6ZoCDK8qtNIU5MJ656Th2QmwC9F2rm1ZZZFCamhYa0xLAZ7pEE7rn
SLG+NWeKoJTSMUzCRf61Vc0bv6IYUPZAX4J0X4A4aRyJlLFtpcsRaRUbWAYqBqUs
m4/mb3iy5asXoKd2X74LxYN6gEYAodNBmqZpi8pmG+Z3xr3bQZKwJoq9mh++V9Sv
lNPU4XmlSeujd5uvupJ+fW3JsbIFuW4bzn8fKyRorabqbrtyfdp14AR6cMujZqZ9
cy8RfdefiRXp8oFarsoKBJci4h2YvavflTSa/A08SXRpMSddvXn8Ig8uM9M8nieo
PXrkA4fAMk3NQYMJf+nHPvMxuSx/bgPfygfRreFkd+xzku9fbmwX5//Cjjo4pVio
7IQt3valv62RvwJoJJCJ8l73XStbWGOTNiKXSx2Ak2x7l6JOuzrF4EErlzR8Yf/f
Xu4PFfmG4Pi4Pga34q0//wq9BUZm5Fv/SJB3pr7hFLsteUqRacOHr/KPWGhMJs6S
ry2GkvDsRLjuliXxZK8+70MdsD1zkIbiJvw9OVyYs3H7bAiJSrcFyUx220OUzSTy
BF3zsCK6dBUKdSezOkhmZdhpnIXb6IniJEjsWSnrlBwIh4JpPGu9E3xbWICY0S0R
IDt0I9GytRVPrxFmKJvrUN7Qc9LdK8HfBjNunIQSdrfdlgbvoFM2pQU9tjnwHSIi
npNeEmV5vvjAGBt9TmI4Iy2JqEfLRU+jBBCjz2b5PiaUu/Oby5UV7PXvu0x8phgy
awEddgcqE9J+wv6ymTOfDc60VJX53VVUzn03dk2xYKYdc59rwqPHcg99WYpAJJ+x
ey9zi+dap+hiqCif//imQMWxRbRxjKTZ2kahZmX5EqDLb8trKGutgtwFWG/M5Ghp
0ersraqr6y+Iaai25FzpDMacAyvCOyDH5rJigo2l58wpW1yO4rtT5iFiN9WzvA6H
WSvW+jgJ4IIGfCRkvccgnPKF+HmdWEQs2u9gHq88w3/+24GGOp/yrsdRbMro7ldx
op+eBKmKgSqy5PN8/89Odn2MlNRLStvuO1G3wqrkvjxfPV6CMFio4nvw2ay1O0pN
9DsiVcSkZjuy0e4BdiNotdIE6rjqVVwWcEY3GKWz9iQLDUSldoLDEtbyAa+Vfuts
TkN61rVl6KjlmEZL6Nb5DANcrZIocYrCqj4YrHVNw6N8Ah2dnOeniABLxAtUjTBQ
VS7O9Dg2Sk4YZaJYSdE+OzWNDVfmLWRiK2zncDfY5+cQF6KrqFE8FHEktI/AQNBY
j3fzvo60W78f48xZwLNwYVGrpbw2z23l91SKPAF1O5ezc1wd0TuiSzRQLzGe/Ifb
wSKT94vjpDBYycW6hpAqdbF4LBaKJCT3zVYzFYxVc6U/pYjUiF96gvXrlX0HxRhf
TvzIrZ55Fm3JrYxN/wHNDDKPfcKFVAG/mcaMSt4RayeMhR9KoRYjqDuVCfOpuMJr
7YyB6WH+wqpS4vr3Ocrr6wqbOuw151mMH5aL87pLxjOKy4IC2bm+NrZ9UAmFIYr6
9T3Kqwkrq7vwEOpQzi+/eYQFEwM8iU/mEw+Px9R5a3OiI9+XgMy5UHVF+mPL1hhr
0HgL5fs5NCBiGJWj4Xdpnz8ERvGYtbiWB+157zKoNckxehvdX8peyl57wqHwnOPi
OBwQsYQYa+fJk+FfiuZOJ+dwEPQdrG0haSgnu2pz08Gxe02MPMPrU13WlufNMc0r
5+TQGKRFJTHsYb2TJ7lGZNyssJ6wS8fkCP+FCyzTEr7XBbHF6/LH8IjKFIe/bBdo
huCYPHAYfxoOAcop5IjWsoI7NfsvCjgQjEjipyeatHc0ioVTfuxMxRQp/4Pg5o2C
8Yy8WXT9mVR4WUSLsuQi/R/Q3Valuc0Ay14iwnySZYSoPuxbb4NwkeufW1Jh3ATb
/Qd5NfE/qYSp79shurWFMcC7KkD3Fy+ArdwveCYJCMMlm0nD6nqloMGSJSGdHD1s
SBB16YaVm/vCHdNV1NnWmQMMkvFgilkNnKoJYD4mROB0Z/Ttf2rErOBi/6cbzZ/p
KqYw/wp7AFIBQNBfMELDpI7wXWvW1Tg00JbI/A1oG2XYmainTr0Dnte8zjolALCQ
3Jfmr/QCefSehzZVeqNvuQPXgujoNVqdFXkDWAJVq+YF2xr32EwrWShLpHXC/SGV
a3loqy6uTg0KJNtUyQx8jScdckJzD/G9mFh4dydWuNexTfAFSWfV6FcX2n3Stp+R
CGB0FP9sDI3vCl1B09RuuFzMLabEPIKHxUWIXvxy9rRAWi2ueK/JMYGzKCLdb3RF
QgVuz3KIEklQaZE7jnZDeuYHP1ghvi+gPLZtmIotYYMLsfSTkU6Hg8Fmb+HUbzDr
4ElIAArLWjxobX2s80MuncWCqjbnpgiR8IETrXozjs6s2whmqtaDFI9ggfKb/Yru
nouGCd1lJ0WX2kpIuK5pBZIMaX/7EBVAiOVcfP6QCR6gFWZNpjcugYUSeB958RQv
DGCIertp1fI7PpQ+sd5bAeLor5J9Q4WMbu7puY5860LxLU1cWmA7myHXidKG3UMV
FRnkBHwad5TyMY+bn8yGcpGKH6PMHiPNmCxx9EkHwhquenjM0Cj2ZHMtAuQApyxS
eAkaUxfG2+9QLAr78shVq4VAmzB6T44GW3psoJEcPFLpPWNvBuBQj6opp60ScsUj
vj5cp6Cp01AT1WrDk9L+As0EsK4Ik/lPOE0VDvCdY8GEvxExvnT3fOmBogHwKMh4
GtEB5QDK8TCF0FCdUvX/3y+Vq3kerVTGVpY8uesxwJ+lwLPTz0SsbUJF6Q855HTo
D1x1dBo7/DnsfHlV+aO3XfbpoCvtdwfjMDFg5qgoUK30lMnIItCFaXrrwqew8flK
YeceuEfMgl5Avtqcq+2ls0ElVH/CrXz5WGd693eiH0nBgGrPTretN0hqYXys2jgq
ATnUei3Eh5uiZxf3VRmuFRq9JfqSdFWHqKslo0TK42DpUEZESgoXfFYg9UKYdu6j
jCeOd/+CmxeFGOllZji2DY6a7dAORiSuBECmPcWyvrXaWZDwpzlhpRlW14lqMKMu
tF0stEDeMc/o9Pc9DEf/98CZ/KlthpzjRdqWhbujuf2eurm8VnmW1nvImtv2icye
HgG51zI7ejPMY98GPI5fG5JX9mCuqxHY/Q2hBZk19+tnhCojsKfoJ+hgxKqZdJH1
fcu89DpDCyrHfHWdBgD/ESrPzvvarsEPzJIcbj9poemfs8y2ZMYQfq4PG3+Kzfmg
ym1/6rvvLwPootNtL3q7lIZ1w6KiKsLt/sQflrYAj3+tRzrz/zR8TFL+yQeDRSkz
TC4+IXOo/e9MlkpBBgV9XQQuWdBNfwAdTnr215y5wnHtgbolA2QG2ONW0k9LT+qL
i36QMfu2VKckL0UKZl5XZixKFBwL4oxDh9MYzd6phpNJsq1fVf0LbhjMhJj8A6pM
OfLdKeNYFfGp2asGYmnjFEeeuY2LbpCupGUhwtcwUqt7h7/ubEUJYGyBldd3EFGe
rbCdsYROnYaxXoJg6G6nGGmUD9449rZBrWFmwloucD4EDRnDR9UhekqIas3JMa76
hRtMkZ7kxbnKGxz0VJ4DEItMbipl3LgTvyAsFiazg6zvR+KiapvAZkKLbT41JSB0
+8LTs+VFcv7fEuSVgQz1WtSdt2ZbylbbSG6Ld/uNOLqZzMoEDza3lyiYwrEqLg8e
mlc9rsSClezG75Cau/XFVEZzZ2r00kLHViL5hGJ8LI/ogFIuKAqvtXfcTpNlNwtB
HzhuR1lgXvz0cE1jjT6F68/0zZP2vcC+SM7E4V5aMUH7Ct+Ov6lJbwz3BUll0axs
1JZBZjh6kKDBBONPPt5QzL2RfMDZuqjJidgDNjr4HisSVIE5G7f/bj6g0KNj/umh
uNkgbfrQMZT9W6q7oRS89rLc7QvG99yyxGMv3L9BLF6qqOYOYaNPhpS1dx6r5jVg
ZFm9MtY0U263PTtPH7+tlsKT0Q93gJPofbt12MqkFdygnriPzMB6n3Ho3gC+L3kA
3rIPuIYyEvaqqET0RZzQUotGIMHK+yM0o00XGAtnD423L9WqflGlR8xt8lzTJXLm
SYm8mkzJ2QwIRfr7CL52Qhl3tjelRZiVCeWwNhFCQSwTPRn6QuZ4oevec+QYFgkr
lb4bNj+SqDErdlnVnamzZfN7POLOp52XOdKsksAmdT+OPU8mhoTPgm6+qRKYtg59
V3cwNA4tU4BHu0+G1as2jDzQjb4OGUXO1GfcWIy9GTala6Fr8bMzF7E/dRapoIIL
Y2J7+uZKnGtRtzQSUljTDsfFB8PrdLff4JYNk3hWufEOJCOKs0DJOpt5kDFSn4Do
zNPxVPMj8cycI69XdpqccPRuJplvs/0WZMA/jPKK54QPy7eeYGPsQwvXQppkTIAl
iVyvA1uR50Q9Uxppm2LboHzCCdeMHGxOqb8qbrBIVWrasedTaT88w4EfqT4qUrtt
MIaaoa/cnXi/GBLktiDdGER+gwb8co7nlITVMOXTd5e1ki/1qRhLQm0o83h3kANb
oanBRfWV2AkSelbAKlk+5UvYHAIQTVSZ2Ayk7dlt7wo/xId184Ho1ypJtQXUn4os
ML6V8KZ9tt/Ndll5qu4Ajv06WGFqQQfquGJ1+rwWcKEDyR6u40mA6aIfXA8mmH08
+UxQC5Jxl0nGhFdiDl5ts45Phenfk6ytN8ySId9cjSfLr4Q/BPg0x8sLANmd/DCn
YIg+hyZ/Yd2YHxvSD6R8y2G6BgAMnFaMM/mDyUtRrafgb3V8oF3TsmBY9aeq6b13
Z3+JLesB5FqqSI/nF3sD+gG6XToauRnE/lMdewG/NF7t7awT/aMpwuoEM9BjG1q7
kED5KE7gTFOYAgyYEVUuQO8xcoBjQrTkdk66d5O1Zm99JzzNkRmtFfB51Pr+AKj2
G5pbHRAEa/tnyou8e75Kf4jZqgzs3waUGd/5lO5et4C82vllx+ZynNCFf7qMz/+0
zJFg9VJyVlZeJAtCD92zXIcB8i0Ctkg+Dzv4J8JxSnmbFPjpz81ex6TNo+lv/8ps
9BueiCPAIqzTyTmPpyd2w/ht7P+4AcpQ/jmJTh80yeLwdZXHg/hs7abZSSgTCRkG
9MJCmFuMlWUFDRZDVqiVFthDWgK6hRKDj5Czh2Zh9gvhgX66gP/2Ov6FdC+7b/qc
nQ5gc7hoF8in4JWOIi7BvNe9qZmRifZwag1awOQpwM+NO8Ne3SelDLRxgZHRaY+d
/xLZ7oaK8zbZk+MJgNsCAWw+ugmH1BH5dbCbq1/rDoH2+JtB0J3aPVuscvNAUNam
kN36/FsW1LiO0jbEXH/N6YUSmPsm8r40TKg41xByydnERL0G1eRsU6yYgqR3xcvG
3mWiOr/OUuByajkpN/YtbYFXrEF/UQFdj+C/3Aov2phQbm7o2dkF9cSlBQa/lnoB
m7RWmQMtgI1rIwNEWyY8cynbLtoJDqZ5tm4plCprhaW1/HEAlvPkuZDFRATgm7GF
ZekGO2+YV3+51pEJn2M+CdDSA1r9hkP/MpiUEeARrBCSh610/rEbuAXoCQkpuJEI
uf7waZDnAHOhRpQB77NxqyOhYPeOg0lTxLWOl2f6w0D6XQ5Brg2ccSzcRVukm8Fd
emc3i+4CPEshOltbNPwyeuLqjy2ipd9enYTPwykBulu7gqe4F9kYt346bHykXwVs
JXmYaOpliXY09hjffOdbPCB3IN/SHSjbUHtFPVboIMpO2N9wdFKU/7Yttq8Sdtzh
ih/lI1UJxWv5+sextmzO4SNQ4b6z27XSkVGT7COucXXiBMfrcBoOHeXG41VIdZO9
gwj0cGAjLNmLsGbjMaoY54wKHlmOQ6HYQIVdIqAHrsOoy4nebw8CEorOWOANjlUK
O1IT6hZxbk72b+KGHaiEUFTsUDpMXv7aARx/3tR54refAz6LYgo9UGlWYKLExhxA
ZH1QJm8Q0Ug45NKDJeC5YY7Iy4JXit972FzpQmKVoYu1/vuLPl7GxsRnJdl4Z5r+
/LqxTGIuTXFWHLiAk/X32WXw2uRAixVOWbprNuAubv8vylJYIIDa5/7FLO90MblA
OV3FtrV3mJi/SDCKIUF4DM0MtspCzZEAHzSYc09iim4N1FelTHQQ346m0XMxoLVd
boSEZyXG8t4qXmZvdGTqqqXaYo63Sw52HR6cRDMNCewrVBm9vjyVOn1K2xzXOEu4
UwWY+2+sp026Zsy/JVCCBI+WhEWGFyVJZqcV6XjgJsgZLb9ToqF15ipwBjza+y/v
I8xaNOClhUax99xUgcRWFBT5KdHpt7ZRBjIbv0U0976jS8RkC2Ittx070GnK+WJD
vMfjlQWBRlbEGdBYrb77geJnKac/0si9Avpbp/k/gWh6Vl3Up8ObaW2QLX7R5Nnh
FqxQi7W4V9wrx5D/smagy2n7qjpmN3tYLn4wARgQ70mGtv6ze8RUuQGmvdssZqZW
sXszfuvkIsnNyzI3b0f/GR9O189XG8NUwJcOSyD9eohF1JVZkZ5z1Y4N7cpQUytF
9LAtD0QXIaO/egjgLqcEAdXE/ExpHXCNvY16UNk9q/ORsVGnZQkQvQs7tcwtyEsF
hlw4OlGC2aRGG2svVff8VsiAy3mA495K1woDIUdHb+z0/bsvhGYf7uLmTjnHJEBS
givNNj6webtOI2YSws7WnEtEtQ7kYI/Tl3wv6ovReT87XhzIHD7U5qy7rsX5flJ9
LfbtES+Ai8/lgktvJb1V+k58ep0WHvEhkg76rpOHWdgWhtuIUNPJ8GTnYELR4/ml
geEskkR/OXZaVGBFd8F0IHrznL0uaoR76ake9WqVI4U2Vspw/Et4Xn93Ka8NM0fN
H+2H4kHnGwcd/IWTTLfEsX+JLS/sOgfOzW8SetXNqdcUZBkPuycwr2i77ClEZ6By
fjUUiLQ/bLbfe7p4eM9AVY1rhE1vaEbtSsP90DWCKAY70pcsxRmIcYgxz4BWsBn+
SE1mRirluwN4GIpOveRmJ7HPAWX2PpK70XAPeAyAbS80X8ELoxjSXjdmJffN/MgB
oCfEJbFPCDTRPkhb6ZAQMnKajccohlQ+ds3SLk0tjezQAzYU0BMzkBoGxD5FceYO
+vQ4av6ao/lbXTSQuIjtEWMUiaZbnmZxeLH3hetWIlODsDM2wwLA45EjLL68vVMD
mbs/a+wfeg5HxCGklkO1aDMPkhwFAOy9F59TsYE9DVEdybOuBkSoLHS6YHKMoPbB
owseOn0VpOFmaUnZg2U646FMcqn4i8C/VwVUfVLISLfi2UesM1iI4tnVyJJ7xzbG
mEygiuXBaEbhO+3eqIKorg4rBpZG6fOq4bNTg6QF4pEIbZSDcIvRK9D6gIzzYist
G4viA3TblHb6x1AQPgWHsEsAsK9mbKCtKYNyYYooEZ4eusOaTjsUzV5Lp+pttWKV
1LvpQhJ9CTVhUL/Nf2ke+BVtx2EqQsVGBHYWhV/XzFhE9e59fL/QvNKTKaIsNpUO
+n+z1MABHjMC9Fe978wuZMM8ftxF1ZQh3UC8VJ4FOmsmb0/44erHzX6eZkpWV1Pp
qq6m4wQ7dlxLRUX/pFRvVqj+Y0T9p8kA9Xni/wFPBEzAKDsrPWUEtkcDU1SeWeee
9MTFXfpAzjSV5rUWNVrMCYPMCQXfX65iLYE500TJxSqEMIsqJ2BQk4SFvqG5XNbA
DaPNSaPPFvzjf12mSfR4uWN23Kb4Mg8z65bQXQkCRzLerSuHpleYIHzw8qMnHnsR
PO7toFZPjdSb9dnUXaaaOT3BrOHvtVW4nBnSmnFL+S4XkthGtLWu6tVhPp39ftN5
kQYOwBTz/V2JvjKSgnVPEqZVdHwQGxyFyMOR5KQcBbr4DQaUvBaMNaZkaQvxxITK
HLhy37C5Qy15rMULtIjMwHqO0mNkN3XLRo/tqFWXNGcUh8n/tFRcOoYTLI1KuAjs
dvZtTU6u2623Xs4hFUCd8Q5HSqAr/Z55po4gu7zz0zEEik3Q83mB8ftWTHyQ4Vc+
3sl/FwMYKL+zqtyEn7IVeeph+GquW81EBqZ4/c39zBKB86LcVs1WssS9KZ6XaJ7l
6ysh6h4xSvvd0Owzl+irDYbP077pfgc9YWlB+VWjkLtHxVdgbcCWLUHUov6HESxp
hncJ3rXcKu9Em6dHSsf1ZrGgV2XgMNfXp8Aig8POKkUtq/Mwfk9YZ9Ju8KGeZjlR
DBoy5UqYwVnr4x00iiIQXt+/PaRDqXNd3Zy7J+b+stAQItdZzlqf8rzxKRQc2jXt
d/tPeRGI8B6Pl5zrLvjefJmglNlIvrvUmXCpIw7BKtDxbsp7Ot4uYGVliZEi5pCZ
m4L8dTSA8ceJypKCXzQuLQzRA1dg+lKR2iPGfsaJm51NMNiRZdEmbQFk265eMx5k
hfJ984GbGMkfmWYaMIun5U1TRvi2485QZtJ0YQ822UIylQKfCgHbVUPqg2COU/IQ
51fjy61k0M2TQY5IgNXYYwtghwAPivM8bxSTBUJArEIQwjlTus6uTu2busdO+Wt4
Ttbg3y85A3JpIm3MAiVnTuWEITARGjWWnlDfJktANc6McRMJf9+yG8fDeRb0AONN
TcbRENUzsqzqyYkc86XjQtJflue/Mbqoh1LoDuayC4RvgswhwzmUuA3By37/G+tk
GB3N+vIqbbodN89Sr9JJG86gkMyWdkKPuMEyrZtM5MXsA9viUgOfh/gOBm9ggle0
fwh2Ww3IU9eV1aQWuH4tyPB9BBw+5/6b/51dOZcadC8YsWSuSJZRZZdReoJXyA0G
MZE3syTVWoV7owiyd2YnhR7aa3EeI0HDBxDTKE6PK/DKkmGmlYUCAWKVEJIGjPkX
xjJGXxqhyukeV23ZhqSAPzQGOYTA2rvDoPIoAmKF6ukxF1abmNoPPAYRufB0aOIG
Bk7PNDXXc6DWiQAG6geS9dKtjtQy7Q0kW4WdfD8Fb2yaccgGKm1ieXu/SM6JTO+d
uXxiBXLh6Pb39r9JJtyfPx0hsS0+XuktapJ/pz08beh/mWOttDlcrQmrhiDoxT5L
z9eZIxUiJ7xSoWXq+nZzDTsv70roP56CUo5P9ZYCOX+X0Y5luSpPPaz/vpGP/suq
gsr+7xH6YdIrjDZlXIu/Z92OtqhmZzPjxHvPFyQbzRp7y/bNWiWNmVI56h4w3eRe
XCmopV3X2yxML5aztEKTqYU6CkUIx3FTxMLIXtkb79PxSSDrtKtV8UYZifs4fd+u
HT7Qm2l8Xl70p5RPljxAMXr7RvUi3/7cOzuWKUXscOINBy/NXFTKrn8GeN/Nuo9Z
3gc2LYPEXYbGSLCAy6TbtG9JMGOLJDG+eBN4Jxhf2Yue1XxOEkYz3i5zyIPUwgnL
7HSIKGF/jpm0YYIv8qH+u6UjGXta8neWqZ7rVWSZYVwc0gddYmOZdXOiONKQ6bC9
Jg+mZ0B6UGoviKp2WSagYt5R7xo/DuqueEz68KYoqmr/jgy2Oa9/IXdLtJ7SUheb
w6cNmoQUYv+oLisWmEWh9Lw410hgqzPBkl2xjYX40ej2ex9cWPeFtFxjLtV2SeEN
iRrTxfHC+L3pT7cUKwwSxa2EiG9u+xvUVTXF1eXYgMnC0NhuVn6jMEqAr96lUPU0
GIx7stPmgPrumS3vrtimhTw93w36R6dfdcsCJRH7aWZ4S2INx0bCIyzGsOWyzJqO
bIt5n8G6EyBCThEB2MBBM1UUvc6DzSMpzsioDHOBXZ8mwcg+twLS/M5aQAbszjXD
1GOb5LP56mlYj+X5QPnlvJz2t2xcx6G8c+az3UbGVEbWd+7AGooNsUiq5J3zaLWP
Wt4t2i0KF5XXD9Dojm5anDjYWZp2gSiVHDNJptPrOuOm3PwA0xYKXi8B2Yv5TXnK
d/QjB3XHXvZuQpelDc7tc8ZIZRsWwEUcquOZg5p6D6Jbr1l+/UojEnixInsZE5Ja
4h4WMTWVitSt3ymLdgeMm0mpucRJD0JCia+dJQhk0ACI+8jQGYIpomOL3FS2bDnw
HO5M6DjO3372qV+cafonbQJ5IOupIz46c6c5jfq2GYSxWwRJsmIVk3P+Uz0F4vju
1JW8bZBPx6xMblWtjBG132yJQ+nAXhELs9kzXCtPnypfjgwSqkQvnFET319Q2g5X
usZMn6l+OzbK9iCvMe9BtuhCwee8DlixJHOZB9qrzLGOy48WI/tLhYO48tBybwB1
YWpNYHQGkc21dePJp27JpO95T7rSoJW7Hus07jCi/iLMZBXmzeBmUcklWtEliJZW
L3c02VmXaY4P6v+sujwGka3FgYRnFbF0Jrn8UXnx3pylSanN+ZBSR9SmKr+J2owH
UFOsa1ZqYWoaNSFPsArhkMQYOg1TYPMJnLTnYR8QN+aqUkNxn5mK/evOYgKI7eX5
OFK0A2E99vB+HKNWbgwuJypsLqWtEHLCmVw9lby+syDFdXOLQJlO/di6DoE3TWgZ
T5FaLBDE59Jb2YWEPPHxRoODnEV+PwMKPBhUd2659LZ/I8HQKHnVXymI2QII/RJC
vZ50D8iI44aff7akNm0Sn/8qzfICHTyexrtX3IMDKY9JTGSEw7gI1IttJVKRyjuH
lBbyksDbqOVssdfE6JMu45dXtcWE8wRaDhBWfLXKt+q0BX105mLh1N9m46nh5P3F
nmK4CVOnsMMp6oSw6B3I9Pjo19MGiZXEHkrl7Uu/rsFjXIqrzcVEfVn7lByOahmc
DXk6WPXWqYy5ujXCein8v1hamQqXKqsQaj9RGq4aB9IM4pdnndfY6JNysMv4zAbl
jAX8mHuJAZNk3c9qUAssXhlFmq/zvcjttLLScqK9Qxkqg8KhiUboUCXPsMtNT8AP
w5b6Pcn38//626xGklcd5DKaVaYeKmoW8OUOaNQqs2z3EMSo5lKoiYIGW/B8NAOC
QWrUoYk/3x+vNbj+mMwYGy68vuddwg7WsGUuFuDYIrZKn7gj8iaCWzwS9Q7L4gxt
lIfD8/f0Xj8I5ZRtXB/67TdMz51gDB3TtQFZ5LtKw+ah/5ovKg6ahvCx5y/e875D
Abo+pzwogeywFpY1J+9vPbsOzbBo3usoMzTcSOBHnvlDwKIUX1K6pUh6uybToRTg
oMiiFkYMc6FdqeyMbl/CHpaBReaJx1p2NHsaT7YPcsfg/yLJDww9xQ5gTLL2SMvq
pd6WvL2ojhWVNvdc+kYsin+1YqNsOscfsEOrftiWlre+WoFaYsJ6JvjWgp0abfeA
tRRn98OcLKE9UcHJJCBV22SBNTuC+P0Lgbjqb8LGO7BaMzNzxHhWcQOJlXGmIvLp
fiOjt19HV/zDl6/Eb3aub20LKIJm4i9bMzoDoaDX6tAdy+z2O08aD9ZStvndnnTj
7jGOj1zMfr51Gt0oRRMFl9JQDQH3jmKOPXx5TYfeTj/WpslNR6bDN8AXDX8bAPk7
t4BBDgBUHCAgyNv3ZpV8BDY9e1laoQYDFthuXWEFLEemGkIfXfChNSBDQZIRBewL
E/hARdLOnxeo/1F7CiPGv9btXhzqFmrhLY2zLPMtO/Dyb8cj/hS1rh554rteXwnO
uGL0zUtOzkup8z+XOXSOrTnoDSBnPzD7B8Nc4b2B0pgEClEjTUov6C7Cf07RiZX5
CNY6kUDWyAnMbywq31bdkNL0CivU8rcXVLc4aj+1LBXcDr7SZBooC+O75UmVIOa3
XgZN4ybV64aFTj75g2Eg61/3w3mViMWt0rk5WbSzcNv1bV9G/32b4+HYnjWL78cV
HU4YC1b21MPSPaz8tstuTOKnc1fmz8ddl6KYGNTv6b6NGhIEnjXj61YqC1KD/TBB
fwPkHTdK0aoeibIpym58ya2DPNQtTAKWMFnRqLegEmq6clVPL2PQTONBGuk8/QwR
UtL9/R1Eo9Q1Hscx20nDYbclBacVCDfkDCfqz0iRgL5zSKA8UgKUllDV5SEgPO8O
zXQrWJ+yEqkxFenYos/xUWrS858YWxDi4Y81NVdyc2jhiiq6Fu5/qZk4GxBM6nzt
Di/TsCjS8VcEWfFHoQcmzC46+nJFH+9I1ZRiTa5HWF/lOEdsV6QeIymwvznK6oxQ
PS17zQWx1h1cZLDF+91sIwCeufiFG7w41145bXwNcmo2T0OCMQiKy3gUz50vkvNG
qMiNGJajxOjVU/wCz4UQst7duyWLbv/1HZXkSXcBaO+hHNg46tP/6ny8rH6k8Y0q
VAidn+F7oOET09V5HQMRhUzsuAp/m7FTjEkd+x8dqOKXMDEa79HxOiZ3MsZt0tq9
adHEAtImv8HTkWVLgDp8+3XMhr4zLQSAb++rk8VhaK5xKCSXjqAJPkwvhTE/bYcJ
BWLquK8f74Ka7XbGs/R20h4CVg8eG6mt7RGlyC9SlSZa32PXC+ZU3vXZLJ7llCuv
2QOFUSJPIjyMr+pKFnyHYNn2mYOxH8E7eXFqIWz7hwzqj2tva+yExvwwIgGYE0Hc
arwVURsh8RX6sWdRDmEV/wHrPG4OxFrB2xL7vZrvNAPhWFSVv2gx5gKR1H4fYZbJ
voYFL1H0+KBWTrqboieX2Id7jegVjCqOfM+fq2EUveqEn/vXUCLOWaIak5DQX6af
4lo15aPJDzEndD35LnARmZnE2A1cAyuM8bqKeB5iz6gErzgaP76fkShs4Pn5tXLQ
tWJ/0BBRziu7zQoR0OXUfzr+eDkaM/9kLAjM2aiiZyEVLbvCuZTBDXGEwjBGaPA9
96wlT80/yiFxC55HI2CSqeMzXic4jBPxVjiDKj2x7pfVh6VzXgsptWMTswJCMKcQ
DNnfmVGAF/FiIpPT0HB7gWQALBr/jl3zTNpyKbB9W2aAnv2Qdex2R4OFaB9qA0cm
9kTL+kesCmU9C7VKfpeMdRn1OCm/SA0Tds3gUBl6iM/UTf7qpjVJkv3NkF8r67ic
Hz5HAFyeeqBlGEm7k3hZzb9huJuobQ7PhoNsim7IRNeLvkbZGCJcKJtaIq3GYl/f
wxZRhgMw1t4/EWwJHnMY70GSxSnrOXSEiCv/ThkHvk6l9RuBtzJ2OmTV27QkCAvh
3Xi9RZuwfZ7mnZtEbYeYToKopzmqG9ccB1b98p0DwBow80dZFZVhWnoJx+p1Govc
rkhqMn97Del3l4jCEPO9Mg9G5lMEJy3PouKdSmEbnkbrzTTiNBENTCm2P5qpPeP+
Jf7IoMTwdXUx6iNyycGgWwnyN41efLlym1vzLwNO8dej2vnJdsGV3VlhjVwIfjyB
QM3TXgBWhT2zw5EESSqEdAEugqErtfCP8+NqunFAHwREEe0qY2BuqSVgsfUpPwhc
uQBfZV2m23JQAJji2Xhjifm6XFW0P1Md22NVYFugKUnOK3SDNcqdFNZNGjuj4xOG
Wft0r0P2AM0wgxsr++VT6GXuub9to/CrxvNcrOIX4GPlxs50kt5cQLud67f3YVpe
ia7QetFpGnZAJah45Uknq7iNo8fVEvN2BvWlYlV7hLSDs1b5+IFesNrhMdvTjsFl
qAbihrJllgADoTzvzR3fXsvX4VuF07a3hDv1DzmWE4Czt1gP7LWPKdrPQrKpSxbu
rBA1znV0/WnW86Lb3G8YlFsw69JjcDtBJWpBIrjBUL70yG6Z7e0Ln/BWpVqceeqw
FfFGS9TEW5KPpp4sW+ap+3H9rJwepjDa/W2j8JyTEDHu1BqkaTnbJfKHnfmH3aAa
9YJmv66y07it3Vomh22X/BGJIHZifYxt2VMKK+SeKzYjCiWoWbqhNa6/ln0yidgM
DjrQ2Ho+eTmye8FeQbQodP0WWS+oa41CrJb/VAgueguKpKfYesVeHIcAg5n2Daou
UR6VaB3EpxlrmmGqTsMz+mfYgWN5I/pEuC+TrkOmWGQ9Dmg+bwaAGg0avQe+AO8U
CvST2JbPqiQKDQLFjehjh+qjJqZvAe5F0R+FaKQERt0f3iRY7jUYFb7duyVD4Eag
MKtXccvWOS9QyzVzsmluc20CH8bgUyGrMxXI8JS+gJqsytXB6rR1GDazYR486QFj
/RvKaOyDbr0JMVeSfays/L47GjBRmDWaIrnJrDuWjjEmXwfbvgs7PwDUg07kH2o3
1EQ3PlLEyhRnDu5RS7lRFMkKkLAQwhXjTIUTas39B+adI7I/vL2T33tWJaGCFjyC
G/CbOGTXv6wRi3Fy7VV2Fx0HhS2cmCgn2McJb07vxoscyyYL8tKM9YtxxkWmvgHj
iVVvVNIMzXJ3Jw8/uQVdgrUIbTXZLXUPrCcLfF0xTS8Z96NjpFpr2QsryyiRsR/9
I7xr4MV1J+zsyP+oJXNPagyO55uLMGBzoEkfrl0VjaEVrLoHEGz/GEKrY9OoRqKR
KsQDvjWMxWDEdlZZL96DUm0OvoThjyHL5oOD9W5Y8LQvaHByBLyJzm5OSro9027E
trxlOjSNHIT6hT6/Z1Tip3IH1vNZe6P9nBUfan1Ie3kr5XDw59E4GJJDzr1HZ3s5
6PG6RmPnst5vECpku0h+OHR9OAhGzXZw4ZrbtwSjfrCb5WxBKEM1YxKz8OyBCVUB
WTLLoD+QdbVrmQu2qooZnxqZL8mkbEz2L3M2RczuRAq09zXvsWUY4UAV7tQiH0VN
SQtowEnoYwgxa331KwUUw4vBCN+jfyD4vWs4Gxsphw0tdVFXvqMaxxiXJAkq0kHJ
9lPwd5bhryusI14jhEom2V4yibffNiGOa4dIrcDnPjRqBck0ZuijdGHyvmPrGjr2
KUDIDAqi7WpG4XxiOzpRvb4iAos5GuT5oA20Zz1P7w4SD44svM2EqHRBwH8FONrN
Puoo7+4yiIihIG5tAqZWzVuFbimgQ0jMx9YYtZnIe5SFz+LhBzZo7CaqnzdkczHM
R8zfIO5F3Fk/VEKqmpuqTtC2+LINmL3VYKzYuVE7JDvQDcWmyiTFLXMIGtL3cLaJ
sg/loxfjUwHzmWYyjivod8IjlWWw6195EQtQYQsPPuWDFIWy+QiVbmUx+3nJHmLH
z9i6co4mcIyI9QPX8g0gJZpMNxLoj69Qbhvq7ssj/HVx0Gwjae9tE+O4nDsaw/Z5
yWLTH0O0LNo0Jcs0rGsVjQua9OskNX9td0VBpkkuxyHZ65cFlVfdVEh03uYoNSIt
FMCfX8dFoxBYUS0Tvh04CzxJPdwEaJccjbq47Ln+JjSLIGQyoBNEmQH9vh5k/b5a
Ano7nLu600wIKXv9gnJtCCfnmVOWD2KqxAyxx0MEBF8WkA5eNqgx1k2cPPzybI6I
ZNjfBPX0FHaMbGj9V+1aadTJGPX0bBzaH5DKBFfB1x0rx80TDLozlD3SPbSqnL9Q
C335q1qfB+4v/+5WeznM64fjQ7/CKWaXqSlTIrY5cLBZ2h2+Z9sSJ9gXkgrQ0esM
cmFBx1ybLRJUg2EVTRvi1/0QIB4uNQsBVY3HuGTHf1X4+FaaQ4ut9wcEJtolvDxM
5xsIo8W/LHqxCITxQ57Og8nL6urTYK/TUYje4/p8+kZZXsG38XXgWArgr/pc0tgB
e+/7dXBEQdvUDYHlYeGAg+YAzzBxmvWAFYNrwwNLDG60Qo4olh2yrcWb6JSd5iYp
dtXbtcHbQy74SAd/TsVYfxhPxW4RUq2QzsUNgKRuBs1zt43ZC2H4rol8+3IlF8bJ
sDoqYrNqpPnvGzxSOV6Ri0KtodN+2IzaxD0mVjmXuEyOo7pVKj4VBdUbcZcEQ8sW
wxDqU7A9YhAHRa55ZRI/kzSkANfmn838OjMRY20MIlf4AkXDdVN3aVZfe9NFwaSy
N2/jqLxeqLQIQyz8VBPuOOV6TZSXxKepuFomm98xkaaTIJRNUpo94GMHFOCq/Acv
FkpxA2l5xlVVptq7K9xAZRpWybVRluAK2KfPVeSv3a1brJVIiN8jdmahH6Sy5RuW
62ZCSh/fdECpGwWuUDJxBEHjqSvquSZNzR3cEAHYmyUIv/GQhd6WkonV+Sckz5AN
mH4BRII6QE0J4J5WpzRzVehkA45W3dYRADQg2i01w5GptE0mT/acb4wZ0spxhGtc
NR1E5t48cqC8ZoIh5y+rogINcm2NfvnZJFmBm9EhW3sovU9k9Y6ZXvM//jqWoEBe
5rF1uCFyI0+tYo1gEfFivbpOnh4nKRQnzy5KbBKNGvHT+FF0FeTTvcKqqX/mseDp
XTbkwyrQthzejrQOWWKIbiybHeWwbYbj4YJPddoVNfqnQYEymUiAq5TV5MKvjmX5
7n2v0tHzIf9u3GiSaaLHGHGttGywediVbxsx2M71o08L1hAgcEtIIbm27+RS8z4+
BSvTUbF0RV0qUz7urx3x+/2uDTLiTX3W0rNbu3DDUhqxtFO2JfGv1Ut5jmsCEf9q
P+f4H0SPUqgzQXhYIF+xxElmAR4trdMjjOYeAhGa65ZqQGlw33TB7Rqe4klAboIS
V1/8LbxwaFnBUOeG9vKkKR4YvIEknQNyGeDp19O8FCpvIpuSbGco8iHizba7cilO
SxGSUyS/KpmtcZ+/6SZ0Nogy2AOIre4vwy9l0K89XRE/J96JcS78RVtNS+8Oxl+c
E3QTqvHuHzIKmtAvQLfpQmU4YrZEvra9gaYcOZf4Oq47tB5sXgkliA+iBrBrZDH9
iNzORIZmWkWT2iZqllGDZbl8TrifG1qRqrjrs8rryZyb5ribmMZSnWIzhyzjholL
/qq6k4WYMbXkGOKMYdpf1gwm3Jk9SV15H1ahzn4KDCQ24Qm6o7Wl7XFrTAPRqF/O
l0k0eEGJsxTgNk8NHFiXfxRdKrwVblmBQaTgXGdW6TBBqb0C8w+hlRsNwNoXKs81
OcuRGs2EGtH/oqWRPsnHe40Cfe3O3z4sUuaAAFhIn8Q5HnsU8pdnlKy86exCQNR0
dtoav9zAI0iYoTnnL4d2vuccZz+hbC812udBRkcASkzPLcanfVqUnhSzIp3QW19T
S1eVYoFALDIYcXjQGyWabyqgAbHF/AJt+AG+A9aCqJxOC/hfTRZjJ8AopuWIktZu
ausebbtbYJpYMq6QYvsSTwcqyVdda1m4Qv2Gffj6AORbc8Q1Eo+U/8dGgydt5Kur
OondXFQBwxLq9l+dLHHG1Et43XrRDJSLfSSKet20Kza5lEOOasSL0u/KR+DcC5GD
zUoCE7erm5irhLHDHtzNG2x7gnYpHMiNFSDeJPMqqMfhkcyKsAfN2AHS0y55+1RH
maXp+Ypn1jd0x6k/d/lCkGux4k2JXyOKfpamnmU0u/bMQIMwPVX9PiCF753S7Ird
fDQHB7u4deAcBo0vdFcktvLOtTlI8QL6hn1pCKeUV4AAjX31LfHMHNjJo6Uv/58h
xvLB5xr5JIh1oeDPsdi/8e5CaMnVtsmReUuFOm2I7fhvItFx5yH9x13wewpHx9Ov
1f7utbkyQpPCu6b0zPUBVsBbFmP2Z5+zCp5eenC4yvwEeFAsvsmc3c6xlD9M6eGM
Ls5XAYQ9MptaBip6qhULRNqQMtBj/tyPZC4zFMNahCtFtojSAmp05Fb1IVl1VrpZ
Gzp0bgvBC0wCUyKBzwP66GPqUM21Ax7R6Y3qwgDEXymZGXCBqz16LuDtu6+yQrhv
9E5HGCNQRfI2qGRWZermEZtb9hjXvyv/MSyrMYMVpIS9rzgB/fHIvi6BDgFKnRmc
9KaVceZa7Yqnf9Ew5XtRTjYB0DXx77TIujFvMmYdxqqRmOnGqUXulHg43LSwrA0H
gDLxagqI0V+3tG+Nv4LqLKnsR7FU1ZYIJxidMOxt2vSBLdR+Zj1Vc/RwpptBJjgD
CLDJ4T99PA5y9rQOJGA0aBqEnA623OkOlWMgY8iYSD+/qDG6MM7EHq44xCIevO2I
hprUsg8PL5yBlDxfIx6gY+WuIWaWLJr8rTk42ArlhaZ5gP4cRGIls8PsoXLbR70h
/gAvfajcJJffWKYAZ1Nq1dOSofM1nF1xt0sQPzjcGxdQulF3wJhBW+eKBTo/sghJ
Y2U6rr0SoPwgSTeSII4WND4fhyyPRdy6Yq17s5/n+I1LpXOoOA1+pMhHmeZRxMs8
VhQsgXqEgrYExNyRzmxAf27DsDkwroLF6mVeLym92U/VglkYagvvpn1OmsL6IEPy
CgUuUmtDtfWMIXQpV5v7sp7jDShi4qYdizpJKnez9KSWtqLIVlLt6CuuQg0vXEj4
SrylhrshlnyR+8TU7xGLNOKXuXJH1IEJ6faTxXXV4vZuFXGKYKWRigE8SmuVNGYk
NWkCzKxxB2WAwOYdGcdBmQprsjvTuWquubzyuTxueot6y77Oaw4B6zmkrSfsf/BD
MM7Oxlu1QCdM6FTECgsirStws5BybCOE8mH/JzCibaa5v0eSx/mlDETn0fefXSmI
3bsP//qFy3yLlcTamNNIb0qQoca184shrkq2a/aCbr7tkrbP0Vi4XaJladOcEyCY
cjKPRXtVIQj9+7tzqDP69qOIqF4lwhDvM6RygH54LFhEMtGonE8998ee4ss8J7e5
w1Qp7r0tqcMaQo0rUdJj+yc9T0i5jX2pPnptqgKZ7H3O0jhrKmmatbtaV2ACSAx2
eIsB9gquHDJ5XtJh/ZOGpBFuNswaJ6Y60bzV85/ojsLGE+1WJNBDa5yG5zREYdxf
zfHYnJ8ufbj+JqQ+b1jItKGWCabCiZOUmbcj8K6RsJKwT7dd9oxPtw5+UYCjw169
2xJ3307RXWTNhlkU8gfduf8EzDBueoGOwwIGZWPsRZmgG+ViHVi1cf+ZRd3aTlWH
MMGP5O/Cjrq3Jfo6i3gCHVl3JjN4na/HwuyzcbXSgfne+B6q8MSa9kFqYJEkqN9v
pgj13wiQgnEbJ/MiBzcDGWQ5DKZu2/uckHBUgHEoOFtyofQkiZfroVzUJ0iQvdQf
gOSEI3T2uCCAP8QSl+lyeX+EmeKzqPdyPorhHSrPRzBbEMLJCjXlm1keV2Qf+hMi
c6V/jbZvMpJxS7LbGgrpcLTo5HpBiBR5McWAoXqYjkBmLg7GyROcgv4O+NWrfk7Z
s/zBvvicmPHTcVkdiqh6SdGStjFezw5BWC9nCnQoeqcXqxT4vXmMKo4y07j3sS8Y
oDSmQtv1s0+QlRQj1bhYEMw7fQ7+/aWQDJYKYEpRZazlrxc73UgownPCd68IJUsV
CFh12iLPfF19Mat/ScI57jNb1XPANKrAxwA3Q/FkI1XE7OFrjIQlx50wx+cMQ87i
mIWrMRZ8biqOfJMsMduMQ/lA4QU1nsot0gWVpdOZVRbTRZL/wTI3lRlp5z+KGzjl
Zmu12T0Bn+hUyEyB4LsuUiGpkJ5tVJ6iesPYHtA4VVKKFw7nmfDL45w8s80aUNkK
v6/evpHRpzzIebFB6TBv25KlRap5FdQq7MAT3ju2U4b3upjgG5FSpCFjEvIigHqN
ynIR2DOTqFmyktg8iaoV+oHOZahwTFv1D4EkpjoWodacwN/G9erpGnbGDrR5vtxM
aIe0SxgIsgsPYkuKuOwjRdhMIuJCB5j9tI+oozHZ16SLKvAoOg7F51kjAJ3cm1tt
xJ0ldh51MqlL57s7sEL9XrbFJdOOmRhM2aR1yhSZSiwI2NKZVxjLqtOMypq1AG50
n/WAkq15g/i7r+beq0qa9v2Tpes95rKL/UE8DHLlhBO5Ok+ZqPszZZgztesGmpn2
o1cu8Zmzkgrc18/vvdmzePKZRfawze6zE966MXQOZkv777fnko5fF7OdEaeTOff3
FrQHeMJsDrYixcH2gE4hnznDJ629ZHKrzR8DdRAgy9MhWB7SUf8bRNSCf7RT5wCd
VwRSgxZ5zBoo8CBEbV8CRBhFpNsTGz3KvdxZnximp/cMI4+Ll4MFjkUM05HD/Btd
YaxbJIDpuz1ReRS64mAYMj4Oy4i/RFAHKE08CLFWY6a6Noi8szbA4rllx3kyPodG
6OLDsdV5AS3iIjHRyg2s7/uBqkz1qpag+II9Di3veuWV6ZB7VI/EsZ6x3fP6ctn9
5l5aAzCtx4u1nBWig+s8qqXwTuBq3HYymiVZzMlzYkx/c8AotTQwHSk8rlXTCduI
rcEFH3ndQjac6op1G0vOCjDk3GzNv6WoDMxmFtJJ/ZF5rkcX6eMutbO8Y4vD/WaA
VlM8EkPVYeUmSEQMqyNbB17ipb+SijdS7/nrk5AvE948vPINpq4uxvqjz/UCsjEw
VTKb09GsnSZNMu/j+3M3UR1v7T4FtT9AXfIr+qVe0EItElBgzGOOVbqmOAwU9rTU
x2aRAErau4eO8Lnnn6jwT5HJvMH/3wFWDsKX9SFxfyt7Eqgp3yHNzmTZ0jlRhtRC
0txT5a+yb8w1jm+21bQi2NbxqxH63XK2QUzo4jKN5WZutEr/j60ca1YW+G0f15Xn
LlDcKBN9z9h8XLVbwT6OKM5EuF9Qh7WEnPgELRttRUumOhvEJ+z9OdlXIJvFM5na
7xkTBR/YcIungEtN1rL6McU27nKjqdCq4iQrgVL7BlCk071v1sVROp26nnpTrn/s
VEp+TeEMbs6rdWMm5qLCSciSpVS5PIMNP9LMFJXFvCwUWDyC86dOaK6jNt21UDA1
shvRbjwWCNJz3JA1MZyJLv2qdYv8kDcufRLij5fjk10zbMJpRHcKLQ4s9JR/1xHo
Y3u1iyT6mBU/17Gv6CmemnbHfs8TdwKoNFKtIqHyIszK8PFMp+2pIbRcZeQusfuB
WN2x+dScm7lNxA4f3Lp3Ztq/JYrrQqaIRjcLkfh7WJTqAQwKbAFnBa5A6vD49lKS
PzRGoDp5FKvtn2+fegLj4KDfIMC0tA+9+S25c8ZQb4bdrFxiczT9dVK7CH+LwiF5
d9N6iX6IphBGiPyMJC2UlJFvJrBf2m9x4XeQBwrFakXHXeEhRHEWFr0srFzmTRGi
iblrAt/4fEc2u7s9+jcqb2iiYtFYE+b9ZHl4EZL51khB1HqBw7QO0Xz/kb/czxfM
/spGXUu3KmhhN1o1YVAZpS31Tuj7Zjx17wVF/mgxueVRYTcADnGfHavMJkIeC3/B
sQ/WMJjQ3W3CPWEqH5HyBb2X41IFWHEMCzTHo3w+bir7CH1+nuyZoyGOBK2LFTBr
2y94flhSU3icZeEvVK9ASihvLor2500qmaw9NVhFc2Af6WIjgA/WfUyGihrwxpcw
snWwgD7GB7jchKvgrrkmNOxnUu4HqQd+n7qEc3laKHdm6HtW8+ObtNV2eWdXlikz
tLGwgDxeVufj9JD0/SShMvQNoQ9cvH5WnaWIVf3Kdy6udoOnAtf8a7xcDMIjd6F0
0ioioT3wmueF/dkyCEhanpRJoQZwEGvPqqFPkZUBukK0kNbr7M3UBSisR/K6iObG
E11ml3anZ12yw451Z0v0bWzpaKwiZZMidy139ZxZ0F6F9CE50Cm/Dx1eCbGc9uc7
uZ7DU7PRkeSG872LRbIj7RkNzUgtaQuhV/ujsRjObuTeuVr67JtxluadOIRRj5ze
ET9/2t5QynoVfxJ6CFbvjz3ZY0CS5WrvmiiW9We1T0ROF4hkQIQxqiZllsPZdv0s
aSgbsk7zG3e44+25X0Oga6sJJZkI08ovnLAl6oTlQmQlezv+6E59N24Z8fYzTHsf
EF0DkSh5H9c1ArkG/irRynQoeQJUidmfMfbClntSP5bX9g31U9vA9E11Zz/Cf2lY
Qyhk2yhGunxSblAFUCHYxiNUDcmOFDSNNeZp0q2hyeAs3AX0cpDL9f9pzfXf76fK
gAcJ30WOhNLskXAtZZG6wiCSao9FpJ0aZvBaSC5VOIIOiwEAkh6kLu8zbeHb7LAT
uNq1+26ypqdWSeNRvja6ZtabZyyWgTrsNYpCrpnLkytw8kDZRlokwyhfPeo0PyRs
hwt67f0iEi0PnaZfNDRyaII9bVMHjxkGR3w5WCrk8rLqlqkGKYXLX0PW7Vd3heqS
7/tlRC4UlIEWkGn/k7lqvDxGPFCf09SNhGq6DbxhTlorebvwi46Coyc6tSlyGcIU
T//fJ41J8MMhPNRvf4xL9TDw5rOF6Oe/RsPIdMrBPtFbD39V/wRhoi02xiqjz+19
3el4vLyD7cz9lyFrHCI+eg8sEdlxRL/RWAKYtGW9kAT7vcy9GdP2RVFjbn3Km+kE
TAZf9qogiAJuG8XiaDCfhqYaU68yTJVGUZGPDvDYoTfGGA+bDU6cpeXyugt9c3mK
URCAH9SFvippWGYzwf3YEMp4FhBDmQI+nKXi/6C6u4T3vWXL/VjcDiYNd5jn86EX
OMbhqGrsTZm6t3EVHB0/B2+72/tyJ9ePQn3nhgFu7FMb0244caIw8eLpWLYsr4Vr
M2bZviz6fLIr/RO95qeJQ0KTKn++dY7hQe2lAFSLcQmwaqi3+EDA6gQq7IzscgeS
sB0jm9d1IAEhTv9vHnY2VEpJzqUOXfUmDFfdz/gdxSfk1M+YyHakzPlDUUJTL8NI
J9XxJoqecmMbqbW3+/tHxeokTG8Yfm88sT35GnPXo/Qdj25EhRKT9yG47ZFATyRw
8OuEf7HK+Mr8iZU+jazeGyM0O3tbifWGLfq/vYfjWMc2ByWp+OmnVkXzScLdwB4u
rA+lpAUxdhkXw9IFrCZpQcagfip81x+3U5pJ2PLN1Q9sW0NcxwvwEwHcV9ukD6dg
0hR+73qc6c4x9CPDy7EaKggx3YmdnjQX9jfUwMy37XOF1q2ZaGBIOHX0EEnk6Dlx
IFyqG67VUmL+AH4J0n6DP7GnRaSGCfQZUrrvNQBQ8TdSPTGqKMLmef4itNl5Scxo
R+/VyN7u7Mn2GEVTPU3owihUOZzgmK3HsTxJIHGc5GdySmr7uyexXy34rTlx93wG
B2tUVpAGstfNVDJ6PJCTzMrN17s9e0rbXApy48nA0iDBIXTNhqGocJ1+JZNRVM86
eApW9DCBFeLAkdZKX2hQjTC3mkSkRuP/1M0wQOXDVTUVA0tpTfZ0TDpbPSKd4kZH
oUVoXwAcYG2Bzq0mWjYQ3sucgnUksTKlC5ISVzMGC5vhYd5iOTjc3UxCj/7PrC87
vFbuel7qAnxk8CzTDgLK9TLHd9DgIcaS+5inaPWI7BH58MSfjBjbOhNeJDt+OWwT
HRb8HWxt0hKx7URt1yB34IWhjAdVfcNNItGqynPX7WykVnVXTrsBje9Z1HSom4Qb
NtPEapdMHkVLc+VuYuP0gw2axgO+bXsShrDN3OOvbUJZhF1LyH1UeiqFY79mx/33
m2pPQwEoKSO6jMWm2/SazPTY1htY7hjBhoCtB/X8dzTzyKfuHVI+UFFTmqQoij/V
r05qMZAHZWc32x9xhRQob2BBuDsyHS+IftdoeZFIN2U+5jdjhiZ4vc1km37MlTOU
0Jw2gYCtKno1yt/U6N+k5QHlfn37LmbCQ5y74QMsqQuPutgJijMD7fQ3yuqKarvx
TwvLnaQtKbx2XZgq0Ds8Zei1Cg+SwneoNtDjm6HFpsoGVF4Y7tLxAMcRmd4tOPmr
w+0V674RC3s1s1FP1AxFytgqjLCbnTv6V6nwjU6eBTzu9f5PRC2Hre1fXhUuLRhf
bJeTtcXUhG1lCTynpZhooJMrQwpVWiW3WcQYhYRj/a2F1bRaVOZuOCJ5+QX96QFt
aA11D6gXqlcfsuHb8drxjBUR4m0cSybSGVBQTR6DKliua+nwd2j/+JwN+h8usJTf
lUIPWMByyQajAVf6JWecmQISwK+wTS5SHQQP67XlpobZ99G2Itf+8vBjYQ1u5cne
cK4E1NIip6XyWvcqJUGcuhxcoZrPuGSGNZZ3YnaB3XDD5ZkDOELBnia+cyftphTr
MM0LFIoZO4aiodvhCc9A0gF1tkbAh0UFOu4cR8ULh5trCKDqyWUHOCsLepo45GbM
GhnI+8IbMOjW4aQd1t76u/nApe1SfydYUvtJ/+AQum5oGt7/83GoEfAglGpriltN
6rbq7WDns9o0EbVNMOsZUoNZw0h2XXAeULNLgBZXzPjIzrh0yoIvGhfkiQEI3SBr
oGmdw0SYi70peLLE+gM2iRf92dPvbncp+/fyOPZnIbHNSUIylNWtl7uo6ak2gN3+
xqefeVl7oAI++Y5Ny/8jVj95aaXxuJ8v7RMm9zCJtBLMfmkt0F2gbs/qB7UeFdzj
rxHhmgcfdP/ZNbMSUDV/UCdzWNgtHHNck7WpCs5PqkOSzqi4tiOE8aoZ2rRdXanJ
LmYHjvYtEYwqNfr3p82jwWqAqL7BlHU5ZAx6YOd//YWmEK2aTjDdBw2EP7F8SSpI
B+VglWm2+jOO0JsQLkaFkT0XqHhWFF496yItuRXjnrf1f5zb83wbFMHWUG9cazNB
2mmsx939iTNWumr9rHE+EorSiomdq2+RNAlIYineuvLfeB622oDbF2ZIbRCmH/Rg
VnXTVxE1PTrVWiJjom5Fro4bOfYF3Nu4kuddAJ0YuT6S1KODK8BR1Vpn1vyEg7n8
m5qo0UebxjrS7RsBtndulXGn0YopFDGQwZj/kcIZPuGM/G4KNqreuGvv7nLDdjrh
hv+Lx0i6S6e4759EVcnNehOgcRrEpJDP+pnx6RtKaxAXuo3FE7RqJgDwuZeYSpoi
OveB+m3yGFRCnn4s1LP7E4HNHYoEh6AQJGE1KjW8WnXu2jJ+6XS4jJkYOULBsfIB
g3gAeL9eKWmUirgQ9qgei/Q8ut/k/ls1lbdUWjzlXp1nccvrYzBmIK4o5dWs9pph
6kNORo6tOeWdgtWwLndbrpcVt6/UsSvtCgIQAXtlWfes+jFIwX3hewIaDt6O95nb
X/MBkqt533m+MeIgljPQsTFvEhYT0LgnUkjVqByk72o4oK7JpGW1DknK7chaAwG6
S98bIlcuuBiIQK+EYtcv/FeTzGnNxG4jDH7VMRQucRvknhtQs7O+UIVjFZCW3u1P
HMY07aDACUyT7xTf7ifkqWlwCNXIW4i9dhhC6NFhf8M9vqE2jHA5kzJa30zfE2Vv
2FfN/AwzAZpxaLpH3dfur1OkCy0i5LmgpSs4U8YmR0alhnAG+D0ObGggALRsIqvm
hzJdCaX7WHD1teRXu9BcSp+GsafMUjafovRxOlzv+AmW2Hy2dtiyztVIXGIW39Fz
EQRtRgd0oKjGZOYIqaVmyUu9HVp7ETZxq0jEG8zHE2ELZVmece/ABRtz2sgmcSoA
6OPlKI4G/AwiFziQbFC7CWN4Ibje5XM6eqngv7hSGspHK1TfcBiTLfQWmNAzuG9c
HpT/jskqHBq07HLDeZnCTwDIpWIQJDADId9bJ1W4BX5yvtplvSLGDnCxXJPL4WLq
NXHdD2zgRg0R77ZEU+tCFPiXjBqqbAOLBhSnVaeRaAGtEIrYLezXjmJY1ySENRY8
H72KCy8T86IeKMwrw2TMqlBmzs6AGkq5PliVb6He7DKW0SolkvrrerSPA5NkNA7i
8ZNiZOQxuKWg6g6OQnKeiaqxbq1aZDDzrWVksOTeBJfK9T+f12s/dJGsX4F+pblB
NnEiuU37PcC8hyzIo/cKDYJbl+425EHISRafalN1S/LdLCzP5nP60Vjxt4rsBZXg
GFFBsl1kG1Z2gTOJPtHP+2icGY7yjo1seiAv7I6dq5wCyWBeRlyR/cQQ0+wBcIH0
l6Vas7ScmyJ6z2ytOQJVXOM+PXZXHh+jKzRQBXXznJGzpjF+cVz/RCK9cBfnPo3e
DfULHb3JUfrmkUfkKsuoaHKonzu2xfPos+smj+FyN67iU9gYVf8f1W988k4RQmTH
XcXaV3cSpL558VywQDtNpB07y2hYYDWOHGjM1d/TsjcQGffXtPfwrvAYiiNQDZEf
QS5BaOPY3ERlMOIGiB/KiPD/85ZsP4qvTwpJz+PO370mSGn5WCnRsnZaIifY1azK
HnfwPESrT0Ht1N0S6vmdmTIxk7PT9ElUMeST0rdSnsNqJoEPx36KCVpUuMIVvMKU
++xtW5+AwtkvK9QQhg5JWICp1yUd5CQ6MM6DMatfSfI/4FuNKsAC+uH5JumCUTWH
nIM/jQZvwUeccyEsPRqv1ExfKEeztU0z/2thsnEuOToEyU2nKqBOVqlOy2M1ghuO
XZ++JFVBDLEdnn6TqOA91dcEJH+irBoYQ8nJNUrGRWyMamOCjcg836Hyv6tCjSmR
c+ARZKaSTqzi8ZopiM8PDILRTEp197xr6H/Z0UoMwa5KAuYWELxen3kraQwTXfJd
BIFiJixzOGYu5N4U59PdsFfJrDDz9l+HmXxTcUCDHr0mTU/tXtskqQ4t312sCSCE
mY4Ojt62fwFnX+tM+Yiwv4YNSOHHz0bSo7Pc86TwLu8pN1HZVh9a4uNAFH/dI1yU
RM3N4JqLojsd342gxIFdKA6GL+dTpk/PA1Wp/me3vAsZJme1MEmXl3YyYxnp4+v1
tOsY8HE9Uhi4tt1yBBNLQ8uyb8llAgl4xewSqWp2jIIKRYmEpmBLEHC4dE6hoy5I
L8EMm99cI9pz9e7VAAeCP1Y94Jgnh4BMmzIGXLlGrvIPUfR+Rrq2ewyQzHTxyo3S
MIfoUPZdQiRRigrINU4E1bchdDsOLnKG93y6wVJAl2u+UKiOQxl2WbFhZ0adRd0Y
nNbpGcSRHpR0sdjYRMpinpxD9DiZdJ9ECE59OTcD3MZuib1TLR1FcEFxLyPDwr4j
1/Cz0GMjXiYGPNl1WOK1yc/srqpxFDbldIg68wXaf2VRC17gwz3klJ7WEH/t9DH/
vX3S4VfvWuEGRdx/OA/yev2L9/tZrrSrBur6VuGYhaLzeJG2Q90n6aBwWh17wREX
E5Qx1WrWAQqubDa9CHcvhjX8zNwkROKmBGlCafl54KLfxnePIjlxM/X2ufT1McdX
jVcotbJdajUNdO3DYaScmbppw88lMF6dAE94LqWLSwkhvqLAZZExSaSaMoajvOdo
LZ8t/gW6BDoLUC1DmfKXipNHvObpYfk4CHbWLshRozRXvaxSrLyLF97tZYtSK5JC
DrKjB7mkr7eSzS9+rdSzuUl4f+GA9eV0wnCEuKBQA/Nis8xAKwzVxMeIKL2Rlpe3
y01zWJ8aGNPnXkZghnrCjh5Z+Ysc7CBeQUqiCX7UiN+HNOf+dB3xT5zSOJihCpQ3
H9QxlToZpHjyBc798VIrKlLVviY5HZOwEHDRsXkDdYm6YbM66vOx8t1EXMloCo6j
oLDKFHZhMiGj94xOf1PsjGILZjHyEOktEF2BE2FOkHMG+g8OA77OERsEdCt1Q8zc
NzWZC5sGwuG59MxULG+/sjLQfw8+ot0gOsKpQE5W3joqfVjf403T2EOKJUZHTHUo
kpBZtb9A4dekcyLV7i8uBqRiQd7hi6UkEsPDH1XOecGJHrqvRP24VxUIDo9z6jS/
Zke7u3MbvVA8+KI9d2aHGxal7q0itXtUu6YXS48wqyP5FL85sLa8NrMFO275OcBB
VecoYV3Grz/4KJBmo9QfDuZsYZGC4tOzZyoXfBqkbvy1UTn04mq/qpQS+n1xJFP5
F4BVg2RujBdnOPkvNHFfdQmjfHVOHcvnA4Z3Y+kcZJ+1EfLx5NeVE9oJ2MtMByLc
PNMywUZWQ65ELyLLAAYtxmmKTBAG6Y3CrzuY5bj65gv+07wRnRYOuGAkQCBH/Z31
OBZKYvHa7h5cFFX8yZ5k7kiURvVLpNSbDfNMQuBLcvYRXaf9tnKayaQDY2JuBBke
i8alkyTIjVLMaCERYCuOsVIZCKvrSPqm7i8VNW1ZLpPfICtxewzIbndU0fe90Wk6
b/v9Zile1vSTCBlxpnGY+6+hpTH1QXR4zp6/Qyv4MO5y0kUf44fNB/+PJyKh6jdu
ytRvTzFeiVUZDg5D/2VfYJJCAwiit3/4+Ozo8LhB1LmCVjiU3LWZbFLlsw3tdeyP
CehPcUSKtiMzKsx+gGY3VbUEObeTk407DL06UATjTCDfrmTLQuzc/TVU1IACf2AA
wVme60SmfnLKpy/B3bn1YgvmlmPG0clJfuDpI/dUwwYmX/GnzDJzuFJ8ry49xR/j
nGIGeYZsiz1ByYO4TbeztYoA1E/WucLzzxM0xiJfndcNzgbYxTEh+FkHllPkclW0
3jzb0qNf8DXbiMmkn1kTBgc6ekHCvvquNtowhHZCWShZlTOJ7Ul7rAc5ce2RuA7c
3tb04TzVNSmISEyjD2fIP8dMqoiGaiDbSuWE8lghllTTWyn8c/EEkq39TmKJ/RSc
ThQLpfBMWazYICtCk+w5GXHaKv29AbwBmbuWfsewdjXXPclDm5NZRvrj2aPdoRp2
bV6AVPzUD3nKl3KSL9RU3RiwrD7Tb0e5ypu1/gWkSj9G1kUfuq4PXfEAwrR4SgnE
gjy2XwJtZRAhmq5Yw1jUCb0swERQqjHLJE0PC8npKdKy010F68BZrTOYbtqQQ/OF
CD7xDTO+SZ7r59yhicE+mzu3xafEbAaFM3IotdupVYmpX61RHL0bHSDJXyxyZD5D
pUkKdyZ5QRrp+drZjKictJzk49vOt0boT+i+NfKIDDCdMiafpOvVLIDF8FKtBdMj
nf933vQpE+GGxXPAzKl5S+F/ef+FxqI1wTlC5xE4NZOtZK3qErt027YnEgZ+8RAj
Q3efZ8KGWuVbSxP/MfWkI8D59PCYt9g36CVLI5JUxfpm8J1BlfYEsDfaVKV4AoiQ
GiJ/o9f9U6m7ZYvr22yRHGWKEIDuflQxJZ2vU1+iz/eEVX3NsOrveduFEYWfZt/B
xy4BVpsWvVYIRc/XLzywSm7Bh3j7HxsOkRND8PhyfBfcdewFnV2+PRQsG1dS3Dio
CJfIh1lUkRJmjtz5xr4yKdDUDR8+a7r3qz33/g9Vw0aHawQUeG1Jshtv0V68XiM1
44j/DHMnjz/6uQyWKiwbJx46aMazjoJ9vrBJexZwubEoqDfD/Oek/Ey5vcIYH57p
v5CaVhrPnnBYvuz/fjRGasM8ZExwZ9YNmMPfQI6cOLWQTC1/9reSfgkPup/FU1t8
/YDEBBuj2dCiBJFWCvLisYdUSFf4W0MVLs/xS9s513nHysSiZVEePUMDug/Jvv9o
w3BbebuhyNn3hTwMkPGb1JgelkcmeJWX4Exhchn2XJbSOGCmu+t1GzAr0c2HmPdZ
8qrOp+/tDwkD61gTKcGdjlliQC9tywZiGhTHRxmxE5Sav9SdkJJla0Z7CRuIKZkZ
HFguLtcyubeYZir/+Dgf+RxGsUuQPCw71cMKkgqZRAPVj1Ql1C3IAea0rfDF4/oY
hoSd3J8yPRvcy+a4Ffd2v21JLdCRx/e2dVjQbtWYhO5/6gJS0fvQnPx9Bwq6kwdw
eYELBbFKYramgA8e9dPElug3Vm0HxJWcUbvvNf2+C0LPnn0VPFhtJLAk1R01hszk
0PKiuQ1yCxZHUzkoARTfBZ03yp3FVEDpksNTlZhnSxqCzCSnpE8w40Hk0PTNp6+n
RI/aJ+RkjgTT43U+tzMx607KYa7PUf9Q6p6MapsxJyjZrbNWx1j3gaQHEomsf/g6
E5gmOYWbbhUuXH9/FGxuYz3eg5yKMzPKNTVJV53/DGh61RU1N4fasdATVDCDDgL/
4+Ozlf3351dqs2oGBL4rbuouG+gp/7AA/Db6HrRV4cYWGcjjbWUeuzol7rMNJL+q
2RyiDd/nco9a4d9jxB6nD6gwqebpigWa6NMFESrQKmJuNFkG2h0FM5vx+5DCr1Pr
nGiSZdxGh7ZpsQ1SUf7tPzJ1OiUyVfCw3gN6GdvVzL5FoxNR0xuvT5sDq8VCCGyI
gbGq5exWcTqrwSejm65Hlzhp3R/EWMFzjxinE7RdpFY8ql+zSPeePbRBxhAKZTMR
FpZ81WwSSGtYAB64EY8OqQRra6htDNPlWF3BLea43cqQGUsriiNhrwzIGyY/bxv7
K4xR5dxOspdD85ba7lwa2q/P9BPP9bxx1JMEdQc9l97+C/8BXEOUDlST2QhvlrjZ
UY1Gjb4sPu828wW1/1OvDOEsQpAsckdOI+XdKs3+OnUgL7V9cQViWybp3JTRHmDQ
lpLYKDLHqIzrvmNisIyR0tjidF1z4o4Xxg1j9JwFP3ufd0S0b21l5ZOZW/wlBOb+
v2LXw3NbtAcMfv8W0oIvMIFWGeQp0hhgnLZZ161hZ297V17l4LeuUwQfQppjT3R3
8KT+gGb6lAEC9TekwCUonufTcL+XdFtkIqfKhxmAnfK8Z+wgA4zhjuAfGJrCZjal
5qavF/uwfdl5jLYgOIsrYLRi2EZcr9FdHLbV2vy0KF5xTg05IecZtYbQaYQ00BY4
UCONIA5dAANtKo9gqQS/wodDvCcATnhACdBIEEIzmtY2hoDmDF1zJcjRa0wwB1m+
SISoQusMqJEhm5QlTaZXeZr4YWRH4Bb+v+B1v5IBXRYOTk3cbEJUF6H7hxntSSNW
e0IyazRkH5qSR2SAL8qmcpCwSXhe96II3hljq22TrZs0dQmorlMCD8yg0yTSyBg9
mjYT/XqkeEtJr6gR6lVatzzFzo50OKcIUMAJMILwyzD8sFEBcXchlQRfhXRktV5N
d2nNUTq9a2exqPtZdQ8FWdQiaynYDPFcMBPhHVlUc1aox871Jusul7yRmkRlrMGU
hb/wjK7ms0yYDjq1RRHXud/p89bLjG1Thd560ujEp+nTMtNNCLOSVV93BnHaRDrr
OTk2PcFETjMa/QZ6TWe9ukte+0iDh2GpYFJU2pfU0sQpnLJpwuqlS5nBgOOvtc1O
J+mQ3RZ7LhQEkp6VRTYC19JhCYj94khNO967bcJqmQcR5Ij+kvkPY/eH5hgHnvci
0/EwYYGt3eCgmrbIL9+maxIN7KadqGupdLfK+6hyeRiExv3Q9zQsJ40nyC5tKFic
wMf9giS+qBHEQrLBn4ylz1UK2cyosSeRV9DYpRlv0QLVDW/DhD57/1tWztHIIGWg
PwcsRk++QRbtKbx56H+EU43U3Ml/uLReySPN+8FOWA1KvOv2I+ycLUUH/53alUC/
xc3Mc4EZHl4X37+X5aZQKGUZBUeVnzDTfIVQ9ZjtV/mF2qB+At3vjRtmeou74Fp+
ChCwETpEfd7PAPxxEwbpKy+KpCEZAYUha3Fvw/TPGLKH44FZKyDdloNjpQrW8g8i
32qBFrjGgEjQg6PAXY7hd+xzq2yOt/f9t8sFgoVSfHKBRl4IG/9qfhqGi8tRItKP
hp7TTMueG/Vpgnp0qXX01rJYFP/Xf26KLOgA6+EJyL3fSW8dsIe6jU4fhJHH6Oth
Kn4jL8WrsB7DG28IHB+5dKx8AwZ/PkffC7tpLQyzcrdJgkcUKLfdZA4+B4N1M2hl
CPaa78p8FcUwESvsX+lxR81hKPaCvDoJtjiZNCpnXGn+7VU9blKnv2ZV7qB7QpeK
v7ThqsuQbaaWcYcmn2JdErEQ3kOHnp8C1j8RoX9j+gM4+CJyJXbAC7tT73tbgeJQ
Mmu4zNo0+Ij2bVE2wqVYYtMUCtWaelnoLeHcJeCoRlbQn9tT6qMfGUERCDXXZmi4
sMboTwq+mwgVndq5R9e2XqRr74NHFGA5qm2Y5gN8vjpsh1kYn/x+wV0R1r/pRQ4f
t4jfzFYfw0VaWpf6X7R3vcyHBnUxDlTBLAV/v31XAqrFjJG6TZ8BCz05rkfTOt2P
HjrMk2ECEbfAqVMvbLxziyAKnZCffDlWs9DZniX6KujDjmb43s0bU9jp+cDiTHrz
1fQjA4SXHmQrjMehW4zVHKA77GIOkULbiPdUclzQlvKQ/6f+q6DvTVwWZCIdPv1q
iT7Vu43LlwzJFKpfnPaGr/F9xpj4oZnAwMpsfKAoQSO2wyIoVCkYRF0Dlic0YUHQ
yyJlunO7xiLzfSH2au40/kjYa3A5jEnopRQ8sPHzuo1NVBgqDp3kCTu0CfTpT58t
uO2Zw8RKVsepZ9PtmCyodalltaH4+tlxg/HJs6uP1shivMlzvDR1QI/MXVqEkQn3
il4GCLDzh7vfK9qSrl97TUO0bw8dIUV0DE8GFuXAU893hm6b8ddo3rJDF7WsMuVZ
FTm5HVPAloezZG4R958bh4jXNBgmhpH/hZS2vOnuFuGCbchb1CQr6+QfIUUI+Fq4
MBYj3nQ0N3VpleBkKvAJ25qnyeSlwwAiKDZOQHFX5XfT+NsdQA+mVD2ZupNe7uF1
saW1vsBhy7GKHK4BWzt/y7qQsSC9283H0TTaB0+bxzEo95cDf31ZuRZDgLUbVhLi
L0g5yMejcXfRnMB16iabABE6e3e+gARG/YJTYlYOoSSRc/WDYKcE6VtrDjaHYi3y
a7TQ1TiX9ArPly7tG0Tn6beyuDeMtqQ+mML3zAIzvqbOdCM0GFTWGhcGqz+OLohx
J1amwzJvd54+3/0kYlnV9TiIv9kz4xr4J9DPYYgw6PVWFwj7wdjM9Gen1ZsxK+Nx
LrZxYiBQC30A2ATjO0AaotCw3m2S1fgpKzlU1cgW56J0agTPktFVFH7DJ86hBT7d
IKERuQ343B1sl1IBO2GQPpDbU9l+aQUEQvE2hGMPIwG+4WwZRaT7FJpTRz1bu+I9
EVPov20SRiAIrsU7RpZFJQbkyk1kR9RS4EOG0n5qtSRjfY3a1Ge8Er3xiYFhitpl
n8NFpqIQ1Jxdh8bhA1OaldjgNNk3B8mOnvM83vwXglbR7z7q2TrwbYDG2O72pWTR
CiiSmUX1vb2lIqYTuKyz6rll6lewzWPvnRcUaFGQvlkt6upaxw3Qv2yNx2ed0M5E
IPSQ6b8r9vFeS76LNh2ZWXddSk1l+4zo/SkiEvi1W6GjSj/yqpKKt0RtLepDzG4x
AS6sBU5OmiVBRrS2pkatCuKKcyuYTcHT0ItXSJkiuRsR3oD2TtGp2ev62leLReFr
b0QofI/SLJ4qUj1HoZHe0CxFYcpxMQ/+V0zvGG97mOGhB9EKEfHQtHYitsVwDZxn
tV8SD+xyZ/ajI92+faIBcz4tDGcN9lMTGM/mlDG62Fr4EfP4nAvapiQP/Y62qIGI
ytoFKpAb+jhYTuIM0+WKb1678yJHWHd1tW/jzq0SZD1eEiapmxv61B2r28M1nRq6
XzZKSAzvXiQR2E7BMG6nzRzUUls1gqjAuh1+wlYDkDiqr74EiP4CFWlJORKDczoL
pTye376gxYMT6NBcN2Ps3dQcAB7QuhTJ8gbX2fgPOWAstif2FSEL+Oq4UTUmO+oh
mWjFXqE3PxvwQ1lEy+w1a3Jgp1LZsL8F/wP3Q8Bj6BpaNxepvio+IPW4LFCMEfSK
z9auV0e8o+uwj0SzLH0fOFZ7rOQYgE1UBxFA+JhV3xc67BK0gZCmlZgm+lWcPbjW
6Lhf65WaXAzqRyu2BF3ur11dK+oOPhVY6rsbLUGUZOHZjtcPBzJQY33S7Fkuj3Va
yTpTHvjRTLhbgJBJkKvWVEBghtnQnNeEjy0nTxPU7fTxdkdLrfFWMcpXk+sYD2L8
qjYNuGSw6F5HJOhk7zDCCZS8Mgq50/P6haeyzq1YQNV7Eof3+pFwadKdwqymyIw0
8AmDBypKhdqYsAWnwpmTnjy+u9VV0kPuW6J08Ws00Xptg8olYT+xpVt+EU5ygCC9
Xos8eLIiLZP1C+9hIbrxcv8SdAokolzb3I0LU1iEw5o+7sBI5jO00MtKonsvw00H
vuu9HJWEHWynRQWPQ+kUixlope65NrYKHgbl/8h0Y8gVeTeHtsFPMxPloLDUm0nd
tn05pX1891XYxHTsJQ27q0ZH8RCiWgQUaCCe9WeTj/YMWERwHUOKeMA3FyYzB9b4
GocFcGsNOHD0lnHyzH5YJm2YLRigvp4k9pe2B1ODfz4hyQ2v4djvwO8uGzGjoyN7
5qMUmPjNX4+Q68tQdcXHiGzweRJVn5SBZXQyVnzCT13hf6nk0eY5aJLXx2RIaso+
1Rouoc1n3pXf1U7JcGdxtwy9ieBVjzpCoiWOBzox8J2W3BqWzzcgZM40iwmkdS79
dcq8KL7E+BLpnX53TETBCFIKyX4XrTaA57kFuifTEzqrV18hU+UxIps9KqGX/GOZ
RVvVPC0Bam9rMzQjC1huRtYFOzlev9Cyesj58ld9T7zw8fiiKJMNHYpqYbi6rWPn
vKseP7kEB5Efo9LldI5p0QpbI8+FH6S95DnBqfPEKn9m/APLvi/nPRmHDcM73b6q
Uag1n++btLxyZujrVz0ph6NOHpyLw09UBpkUadumeNmth0LARDEDHODaMOoK1bz2
gc4v1dJcI8VaAraEYSrgQ2ba65UTIRbKkRu4tayRF9Ayn/O1yOijso4/hjZPakWp
GdIXD8oiuCI2M29pgJj8BkHPHbumlXwBu1QpJuHkrB6wbCCMQrQBNdWqFJ93nzrh
gBzDPFcWSKxMuyYQOa9noklARwNYOrd6+JHr3cVcpXFEh/hj72UyJ6ZORyhDtimY
Tm9Z8sKnyBA/fCNe8tJSM8z4Wyh6OTezG4BrRLOg++rBCEWd8kLOsMFzRqqCz/ud
NHwX5sHFbAgIEOp+VwX5aDhX9or2BpawAFcID36x7TEqbShvc/6xdS8nN236r9ED
zznSSZzzycTwsBa1iucEGojTj+RKMkd+2jAWd/ANJcNnn9iYmSZdnl2hJjPsuDi7
Yyoh9xMvg7aPMHtvbaPb62q4MfZW/AWX6uvTjVsHur2pPP8ppDy1tnTX0m7lh1/i
HqblyCT71YN1UwsPmJjZDB4wMnIGvr362b5q0LDVtkP3NQXkPIA2GTIE7B3TYLrq
LAc4TYgw/Lgpz9yedzTpJtDH12L0JQOayNEnK/d5nBFMvk6j2Y6KzGqxag4391TF
7vPTvyO61FMzJZmewbPA6aiwATmj013NaxhyaBAgeriyfjVjegx5us/zdwsvD4jD
kJc7P6GmAPOLPY2nzlAUgVqn5JW2Qy6EFkCk/LqM1fdLqLTnTfqajuqVrbq7l6vh
Y0SF4lK1uGa9nC1ggb7rHE5U4UJT5iYRiz+Av+PToBdek6qOQTtqwzU0mWnFo5r2
fSclb0dKMTP0MWGqeGmD7tspPY8bhKR0Y9SeGZxJVgD7wfHbaFpFY5NvIUukS4zZ
QNe4/jpd+sPIXIKKdnZ9L+7HMUfM/toeEa1ohb2MZmVwQCtyvW1lGSdWAnWluRBk
QUzXiZDQBM8SY+RTTp/R05BC7lUTyFfLH16hHtBuo2ox9lSbIdX5ENfm6Tl3OrOt
S4u2pLxc6Gwp3Z0W+XowQwzmhuqwuOsLUHdgl8KSq7qF8FpRZxJrn+8icFtmHFKF
KZpqngyppD27LdGwcHUwHHcjpjMPxxWy5BTibBTbLFFjQy0MoOIC7NZfLdUiYN1W
ZhS/ihJWF1Lblp3yw7cysqdtf4ubwJw/rnYnmo1Tl7ihKfG3pLJuT5aNHW5Me7me
lgk+MN1no2BYSoy6CPNchzdT0gM8r8kVaJQlS0gVaSX9CC+h8jpDRm7wAw1YB/gc
BoAW9CozbiktECPBWHtcHKm7zvM1ZEVISUKhEfCalT4ZDp20nTSCdNGM2rJGg6LZ
f3qj+V9G/PG+cHP5NqUe0PUWoRi46RpFDaDzFX2Yflnf9Eh0tOf1D7/l7sUnM8PT
LUK4yHR3e1TOj/BLbhiq7xjl1zcMntQx1ghX4i7yWkjDVpQcx37xAm1ahjBRrKfK
WMzN2XYQiqzBq1ybh+Nc/aw3eSG2lrXD32fGpbnDvuXZOJzZjoUutAxC2v5qM9MP
SdVJboA0QoPQtNS9c03vgf/MPLcjwlInzWIv6S552iopcOT50/2l90O6bLsHH35q
Zp8dVWG2n2gKE4yrzWdGN8IoZpmPz+h9js/IFgMbDSGy6cX0/nkvQMmitfO1Stlj
rSXAw3ZaQN1mx3Lh3bFIVIRlGh98lJQpmvfvTN3PUT+pCwIhQrBoUIIWEqsARRo/
4tmh0e4Dwz14yiZm+KoOqnvx8qUWpk7c083/GlnZa20xAQkgUne98i1o9ZwGl9in
9z+sLa8QBm3BKOBeNB7me4t20ARKVRZH4ozS7/oD6lca81CI74dZ+g3uOAoQ5Il3
7ewpieuGnI/Wj2xlrQTiXUtpYAgPSyuYamW+qU6KiRes03fps8UTXmF0m1Y+6F0z
6n1XizZCEypDlDItRI/c3nWdF7bHZ1QBkO9MTul2XWzRuvf+/ZvhNU7HOpy5mLM0
lsrR1uAXEmBQftf1BymiQUvARyoowXSA7evKgM/GsnnNflDposj9sBSISOuNkrmb
hgs97VTSArOtbp6WXZ8nyrNMP/D5GO99FRXjKJNYncUWy9Djo53B78tPgivvPyxf
qcXymXOsNpk/Wez7iAtFUgHW/lhvn/Py99lWQqM3hpauaK4J33EKVD/9edvyuYor
cnnj1PIjNP7w9m25JPHLbW2Hl4k4AhvCQPFfABF2CJFaQKOl7ONHLPYV0wIzx0Yo
YaGDwFMfk+dnugbcjO+QP5BOuGGDSDfBW2rWqqq5H4zoQe/TC9S3alrGDPzV/kIu
GCCHyXT2NparDNKPzKySlz3S3dXdw12owdjMNwD11M/R1Y1BfPiuRLLIa+u96pnW
5CaKNkNWw2iJMkKUE1mUhIWXlGaTsLW+OvljvBS4BfzGexBVdUw7id99qGZijHQb
EUcgD1cIOA36Bc0hqiZfgKP70hvDC4VlbwcXKbmGugTYi+5VeVfe8rNSxs67/a/m
2rKzcLDXS5EdFwK0/jHA5ASLgpyaCdhpFa3EHkhiK9uO95bjBuNU02RQWImfh1Jb
fnxTo3FkN/YSyfgWCUD8f36yyX/GTaVgD0DvyQgodb04k5QIRTdGxsBuwGmKlCYa
zdiOgHbEXFV/UpWurMkuhnWzVH2t0nzpmRfzrkGQkQEVQci+sVv8h1bBooWZALcn
N5Avv5j0ND3NPfDjb56LbT2ye7v8EShT6Caai4xm1A1Aa6cNQ8dMU8jUefWwn54c
lFNTrxYQy9IOZIUSWLhxKi44kHfuz76/VN6AUdvfj1raZSwr2CL61/BWvjw6UWW9
oDZ0fMla13+ewzqnFOS1cGqQvEZ9rI3odXlq+RRm6YGwasJ3TWvCpk4wjBOM1Cpt
x7Fx47cmp5uKnN8D6yeOlqQgB2Aj4oNCMX9jNC8RrAVds50LLk6QsAq4Z82FDsoT
wT6riBtRw5J9ODX7w0F2Q0TzBD8mU+EDglurTsiqqCJKFqH4sgQUE+X7CQJIMe3l
1ellirhdCJbLjERXFSu8aSTlQWI0cJ0k2CVwlmrHQ/jipLcJ6MVtB+5ExzHgcVba
nIfnTJ/s6CyFMb+rz/z+xtzKQWczFvntMOCv7rIscVeE1jqpTi7doz6HRx8bvLCn
ChmoFa5fIWUn1Yi29JAD6lM8koRB5dSxOvoi3PBXP9F9hainJ8iiLkwj2Uu3Lx4D
sBiOFjt5NadfbNqJWO3OGt91e/iqvFcsbjHT+nbmNqxDHtcYALgGJK5VR8n1ewi9
WtZaMk27uYS9VMOvu2VcpjVfx4sOAuJqAv/s4L6SxElTMRWa33FWoB6XN3eUCiF6
v5xcxisl2fkhfH5uy1/tP2naO6AJDlLdG4WGM9wdvmTObkaQj+qLiOMa5jEiM00C
T4/VMl8ZRxIyHRrdWJ9cDgC0PMuBoZBtJ+y0wNqhpxFaPFT98L5SKQxOeY8nY4Iv
Y6ItuoiKQgUHaWZ0nsNyq0t+ZaQL49HWdSHNQt5hTjYNosoTa2EWtrQc36dpdgqI
shcXqjxpdYZnbmcRQ5FnXb6Pu9TEByYsqhkLiwbfNMrJWprnGKRLtp/3P8m2k8PK
5/4/cmr7/oJsrvJlOz1ROuWvOZfwllFKlG/GLc7KXbSOlU9SRioiHI5SgCg5gxz/
/WdSiDqsj1zdJPfoDvSjB5Zr9eijACN/pnSMmYjmyHX9orqcv19bkc7xb37EwPf7
LO3xiUoS5EllGRknoQ1GXBwAZWK9E3FQE30FjRxHG14pX30L2FGcuraqRW4ZHUVa
Fp0xAW5JbI0EeZOOoSrQt75lw3Ay0raxA5boNGDJLvoWVlMuYhN/CSTMHGAzln2q
YVf4j22DTxHb2cZAOGZTDqFVrCa99Top53nzNIHDQyF45rJ7HhtVjPlfkksGvNJu
vZL6F0aXfgjzJzajH21BqriSWOWIf9nAgMd1iD/qtr4hX8wlhy9UbXVgfVrYtZ9K
JjkUZ7euekrZkuX94gybhFoM015j3LO2gNjtqv/HAQH5PV1cItyUdtG6yNJW+njD
od8nMfvyrlUCmEniAk7Nte19UNI0JGQtRNch/QZhLK35FL1KOf4AMf/BRg8GcwRQ
z80JJTnOyhMSumgUSNm5j2J3fbQ0kY7Yk0PHfrAiV8wb8bpNtAKlpovIb60bAkZ4
Zna2uvZySPwQWZHn/00Rui902kz+qOBsJ00wubO8TIP6qf4FuyxS463yf7DtsvVv
9EepRtpEVqxdBm5KpJUitd0TeJ2Kz4pKAJXPU7+IBCHLZcyY8TQpqTkUlSjcMy2H
Hx7c8ST1lKHVkYfvmx238Tl6xhX4Ly2/ZW7Up8WyAhp5Rty66En8Mu0woz+P+yXC
xCGQrk/bYftcNHrwzNxddiuBnZq4ea7eA1caKtfVhgdaSK/Rrkj049gUxGCwlncM
fiQpqxJcAYy67YXQAL+LUXw0fuyTre2VGLRtHWy2DKNb38VFKXWHeGrBUwHMCYHV
SQfUFxLJub8LoQjAlDqoXO7O1xk+TZYWMILMqcrkfb8vvkRedUDpYZZt70oWSUoy
CtB4bJP15O5HCgkMuLkUAisAd8jLk/UeWqWGhZDoVDDMUefc1iqPxqJ3rFAneaBV
km5So3SntkJ6n4v3XLjhODAnGZA7IzNGwpvfd0Qovckr//clN7DFj5SG8pWceRFj
SolzFu23dNAGCPduyyfp8JnAxsqsMkNRVEsUcXpFU5n/64QEsfRuhX8NMc+R98/m
DWJwokxAB5l5rBX5Vho+VBT4Lad+TKhvwvroFrv2k+5qVbhPe7MYKjXpC56ziZ2l
BZZgR7j9RUEYo1VNpf8S1SiWPDiOA2lndU+qiHG4m4L7/U36IUr63FyvRJEQ8cPM
qNMkesKi67t6n/26tDPtGv2mDEKWROR+BtLzRBY3G4fEM5yLTEW63CfwWqnlebxU
kwKuP7QZOPCZnKqLDFRJ7J/bHr5ArGDGcRdruWWZGENtbD+EGN6jFc8VXfRp66UO
jDo9q6cgmL0twIx1bXAhkEmlAYcmKuPMcVM829IUcB5yMGtbtEp323epB2e9yPHp
UdiIZy/P+Ks2Ft3y/fv2gJlcL3AK3Y8GluEaDaSr1YmnL1TO6CXJHe8erHxbLznF
ULEO8L8TSHEUpgxcsIRma3mV1fUhXFN5TzBE3Ya4hfAPu2jgxk9yknBwXSnIMI2M
psZ8EZcMLC7nrLrqlbjfBj6fRHp9hg+tTEehdLuMsEfsSKXfV4xf9kdsbRV3k+ZX
Vi3dYznJpr5UlDVYmre8X0Pjym+qgDRjkheeRvcFXxyX4cObltbMFnBtvz5XeToG
O6QdirFHoRat4bwIyq0rOBVhraaNHR2dW4XqhH1AjL+duY5f5qIUm8N2xN/ezjUl
AkUsXifvykSxQWyDhxrIDT9HZ/GZHRljHPaAzO2PgqS+Xcz364dIDgzFvVSnmEAA
gytEa6DfETOOnrjS1wWuJ3bW5vXqHMdOYAwifVeTNDtEMrlV0V1yZr4/jHpz4byu
p3y1t6uWGBf1N1sPIvRXolQjDqSejrlZJdnQtmsV+WKn2FHs+Ule50YktbGwMJ61
psEI5WvJLwUf9RbgF3U+k/g0U3RHssU2AAnzMwPtMkzig2KT7BrjO94NRKN8lmon
ujqZIrfhowQ6tHJz+hGPvkTdqeYvzh3J9uUOK4QRvxmTyY6NoHtqvCrH7vM+Dw+A
NW0HYjEB5J5hIPIBj1HmaAi2P0joszvtufuxcSl0zPmdxVZ/YLo6pyARHmKf9AKm
KCOTBecuBId4q7gX43hy2wccCpH9VBHswpkHaoXzvtp2YH0EAqaxcZl5nPojQD3p
B/Txnh3LYI51uEX1MOEe9TBIGM2XahZ3bVtpDATbZu4dF3dLy+thPJ/qfTYRuAfx
EXeOj3RZKMyRDmi/WAVR0V07PmBWF/5WQL9wuxD+AsMdos8r0cosTc4gRhOUeQXH
d5Pags00xsGa0ssCzD8K3Hs0/CniuS3NQSWk2jtIONljgZEKhQDerGfplICx8ehv
IqLBfYn7L/SQka6ZX/xzvnB87OJF5JsMrRRqOjY6yhSQyczS43cYAPhKNuck7Z8L
ZUYUhevZtz04jiL+x5NvuYmibtfGrH+o1r/lxixHttgnGOJceriJw7CV3tRCV9N8
Hhi1CGvSOReGD22aIiZR7zJ7T+Hnr6E+74IGBx61uGyM83fD1NiD2euAXuLYLwGC
A4k63E5rSwIh9sK7GK47js6H9enmBkYyvYH70227KY3QClu2RTjUwIuaruG6awLx
zpt1SijVjq7lN3qUmqmnPfjxrNryunnx6JXbVzs9fDKdEpdf4HXQKYB9qN0R3SRv
XiL9S9buhj3/PU8dzmb5oeLwgHaV2xI5vAhr9w5u4I0oOABgsQoErO1jS4k2Y9vx
zkEEV1UmO0r4xs3RSH5G7z40yWCt+n47YPBwSRofhxUvkVKcqVDNLcMrkJChDGUH
1tr8tJV9UWtK4/Vyb4ZGH8YMQIParQO/rHUuaKQfZNxUmGEIkiMYDH4yj/eUkezL
WXmEziBorJ243orfbi4CZpCwiNns0+BSHmSReIXxrXqEKCRCOScUFW+Nl1fxoukh
5BtXHWYoE302urnkDvX8pQA1vm1RY3DpN6AvT0IaLYQL5C23bhflLcuTE8KTPmSX
F7XrgXn4Bw3vi2BGQBoyp2lL6YSlB0PAJ3SEB6hDVZOXrRneK3qUz9DeZh4IkOLe
Yw4yS9SAW0UsaGqLzVJFeFvlqbAcu3D1op6qdl1A6FkHWQjrk61cTPeHYziPHN4N
l+jVldJA4QtfR4KXt2KBi5e/MvTTaMpB2igMmfRSVAjVQwIc6hE3/5EFDxC2pdwI
43lElG5Yy+I5v7tZZoya4J5P2Vcbi3dp82A84mYnOM0ctQI7HPzZXFW/+2VfjiI1
esmtqpkhbmDDvXZ6UMk594Q2OVpWzczPjDJrIxLfkLbysJxk0kB/QC6Us1pNhgvD
Rdxtwj/1TGVG+OdRv5tE9gTKAoU0Tfj+dk+cG2it8YrSZBI4DUmnxK4FgmqbmY++
RgkgAh/M5fGNJOXE2E2goHyJhHe+TyN3bH3/3JgOYZcopniJaXWKQAn+0W58oW1w
AqMRwsYTLVEuNVox7oup2FkkMOEhmToop2QzK9gVQLIQTJOzEkUwRZv85bgseOs9
VcGdPdEXvLq/qsXOGcmeFpZbizkbG9RB3b1GSYCQdsMEI4SdtG7uO2cD6B5UHIzs
Hpf8i6yjPuJ0GJOEXSchPKRpdb/TfM0/dRC+ww8Ju6P+FCzMFdDRnWprg6sypFT5
kXn6i5ehcxV5kktawspXBtjzpnPcfoZO6DpQbeT+iwwWS4V3ZNrV62eupD07qVT8
UFgdWJ7Ywtv1Cqg4dVZGA60d44y8+6HjEIIweurVoMbOH83yWVRk0K5ipk3RMc68
gX5lsTiSF1IIKyr4Frn+XelDL7wHE6IlCkZPZKsWftnjYeSYlcqDK8IxiF26LMZo
nXN+DAj1yYHVDBuTWNnL0P4XvMQi6mXW46IqFZ97zhqeUJ911ewVcoyzSsoRPGTn
zOB8MzVafmhxmUQVJC99Pbkn9exUsi8rI3y/uC2U8cLD/kh81933MrAxcxir1Dln
tOeKTEAP22ec9I4XaBzpdz4mn4XnYoTY2iXNSy2eJ0A4SHC2pUA9X82xVyLjzG99
qXATGzJ9C9hy14xI4SuIQRUuXD7BrVBFGb6IfcX3S7Td9PvwUhHCkeVj0dyRieOI
0MjCxC+9Pc0oY0izL+AF+Xnmfd0MhIMvI6S/FSI7kNhARv8fPQCpO4HCQHGDRoWf
ldkzYNriWldU2bwpEfajohxvBOT0Xk/6UGBglSIMlA4B6MKWgT5ppFY4RlWrV6RI
Z1k1WrElLDNeUiAzfvcELkYGARGCRVyF/zpSVQVSvQjGxeeNDmQZyuNUNNwZErCF
6nTFlnSsXpfWYAWWpMX0MwlMnA1nBCnD+f3NPCLJsOUWOhwIKMtO9TIqgh59/srI
qlJVVyicWBXfuDgCJ4rTowMsqzZvxZGFO9VxtyoDLheUYpPGl+LAVLeypHAYWTQs
YFMrryZD6kUL7IUmGoLOjb7Vd8FZDv9CuHySZIL1Z0zg2r/BZeNoceQt5nrK0iY/
k3JVtQhZM9PrQhJ4OlS8fhYhzWqKza35gRjiLCgG9/2o1KWDlJlLwqNiVmmLAoWo
gCpHlkgmX4x3TmbQ7iCwyqla/FI/qNZZaycvx8eBGq49Q3VX1y+FLH6uAWU1kYso
Esrcjipa43YjC5CpbFvs2EbHtuGqEepd526C3ECygjfvxuC3BRSNEOTsN169Q1HL
H718mLIETDW/3xrTlC2GYTIBCbOR1P7dm1GyU90gsrdGCotHBFPmwdH31jw8ZitL
VThW2h3efhOzj/4UzNrCIurFfJTv4wTKuIIiC+DemjVjdVSEJ15bbAs70RWlsiyG
Cv6UAgF+lIxAi/4tzbGp53hFofwiuC3m6iQ4ga7Kmjy+95vkYJGOgG9hcz3nt5UR
ofTvzbbQmm9Nz3YaTSDl0JPSd2M3oZxbAC4ese1JFw1+YY6rJlaodA47Ydds0xeb
0X5WxHUpES5L/w0USI27GTDFRDBzDG2W+m/6qmeFxWteTM1p56d8T8gwQzsqsmOK
j6cqt1V0eEqhV6xZeigJ6jTyhLBVVNAj9ntkJJZk8F37hCFAVYgpCAHJqlXzpHqA
eaqUWWC0LGv5Nnx05TkuQGnueMb67JLSWv7uP9D6pyf/BxwBFPbPISEYwXu1d46s
/OWpnTN1f3YElaUL8wQDtsmrhdtBhPLAEm6lCuR6m1dhDCNPiN8DYZ4NRaOTBufB
lte4waraJWZBZb4xnmilFTiLvlN2Kuuk8l+RbOkP6hP7K7Kf/ufT2db35Xt8Fu8W
O1Pca1AUnwQD4fKt0Nwbm1sby46g4w2kjiV5R2jpf61//bRxNKJ7a32vXJr3Ri1l
rfsdhKvcbVqE5UKCKc6kv+rM9u6ySAITJgTRb2np5YlfmuXQlKSiiBxlSbDdHpp0
MviSc2x7UGQ8S3or/VF2D4k3q741w6tOY/HiVZth8O8kISA1W9PMZIgpqv+gARR7
cqxFAwfsCG/BiiQ2ZZ8x9+Hf1chUJyIGduZkGAnzk4JmC/QM/ek0OBietelv5nCi
KqccwAV+wJSCDK/EHmGmRHoRZy/B74QcQ/B+KHJVPiwKI58UzYZB+cDY33mhcEYw
2TaZPljozebzKCaTNdkRruI50ZcYzPoTg9hZFHmtjZTw9iQxIy4dZ6UdDoxsnBhd
/guq8aOWpBNgbWQak8dILl25bzuv0yp5mqk+q/8ErsezC7eSa6p1sKUv75z2yiXZ
Ftcg+Ohy8WK1+pvmQ0IfDQbMoDuOzJQgi4q/nyWlRm4CTgqOJX4C7Jz9fDiTUIrm
vgpZRfWU01U242+wRBcCZrTqJCkURKE421LAuKem7diEGmJpyekg8NglVZI1piBp
4ofAGYCEd5/S6yvmaBgT9pyD+j/uCYulLd1nu93KtMzYG9VJBtksdGtNYCq7IA61
3cOyZCXPJCi+V50mh0wfJbSgcGdhQNkM+VvSALkLp7jxaxZ7i+jnEEGEwlJ9l2U+
FGfk4Z6x6XlUhMRIBQ9nCZmwqklp7FeWCJnuvS9YDaXZDSe6jFwPZB0fi06Oij45
zeiyqXsuhAEQpThg0hkbKPx6/Fq/CYM1u15L6ZWehnMphqli2hsqqnCVie2C98NO
09jgXclgWEuWEmRtTMYY38Bx8z9ujqfpYP3DbfrBQNbMUmF0m5UkwFML0JhdNUEy
Opdt4tnDfLD8doEq6k1uCJQ1zjnTRNi4lNn4sOg+aC211lj39sF1kmjCK0E0iS2l
/pIBA3NjmWTKYReuktrM8uoKGlqy2HF+2o/BG8sqUXywVfV8HmzuSkQeNQNEAn6M
h9qoCsEMkmRJW3r/2ycAAYpcH1NWAbaCMmOiX8w58LWzhu1UdbtJQ9ox9NUlJycV
FNrux2GR+cTHgMpXx/vVzS8+VdhuYMd8VGnT4IXK6Zxnm5u38mZ8gEzHedvVq+fH
tFaSh39g2BQsomFTkHSIJG1u7QWCfLNxMqP27pgc/CLcjclAEcnQKdGDKF09fbkY
OgDXRQd2Je1I6HFazUZG+y7eKvLoVqghrAz0tPXU19RayecdRF6UWvVqml+ZHGu3
RfljYO9wwJD3hCCMP3jF1OEeTyOPeD1CVCGbqPenD0na8i1SyYFq0dKqvf/x7uf4
WPOHDpPA8xCjNi/v2nMOyMINOe/VV7oRCM7KUHecUsHnon3bmya7PTEbRFjN0hNm
7I81z/wAJzPy4UrclSRqXmPgPjS7GeGLp5gdGqdnFi11FSv80oe1KmwhHvYDC4Dw
Cwy/f3+MxZsrinO8SIP94Fxuqp7njiVYP65mdR9Ol9GWUSaP+LzDckvODagn4uiw
uHzrB9dUwrdV9lbBiDolb9vDO3ILN14yZFTxQ7/v4XqpXbyc42AqsiCQkRs2TX92
mZww8hwv01HxMWra7uJZCbwDRlJCEIyOQI+xS/BnMkYV5ZyXwER84qSKiIs3ZL51
fO6KVZffkRVP7YPG+zxjhMlPL6NIPhIeTtmpEMQQnGlE2r2qsaamM3e6gguZA1or
9MlUap9IkzJKX3xJRY8uc85y/QNfAgiuZqiMQPQJVv7v5vf+zzDiNwdAlAyrycax
xFpdPl1/mwIgE3nUAZh6GJD92NhCQEvEva/2UiSfvpH9qyX4ZrW0Gv73TlQgqdgY
xLf7Z8SxTwx7hVMSfGC0ybH1hLwk7s7rdWxCgQ5TnZ5bAtsGTEZ05l8h+dTfLk4Z
GbNLJH544A0zJMgY5opKpFn010d7lYLah1VPXm/aTxsdQphskqTPcawFe66cyGpJ
jTSEUw918W8rkYqIuWGqXHLSF87Jq8FroZE9V8sZqVvVh+zf7oZIM35uZnc4rvBU
LvVZFDrTnJxZpG/rw7RHh6DNzjDXOyLYWqu0sOgoaKMRF1HSB8YoV6IsDCRoMCKU
38r6Wo1/aLx40gwYWxI8r95Hk9w5CvLIIA08Yz4pcyfnd2w3bppztXU8gmZjbxbh
y42NSKVV3MEo7o0iCNEghImO97U57Pw94IXKyxzfwpy2CMorUK62PS+IPxt1PfTU
YvrezznXmZOYBSZsBj4JqXPNv7or7029rqwkUWfAHeZT5gb+HlYFhqBYJLPO3VRp
sD08QeKm19dJxJoMUfAExyYkclPPtyHQBG8atpcSXPG0LRAUIVgFFy33ZI72fRhv
liPROXakjU+Ay4nuQYSRH6o/X94tSGt6cze4sJCE5alWlcK4kby9Up+L78l/Jeob
uK4AstUtLkG9Gewjt0QuC6fXOUO0Fbx/vUN37BZU6UZhBBns/O35VIrv7oLol1vb
/C89Q2/JyhzE/w5vVK89rFz5FgA6POQVOqqBlQzaKek2o3vWuurWcqfEb4dt+hFd
r3y10E+ho4LctrL9sxSLkMj4WSlRDZeP1f9F5J4xrvnp4AwSMIymMmpGG6b+xJzL
in8X0xWQ4OZPAS6ERugar2vhboqWrETs4IO5lidonEqC/Y1AZWGU2HmnoxS4/Wos
cg2XpSbISPSYwAl/w2E3teCHjj1GWtss+IOdWNtZAhaVEQciuBjDjYWJwyRKuzDd
Wooq56tmxjTPLFZESgIHbsmlW/H7kyuc0nvbjROqqs/8O0vxFsYGkHTtGEk1MMrN
Mof9cjQFJPFFbpobm7kG8M1BEmRHGP3KlLAurLffp3l6QNTp359Jc2O8O56VmOJb
RkdJswlQaOGiSy51NJKcqgIGe3Shm+sebA6dsSCUgkrn85QJgskxljtO9DQUozGU
r+E4VCJptIXFrocfnRti1II9KUgp9ZOnTSLI5YWvAO47TH8tcy+UTDP0u5KFb3Ed
eQ+++a/6n5igVEtPdZwOqos+VMLTfwWc8aZqCVVYQlUjO5V20S2QBtV6TPILHBVl
ICj7GqfoaNUB8/BL+LX/hx+zyq9unTbGYICI5LmX2g4oQiwk/tdj1kzbJQVwE2dQ
lXd/Ib64VNpS03LNihXE5Npd0HBQ2wsCpZI9MI1HLQW3nwKIGKA2+4kv3SnO7HLy
u+nt9z4VheHCGb2iC5df5P3NdrrCaDMsAakClEbYU2BAe1tH0qrKbwk72FS0gy7S
vDIMxFJsIMOPyTk4eTgaDv/1Zno/xx5PUX1na+kPQkrTX7x/mUigmQIRBcK3q0nT
UMivsw6o/JDFSnuptU6MOl5YDFoAsHWzCt5r/gjxz0sKR5Q0R16+h/OIrGGIg3Gj
rM7Cpi8e7kyVH3RHjsyGLV8v9AvZw6xqq5QNtVl3euW/3CWqKBfOS4JwPlS0vbDh
8hwcV60TR68UDhXWF36HNbHDVI+A3xsK6dbxDs2ybUqgGJn6+kJfqABbRdFP2WRe
Qa5QaUw01dJDwAnFVsdu8qWyNmU6xLjFDivSy2s+hduBN8NyR72lnE5oghkc5lPz
7p1QMEjkuGUwd49y0ZQHyT2jS/3sItvw0oqdyW8iRcVEN/2ZJ57IUhNQHnxr0izo
LBfr3GxR8rR8dFlfKMpCZPklyPQR0THrMPR3s68ZY52dA6Ad3+TMTTFuS8m03Ek+
0o6EDBKdHdc/UggWfPvFfD6tHQmgrh3Xxh51GKvgJFfUjWfzUrDnCgAWZ+zWnMcy
PsqKMwtQK+GhGKJfNL//L+7azRriPX7tNWsWptBSV1/xr2HuuYIf6dhUKDsu8dht
dluEVAh5IHSsz5phhVpSLsNX354BhQQ5H6qnkSWdo79Ut+un0nPfOPGX699EHwJ4
PSkcRyZx4CP2z8/jp88bNK9oqJGaSdTZDy2ImkoLIICHYHwyPbDVjgOAi3aYAiJy
azT0T9z9cc+FIlCk4+ow9tgQYnJqGphCDr5ekAICz3PldHxoE3lluqIc2QtZumjR
U5E7kijiBxOdMSVCLoNEQ4SZypwyMGrxXRd3XA2S8A2axjSInMs0ZzH3gdA878G6
yL2d4h1SyDh2nfURoc9kZCjpQs77ceZibU6iKeO0dPrZwcp++HdmuzFD7td77/qD
Bf7p1uysDupvLpRlLOuqMfpUwBgUQG2gK6Vf0y+ZCnozqYHyv320YP+dE+O4eYLS
po45y9hiiul5esVhgFIoC+5Nblo5ME8QYXaF7ITXlLfqe1HqQKplhvpD8zDorp3n
+I0fp7jl/FUrAEgl3KrJfSADtwmgNWIVAhAAKGD7H8I5M9ZivFDVWohcfGdmreba
PzIWrMLVkg1L9hv7sn8yUnrMKAETsVMWuYqmvaCS1/oeQ7LVWrjpk1tDWyfX0Ksw
8rbmXpc6Fb1JmV8ITjDe9/6IqiBjMbUUklG1gcnID652IGEGtXDhoe4JGS99hgDd
sEn/g//mNQ987V2H9b8F4jPY3O3vWmvaL6KlJCbZn/DmfdktPEF81RBKKpIdGEaf
QqzYRXUqLgeKBJC6TdfxvQzuV6hpJXJ82y0RfA4uCOEBsQeJXAfbNLX/gbmxbhgm
3JQRBeTWtT1YZLJJh4F63aiWWOZv0hK0DLmFTEVJdZ/79U3OaoeTU+Dq60uR3SFJ
HdWNa0yk7xOgTM4j9JAYJRYPlwmQxR58KDMjBs6vDtbPew8DoSV4+ylC+pLYhp9O
9VzrlcdZdr9kd7cDVsCmzXXdLbg1m5aJVzCEzVBuQCy8x06ahUZDz51X9hqyEb+9
1DMshTzLsBKjF98351eJcymUeU3EqxKuFpl+9e1PWEfP5Z7Vd3Dk3qD8DzqX5G1X
vMAstGcGpa2xziGN6868Vd9I3RDu14UuU++bsiEQDtznOdU0y7KoE5Oshx9bB4LX
JFklMSubuOav0Xzbl1X0jhlT7HXL77DwLLNeWGBuXQC2awJqnIQ7kPl77l9t8Jfr
NZ6mXD2keBaAii3+GD7mfBYPl6LpfL6F05fhNIsgYjjceWIUXr9PKD0YjGalRJDh
K4FuKXPswSVZqxEdlQTGBkjk+yiexIhDw8qDrVzslDOhLnLQqqQIHH6AzJ4i4xkj
sZqBFJOXMDuK4d6HXGWbVB/8hn23uoqc1PzIAcEtU8tfvdC31wCpItnkQrx79lm1
W51LfDeaKTeC3scxeQFriSDny7J5RuVoNAn9EXWaIiPtLO7Ca+DJB+aUPnM62X4/
YpzfKEXsiPwJYdCwJgoI3V9q9iFSZVMKEKWhSLsBWYHP8cJ7BA9rSDLIFBLhaHyV
g2kcee5zo1RKECX5tIwM/YcwyNivpttjzk8K6JQUJ8Yb7kY5KG/MTUL55mtRslhs
NMwS4thLbUOP5lEm+No0jDJDrUDdhmsiTKzN34L7EQ1ZGP6t71F4rzDx19JTqUaw
1rSeZyYbhTSOmFW4Hc4ZNraF3FCkPMYcAhEYBimcLCCVDmWX/Du29yl/gHWLjre8
N16xghhjUMO6m31xLaOt09jodFlg5N92GRLaxXI31Ac8MU7svhwIOCrTWpN0OMI8
tIImOUx9QrH2lxFSkNIO+9mo0cFbgXg2IEQJ2KtGPul7yhAqHyz+Klk/PEHx3PB9
p4qHAdiU2HltlBujXQl/amVizkpuuukmFL/9iOu3Vh2SSw0MHqbKggZkTCNge5Ly
L6OdlE7IU9KMjcE8onEfCo49+BaEEqhaHTiY1C9IwsUUzW2M73eWuVbWsa6ZApbB
0gZcNuv5PqUQKt80rfH9owUGHKvYgavOIcZAVVKlAnUdzBsOmMrMLffTRLy/Jzzy
vbVryG82vzPr4WNg4QttQRjZznDPzSTty3zw40rEOq8t7opSDiWO76n7vXcTsrZ7
56g4ZOlbt/SLVuAW9qbsDTNJYE2GEF2sK5RBcT6KHn9KuqSZuoDN6C4Q11jiGDly
2YBvXAVQjH+f/2PFZP3r5ourJJEdkgHkJ+ZSZTuQSXMH4AosCsZisE5zgXw49bcc
7Qxd7HGk9PbFozNxTat5mMNKDPcJ8Lun44EE4W7DXOq24YncUbfwAIRiN0g3U7vz
mRZ2IDF/arxFM4R5x50z/IEnPzQZlOKeSUP/TDLd8ARY5BBF4v8lO9H4zSd81DPP
HPgCUqiZnohicAlnWZItXjWgR9+8/V9RRoE56w+QM8YkHh8cRCS6fW+5MNPbk3ZU
N+8sNVRpIfOhhiia6NMLR3WGv+IiYQoX/7rON2XcZq9zJynSxuSPwwcoS8i5P2a/
NJRtr3uAAZizozGdqYtGFu/5P8pWrGUpINIiH9bAqIOFzHieuoWyY6j1IzBE9HNT
zBt81jR3sVkusCnjN7KGCG4dbvVqbAzCJcCVXztnw4GBqq8K8N4u/SVrzfhmRvhq
eeX3SM3rygTbeDRYhN77v4ywqevDRjp8wQrn5Kvrn9pPeMvKfGngXyMAqnkDMUmK
zqe3IEQDkLEKE1+PJBb87GA2xXa8IOR5vpmQkkTt5jyX+tBwU3lCr/CxeIIORhm5
ah+bHc40i89Ua8lDF2vJZ8AldOYdSi/7BKv9ABpWedkGmE1RL/QOYtlLmRpIueuI
o1DQtMyYh3+l9uM8ja7nciPrSgx6dKHGgFqlufoazicIxRpMrJr/huFc3vHYdfGW
MLzaV/YcOmLDbdg5CNhy8XD0BtqhbpqQBksSGyheO7aULCCh5L8W/N9b/7DXjOGR
KAM8t7EE+k3cLC7x8hft6xo8IDYk4FfY6LAX9MZWdn0NflaDVmPS9uT3F7MMcRYa
BPB83viVOtne9R28XIUlJgS3EU2TE2EdQpNtJH2rHizRsCwUM3dapHaEtRKvuIap
Iy7Gs4SO5cYhQS5KX47wL3DhNt6LSkTJFFH/T0caOgwHpu8UkHnR7IyzvE9UIDtn
cckA7cmg1yMVIBGpE56p6p96LJea/Nr+3CzTcPjfmp08aQH78LLFPdNUXCozHf2Z
PpKL5SbLPT81pRkN+x6uTt+jdXRcXaYuAUAH0DDor7T29uYgGG0dyv8j2AXppMTt
7hvue28BNKFzHBduijccMdCLmidLZxeT0J1Io0K9aM5Jpr7vkq5fuMurL1AntKkA
kXbynfPs0R9B4UyyhWdA/Tj/mn2ny0nyjlG8toUMsyE9yfL/1e9maTOx9MsmKUgO
M2pqyb9YhYsbiGkXCnl4uDCFwl+5ijx/wYxJ4yIbj8PC0a9QhS0bg0r9LbdjbWx+
VOms0WiePhDP5mZTgc6u1wWIU/5XZ/FEnk+/+wtvudPO8Tf+E5zmVyOMuVkQm9Jk
tJQIC0ENe89kat4vzoTzbiZLbH6ziU38cYysZxnfA1gi63D1U8biGEl15ZtgB9En
ANjmPKHRAcvpf1HK8Es3tpiFxwji98FBJJ9Hkru+agGUWKFad3O71GWlgk+TrP1W
uJ46JI18ljTwRVWMQTFNus4E15qIrBrbdOzV8RfnSkaHBYx9bW4U0kzgUMhtPnFo
IPCorxpS5hc5/LwGNvMKuK9x7QXkn28j4KBu15z8dYFhlLLrD2w52JcbjXQ2H7/X
SjSL6bkuGMi7aMeVcFczr25vkw2gqXtm1e3YSSdMFUY7hlR0indTuSn8N/4Cio61
iL++M00xC9dfT8k+7qkfeWzwAlISMtprWxpM3EO+xcxPmKMv6aH1u99tOTFhGQu6
TzLc6VXzOoBWNVDDb2A8s5c1TP0irUdFazrYsISLtH9bdXyiHg1oi89nrwiND+se
ekOYyZeC3jEdmXGSEcfClwi0RFBtDFesr9cBfiinnIzQkzQWoUd3db8LjMrBQAG4
XfW3wKPcZ43KEnjBWRvdco7ud8dyEnODV0SYaxRivgZS3RiWSp+t9aVji/uTldle
fyTUsKmBQjF0J5SSA9ihp65nEYUYDYd8NGQku+ZrEyJxd9pnjSar0kaAweY89rKI
8FDjylcLx+jmg2G03mLomk1XjqpQf6Q2oCAnrh0ZhZT+N3b8ArcT53KwMKTrGqoQ
w/kXbydkGEBC08vRK8n2WN4psoKtDzOShT8JbopUePXyB5WYA7rgV0oQRcD/rCGI
sq8Z2A+JxDk7TIxLiNxt767rTkNqxZwBbDrcpwlXSteUgkJhuo1spCY0epfFJqbf
3bqDkMhcma4/GsZLMgOkO2i/4B2P89Ba9/y36hvcPsfqIbdoNxOWWGc9ZxxzHbWk
SYvnXciq+bfjRI3Lgh/jU2yxsrAIBJ4m16XfA4xuAWUryj+gFCX7teOvF2vsIbiE
qbvbyqt21LF7lbkxJhvHEs6Gvvm/Pg0f2QbNpTsQX6J9o5V9k66zswcf8K7iQ7Df
WtAHHSBFCFXRsCklLPiWb5/TV36yqXj43x+slg3TFj2JtXYcZ3vVaixQ/nszjT4s
hwC99jEFMZk4XNXFVvQtp0hcgV3cbtxKp0iEmKoqpbz/uJfWvs487AVSiotMJ3G+
2naCSLHMKareoSsA8TvzQIddxKcTcYau43wBOsCFkAZzq2z6PyRcCDk/p2PGXd/4
SjzKn/ib7eQQxehVe86N5y/mjYCVCEhMBiNxZn9aUlYonGb0shSRcpc60Z5Cwcd+
ajvnm1XjwqJEju1pYOsimTFLdgPvl9Ba8LRpDAvtu008OiRC9Yu8xctxz1MTPTqF
mrE+BApi1K28+UwXqWwlPi4u4+4BxhyLByN00FAJZ8tNwPF1skK8p6p3t8L2Ymph
RpkTVX6+euX+FpStAZEw7OI/jIo1DGGS1n06dYHwWSreXO7NjojhJp0EQ7a7nJpu
H1SrRCrxTf+5u/Hj4EmsKcAmro+EnEHSxuAaUHTBgaZHE+6AwsY/ewltxC3BeTNn
o8HPj529NOK4FVY65Es7u/AnT4kVjvoMO98kZ8LX8wY2I+3mwF+o9XKG7rnzugLi
nhj3AbpIozPkNo5IpTH17juobQtVxOcXkryktYtihRtCuFSNh9tQI/hNMrB/71xi
aigGAM2SBP0ItlO2ejTHu4zEEfgP18MoUQtkklSOuCuv/mZ+AIPSanJ3ta6M5CcO
4XX2Vqp3XsMCvK9aD+5OfiKf0rtR3p0zc27UDz2lohbzN49BVg8xBcfIUamusY4q
K20cck3nlN7pEZW9p1kXsj+ORtsQcf3X61SMBUnwwIpw0uctFK0lUG6Diusgwtgf
lwbM2JqzE8MYseI37azsFkbeHtPmo2NAwwchejcPBl7AWQdjVJW7W36oZlFmqW3A
w0BHEs/dinksRTWwdbLpe8Eai/Fop1FTRP1WHpS4qdw8RMMMb9JzU+/kk00WIMwC
JEscjaVN9iZtYSvIW2Mxee4vzvKw46OlQgOHteojfUa9OY4VYd7WuNO5uH2ngxib
WzkpYm3rI78UAlAxK2CRAjv7S7JvixtkiBQKoqxgnUOtLpmZCpyN7gUucUoXoYAz
B39GQEQ3uBZ/3EO/R5alVaHuwef8jvi0fQVmXznhiUyNt02XGKX7EI0U1ypAPl9y
dQtTsorDfcqo3+ozfPc+ApXiAJ+/4KmaMeEvMzl/2ypfSumw2RFA51e4tNiQEhJ+
VQ56HdvDy5sKmVjKw5oQpjI4tnxgUKn3udPZCIfBtLLRCfnYs4ovng5J3U2xm1tB
TcHaJYSsyduRyqCeCukEQvgXX5CWM9RmP/C1iCmniraf+B3geoGtFCRqFq91ILe5
t1qbVX0U9a8PTW4XlCvEdxzGfLyprFtHmZMjqhMJS2Rjba91QHVR62VVqkw/wolD
8MroACrHUGmBelasUHEDvGiZKDg79X99KrZje1cIalnrWxxNRSDWG60hL9liyqU/
nF/buGCYDxt1B9pjYJKlWANSHONV2xGyYrH42HEvwEXCaP395YUHrPLh4S78QVmP
zJIevNMQDjqFgX/GQBGMLTDvBk1a69pBd+xrCqC3Rmea9CPu27nCt8TL0pwKCH6E
Q1rR8qE+q7GTK2RMM6KOT5Bo2B2ePHRl/4QwTesAVIPjAD2cnMf9TRuDQl7tHGEZ
YqbrmQ5YJMjoUQVQ/lDC/lZ91/wHcEBJn7WcY7qAAlLjnCvdD/KrArzfIp0i8LUF
ovSGV0DURtVQdDwoolk+kcFZ1sBT+C5Iupeht7HEvhysVtFDRJNkdR8MeMrT8e1U
HqA/aB8qSe2xRLWSBtMutdF/OpO3N0OD/pX28VBcU3bGM1U48/7HfESxDag2hU91
qxrSy8CQE4ZzBvjsCjlb4zT1vlstKjV+bpZgUC/Q8gm+UOe5qgf1pp9IhF+x7Qz1
hhID5nX3ZuX1f2pk0Yioom2ihT0XXfU+lRpcJCjyADHFnPTHxAzbcPT/+UfkWV4b
jGW1tG0YNQNBpvZSrHhjpR7klKzkKSyBoiRfKjZASJP0L/CIns3OIzfSz+UuDiLU
+bGcT3iuQjP3Qp9csOhK+CHvcFE2FHPq/yzkgz+LLges4M8BW3uDlZj07AI5UKxB
GieLWcTyJiOdOzXi1Yw3sL1RDbd89G25BJqZFOrcndHpOz508S02hsiLxtz0Qob9
5ySDJGfq94ulQ4onZy8wVqhq3TJ3WnWeGUApsMiSdBgp9M6QOeZ4g9WZtVvPhsel
qFk49cAY2C3B+WpLlUVXlPtJjie62uWeQZBABUGQgb4KTmSxORVmQxKdvis9Ivw4
dq3hWFBSOu9cal4MRQRtsFRBikJBcflQlyOAH4HYsNFicUUTxFqdYkiq0vUyr7eK
a5GxG9auRwWlvrd/vceFz5PlGvNJ1fcMLoZdi1tbm31tO1FIslZFPxibLpK9XxCu
3N3NNPQldH4ctHkrVRrUM4GYjeabqH7PbXc2XwdOJIog3xR+BWqFoP3JThwQNZmS
G6nT4OuKIZlh0hw9FU80WJY0ZCfy8+hretXxP5jWdnaB7NOwqk4c0X8yiJEVrNzN
e2x3rt9WhK/qlBAm7c68e9lHAwKZWj3c7H8HZHCv13oZPLTxyfP4RRdQbT1SkmMY
abz9FugnzG8ifOvZ/W4ADPij57QCBYw7l2OTRN2EeF8jBSW7Lv935nJlrFiBQKAD
zKVsbaFJRCEfT+3LE5fDmKVQdTZdWzc0Ttknn2kxBxVJsMmMILRH8A64PhRuMsOK
sl3MJFF08Ozfs2kezifRifeZnbf29agdo5ypSsBJuPCVhPiDleDMv/Pbl3ldisVX
7nRUzQYQ6XfCgk6xp9xRtVRnXcdcSZ4V1RUXUNhskBu6+jtFHZLfWQf5cLG0U0p1
OKErXxkOAfwoI615/xt140A/gJHkx8Zs6tKYectofrhAiZZ+CyeO57dhQcelLG7z
eWj3R/4RJyYZCHuCmljfIJYCtXLEFR+1f1FquNoOUxx5DbdqhbHA5duC0B8USWB/
B617S4XFntIz5fu5zOBqWv7p6FNWvZMOwuCwgSJzVH2taFw0VU0AXmjv5d455xgu
E6apCXePy8Icye97LurpDE3hOFpgtSswsw3nk2BEshvMmNyLqBXExVP3haWSAwqK
b8O+yaW671BYD9YZKv9031wR3llAET+iUhubT1QNEzp1cwajy9+7sbUg1/AzFNIs
vO64jLESS+pQ7DMoR02gPEN/5c4ox1pqNFYjRlIaIdBIqu/AukU2NetApU9ts6oK
VwtJYEO8E1pNYL2WqrFlyTjRO3cRt/oMXEDHMEGmcjbonNGBnMo7B5wQd9PuO9Xt
PLMNKwzGMrTmrAr6Y/30FcbTpivmuTq6pBSf2/ONbMauF1wKIh4OODRwLVs1txDv
wLq2fujVc2DuVjvpgHpVTEyFdjhtkIEVld3/iMqy7dnmwfYKK3PIzZvCwKaysQo8
Ha3Nn8ny5WP0tsUMFQrXXVwHs0KKJbJfBohej4+AbgwSofU5CVKY65mfA10R+9EE
q6qPbLTEQem8wjEFLXbKdLdlDFUrnB57HIlgVAHxNOF35hn8QOk55fjwlmrD6KZn
REuPWn928CwjIijHVlweLgU4GJsLtzUNLRPT0+qWcwX6YcXMoBc78UMavINReQQ8
Qn25OERDE7G9QGbREBk1emNWKXM4HjOYTzt+3QXbDNuVG4M7yE7Ay2U1Md/B/7kZ
p3I/aZJBWurezfPqNrnai7tkVYJWqaQzzi3MjwxSdXas2Pl2nNOhiNh2w/zsafxW
w5hdPLPVUGG9fep19T0zxleyNNLR6857VD3zlHvek6sf5WkFe8kPDZuAqrVCXIRg
9SLeE/asd0fyml6d8WHRWQjxxzaq5aJKomcAff6DFerhrUBdrfmkaWxSUviWzFQ4
afxmVCVAhTPiaiz5T/9xHmxqSGOXCJ0uC3U4dr4D/1C0R9lLt4oWIQrUQA9Gxcar
EKEE21kybUCLp9Q/hJnT4+9yKv6BFQdJJ4E0gbQDsDXLnAuKZSkP1fCIkJ3JELBf
560Zs27QggtO60+h7E1rN/uoPMue3/2JLJc/KjN8/M60nthxilcpWf9yegOWcfLP
8HmqbaJ+ZoUSKtB+swmNonwyF7rg4IVlHF1TCzdtV7ROS4/KJHGgWhJIBfxDYJzn
adhe/j/nzaqy33KFULEcF8XfLw2bvfmKDH8QgsX9r4fwZzcIK3y7N7mvUDGv5dJs
e72bpJaEeNpyvMON2yypdGXEBHdvA0JT08pgiJXHpUjQ1oVQOmiYJlQCtMeVr8P2
mAHFr9cnQRoT0rcGUdn2klwJcy0Pvbb9jdDqN/J0UCqb5BD5QMpHmajbUYCxiOH8
nMOVgTidAY1RMPg8qUzNfh6wP6jScT1UPEwls+w2n7q7MWJufYmpW8dOQ2nUoUre
JURScQyPqaoA5yJppENqs2FnQDjQeqz/LA/S6koj8Bxw1KbefxlR/rH+uZFU4QqG
vvElP+Gc2ZWwpyeX/ccH5LFO2QD8GrIhLHwv5unjHmn+fI+MMKXl3ylUAnEvSKHN
2F/HscfOWdGdqYQsCIQaC4vZm0/DWcnA6NTj1Iu1o2CukxUmjYo7xY7NF3dryHiL
dPv3mQ724JqCK4kTgw3UyObT7xnkTDgS6RvhsgUDJxeRDPJAhjE6if4/dtd2mh2a
hLLUyj8sa6O4TO5+XOazNX7fj4bbnE8jDFGJf8SUB9IZLh1JHaT7CLeJaDJX7IRO
kfZ0PvBvJtEW+U/5tdmY9pcktjs3xQ+2289ZYLUBZYEX2sI8M6iIRxYOmymFmIsY
EvS7paYbQYPhlnLFpHHIM+exbo/PirqmM0LefAdIpjQk01yeohTk/cto0sKyVslU
9XlpBnG4UozDNZWvV64/whVv+yaTGgms4EnT82VTmuoHSebTKF3FH7KR43a9/0Q2
7TRm58mbZbXmlnrbR1J67ho8ZH1v7WyDs21tf3VCfRpqUYizk8MVUIVXQeLUE/Hh
DZsgcwY4B99vOSMDuYRnZDF9zExIEX/Phv+sg2ldqVQtkHruXBFVQla724NPLEFw
AXrF3YJLF2BZoJvCcImNRixBbTOGyc3eUX/zK84UR2vTDGcPKIXv3fA3pKVyy+iI
89+NYRUMaf5HwkYw9sYNM4ef7tbI1aQyh+AEJcLGjQJNGe9oA2Alr+xtdFKlhq2x
TGeQ+ke4WeAOBxnZTPVULkg/7WdLipoHc1EAEdJuY49LFYF2TAyhbCpW/LfRauLg
5FFkgokvvyAh71n502zT22igzezikP2PCyyhK7nJeOSE+md3lVwPT3XAurCIud/Z
INCP+n3iDrFBz++8fbwqktoH4Xw1p8Qk3Z2eduavW50tgLx7vcHf7o+5Qzz8/TNr
/vVk5jgjU6wX4BIDYmwD+kBV3//FtN5RPxbzk6VQtVk4LmgQOzJ/f2oVlQfRzoEl
eaTYuXwrS7WEsnppM4vEoZs4pQltRAMBb28K+R688k19mClnZjN5mObX+g5C/zu1
bGTCbaKYbd8WJepniFSog5pprT8hw0hGdx9Xp9jcEn9vnVw6ztQ/X4A8BVzIb+5V
ypSKfImjjMOL6NjPj32l7vBKHgaEb8xdQ9PHoQwzbg4ruBw2lXnZzg5sJhN1cALo
CDRbBt4Rs7GrkmFNqObB3W1lPTy5LzGERa16XtcCB35GskSoW3ddI3QrSq3QsTMY
5oZer2ziJCvjAH/+UgOnZ6oscTJ+1sFjZMt7bs3lkl6IqdkgzL3xdCQo+/B8QaHf
XwNi3DM79iilaEo9k4VzSvOEMcUMlWmHPRW8h/rKy7PopTZHWooqLMg9U1fca1QC
dj9OlLcnn89Abflwn7oDxTXkhMRgrS/3EF6oJl6XxDCAIy2tMxV3jqJLXoNdAQ+R
15BK63uAcQ4kbzVowzrObI8WDIuh08W6M579ppdOidkx/cgjXvV6paMjd67bESqz
mqf4AnJTjwAA/x7bQUzsS3cjsr5DDGIEYC81775GGb8kb/VBN9SvEx9wR3Bdag5l
FSiHUhgoTUp5vw9Pbfggag0fnnT5rh+jaoUauojUfByxClGPPFUC1eMNuwzPXCNR
Lnzq1OEUk1NBI+InbpvvbHeHHO8wERRxQsIyBjyKLzlclkThBpx+8JqQXQZB5i+t
m6U0nxa13VxiH5iPb/r5N+PvOhmerwCLzKLzX8Yp3DDD3ZA+Usezrv8ikimfvcmw
jx2uRov0Hlq55hNroo36gbSzgrvh5yRSZx3FjnWrSmvbEKKJBwyhKjK/oE3ejbhk
Mqc9ZHJeoDn8yf4Q0y0lnVcRvpHMHk3qL9nNljjsFjdalqzx+UqhqhVTuuetykBU
x5S9JfdCZpmOhQ6hhWfHOZ0BnDecyWhKP9XpnJSj3z32KEFk/IAF6d8a6jjy6IYk
gSnsaM54iHQycA5JMQkPKqzkQMLAgus4fZEzuSJQxPCHwqzl3KXgXKd6+9Eh9pQn
ILpJ8L1LrhmlhnBEB8ZZHlhTR684x4NBQYBBQMQorMhO/LZQSsSWvYwHTSMXDXRm
MOgZQCm6DPat2yjbz2q798kcoStVd1PhFSLFcxIzAuihxA5gkpPh5IR3SZAvQAQu
nP7c3wdjqOhb+dgINeROhUc9PSF21YjMy/tzqAQmhig+GJAlx/neXcS/709lNJYi
SglNGjXu0CmrCOCiswpj6Dpp3836SPcaq0s7bMuESxDQLq4zz5Y3I1UGaTh14g1e
fDysdBZXWnbHPZygoJK+Aq1Kpn0Ll1yAQQmFPYoqldfe80JwgrjQewAUDADvFqL6
M/MJ9DcyVomDxoKAWUOViHPUHLgp5BK+9a3FI1GtkSGKVHKNqxhLeVvK1z/kXBEL
umr2/ga4u3TiWmp5Jjl7WdARYm7VTSIEO3DBC0Cr+CTVk5yLl89q2+ZCiW2hqLNj
kXj2shpayWM9RM4EotSAcfSKzF3xN1s1l8FWy/wCEZFZ4VNqrF9WVOitTrrIVYuP
1cP6oENsV3FZplyY7DU8yj+kSPKmy2vottom8iI76wQxi5mQeed4kOE42aGy2RGb
TCmsZxq5LNivakmWzNq3htxnx4dSoo7iV26IAvrRbgozX1HMI0dBirsxjUaDWbyn
Ac5f2qE3omLh6tUqt0+V7Y6fsn/bBbEmTVkOfMbAo1Ivoz6tcMe3sSRo18cgnHlL
gvveIk2Nn1AhQHBRgM6AJwrJj5b/SJ2FFI7aLFSRbWgoTMhkw3i1rWhSmH3uxj0o
Bv3+Nn9bXqNqYAxJ292Qjw76aJkgcREBjS4enLdklW3HqL3lMXLAtqbdGzthbPVU
fQHtXwk9q6/dnmo+Pg1YKiyPFMuZTvNGmNKYjgoWgy05Jz4PYcLY8bzuvK372YAD
fI0fDyGjMGtBOZWSKwRaifw5g0dio6vpPDoGxa+uaM9wTtIedPJAcCZPF6rsjCiu
GVCPteb3801KZEtJxhQv+lbrsY0a+SMQqtztkZkPrtf6jmBkNl7KLPxapuECcu0i
bwu2nd54frwhX3AaJwnYiJa7HUElnx31qOrVnEVFGvtHaBe6iaw61TqPem3DU+o3
LlLZaaXcgH/QWCH4b4D9cSxsTM0X34fZN58vlxT6PZHvmCML1qyDJmZSukXyodn2
iHc+1tuq4gEErfpFXpvvXrm6j3ChVFWZbzAhFlA+RTMu51yxHPDEXi6gqi+CUrQD
+PBpy+KAhBdxKDl85BIEWP/nIjFS6Abj24FyhK95pUgs7xipmhpmnfLyfB45w9w8
s5p70qVdBbFmpvv4Y489X2Ajgitw09qHwxszEF16plbP/XaYAXgAWLThBS+TRxPO
UBt6zBGuTpRAoQMrF2JiwtDUfscpvFx7q1SCMmkGVahjiRTR+5O/TZbnpst6F89n
8QAvZVxGFwVtb4Ryxbjifv2WS/5t0yecICTDsTXovOOV961ptq/hTeZnCCeyJvew
zuOB5VscCMd/b3c440IOrUxkr28GOLnXPiO+xV15S2P865C+DBy+Gw5kpP3VdTNk
pir8P/mCqg/3CJ6H9OIL99lS95Z9nbts52l53o142EiYcTuKoBNM+qZGJFeghCBV
1bhJAiCO8tQaKdqDK+djHwYLMsOffiQRe813OUvpZxW9TDhCPAnzOCJhF2V6RzFm
DJQ1FuwoQbhdqKzyFuBZXP7PP2s/xGYfK6G9K9Iobe9tLCnY68pKucVE0Dx0Njae
mvXc46o7FHKeDuWeQwUfjT4jCSgLpcYZCCWAHm1QciT0xSuxYvbLRHPAvDjOSYj+
z5H0Vaf1Jj2ntZ48727n+r5kHm1yf/TvsBVBX/jVb1WLtB4qrv/tQ0THZYpIGi43
CQkCq9QhPecBMzE5Hrzro/CzADhULplCbEr8UNNCnjD60tHh3T0OPrzKHkfktzMR
P6kqnH/H3HxmHsw5JGN6dlvL25uPY6U6D5oagEPjUVPL74KHWe4aim+foR2A0Vz+
cx7+8mpx3b7BvUFxQfknE50oAYh75NJx87VNBM20k+vmaYlfJ7pCMIqZq40lAZbY
yv5ow6khX2OcFz3OjIAAaolJxbfSMZnXkSE4nDNuE4+B8/YxuDSYwWSZyV1jO4qI
J0NXruQzCwgw9Tw/nYmoM9JUO3Gbeq2SvRAlRO/TaWFFTG5IzO+8Jg9J6XEd91lp
evhD/ZJS/DdCQR46UdUSxT3th52jJ4WxOi9QaHZ5seVC5cSaV6+zbXUFPwGuo5Zd
Og/aM5VGVuTTqgJiBpBJdMurMKJNLrZC78vPOONxk7+Y6UQq6qxTwqf5UF4YLpLg
VN0tkCACp0zxL1x2qHhI7L86NXbOwtEZIoaEnnvA8hzNnj9v2MLWPUB+MFVw2rEe
EKbHSDYjRKjpnJo6R/p1JB+Hbz1MvyIVBzaVP44hf3vdg0J0ds3plGz5ahTR5b8V
QmqacUPmigb5nrq6N9vuGhp1xpLgWZavPKtUp3jNHlQ7wJuWWK9zRMI8sev2QTdC
ev/yc+xnvxGjSscW+3FDzFsozjWW1DL/0bGxXy88SVE4FBo/yaebmYP0EhploZ58
QfoHaxBHDlHwxKSBdoT+D+IYCWwFTgyHjncU2WidLHeIKxISf5Y24QK1NSc7cFTM
znGHbImnS58FNwRTl55oDRmdZr/CnwZwxCIfRxRnY1LxKk1uREhqt+DYb2TEep4v
rGk5xWGe0091SHi0H8vOewgw0AqHpwUELopBAcSDD2CN9BnajEnsi9Sv0/esOQL6
H/9bbEOxmx+ArkfNbwtHh0/9dl+iXTb0kOZpdOaPdU0xs9BXizIRz0DRnwgMvT83
fZox0qa7BsSdAvhOtM1dUCBjKCshc4jTSaEZIgkAI3JKMoluGTfOmeoj96AbBoyX
snOaxOI1DCucnSeMOyJ4MJdaJEnouQJ/odi0ykvtqCgu0gNUhB+3u7aUJ9F89weR
AzLQ3hiGrA+Y8Rsmb34xVpR9cZleEogpFTy4EkOIH3n/SJFd91AjFhawqBLx/2k/
mgm/LqhzciKMDejIQuP2P2Cs+E5sEbxzMQ0+3G2TywShBtf5d66xlyg45+4i3+9Z
G5Df6+NqpbGBADGnSEI5KRuwk+S8qNCMid8svPk6+RcuHf18+dNZX6hgxcJYao0h
xSBpCkQjMSMz2lmFJPqf2dPwsgDaroYSwzZXUXp38Z0z9SJz9KUJDOQvcxx+nmyV
YQ7Lc1BxJ6twM199nQh3Xs+VJJ6ngdHCJz83JFfg2yBWgyztCJQq5vUkUi2egtCO
0BtRv/LuCao2jUGrsnIHlHfJTWrLnPpXOKmLpjFNYIslfGwflLReIECiDWp3Z5N8
Cxuf75v4Z4tJMOLX5RRIFXgTKCLLcLo0GqXBnT14+8CAaaUJTM9Ou2MvFTq9RVq5
Is9Q032DxjwBu85zu7+qKzkaM4mw2auD8PxeplKvP05V7UPR+5cXdVmqWrxSDhMV
1fQn60vZwNJJrToOQ1gpmgJse0WDRBCDfywxNgMgZs6c0qLXBUty0K9b+Kdf7FgR
W0Lq8GlvF2AtrcuGMEIZF+a7oUWv/NJv+vtz46Mpvl7LhZfEz1hrZrP2YhDysBHA
3kUmkobiZPBq+SeT7VHKAJGSExC+fdUyWkVJt0WLJj5YQhY3vHbjchma1vOrN6dF
Uh8JEsfaG5UCHIhpD1YZw+GGbhXgk1i+GgyAgK5TEjazezrXvABgdjUn9O2jVp1Y
mzPNCJv2zdOCy4Qq/6COuAF0mUvQztI/F5XQETn0K4srrUbApsdIEPeMWnEB9G08
CgB+U2rqcxDGulRDsm8MhY+4BmSeUZuYxhLUVYOMdj2ljgzoHCvz9sV3OpEW5TQP
yeBSRlxV+odl293xyBenzm44CBq4Qn+f9Vnxlt+9YcwvBHrX9h/kMqMBqGXCUjfo
I/aQnXR4KuyZRV9qzVLFmJozLVbaHd8pLD7V4JlBpoRZg4zYOwhhFqi4s1uvNc10
h9rj72BuRPxuJ+PP/4iWiKocaYrKkmKaZln3A4EspSYwFxVJN6NLGfnIxJlrToRv
xDJfc5PxnDGegGLN81nShLzp+eQddVPahUPwDacAaJyel8pAI7lnVzUfDkqT0Bq/
ohzbheTzgM8NK4s99/rLNvTqzLM7Yz/C6CrNmvBU4IohxdYOJyFgg1eEECmL6S3l
QoXNovNnHbOD14KYVvzhOJTbL1UNiClZKWuwRi/QmVVjnbWw6ODqkSyPGAmskPSH
4IyV8e99hsj8MKiu2yGGlyT+k6jo0XJzPZft16A9x482aoPluloTZCE0SXGGDLQZ
KtTLtY1URQ9ZxK1YFxCHZnNjC/FI6v1sULZcQaM3SfypylGCejOBD88ybdTVVTCR
Ut2CvVsDeWorkYxZCq3QpbzqgUOXn3nftiwMXEXBJi1k6scekgxYCT3WFmaBHFGw
pIACp0tm94tpD12lMA0+XPehxHmgojPPTtWSD3sdfuXA8HPZCT3TrU0KhLgjoiKD
S2weqAVIoAR0D0oGfsP/Ckmc4A6+cifKnpnGajCP0GuEK4KvPgWgkNuX/yNgzmDL
mjHkPWDbXDAV55p9UfD34koQFk+qEL6n+SsFyzOIuuKGwuIhtdjtZoFtrcAVxB6F
XaACDzPjgBRGC34bf9QIEnPBpQjIR+u2SSUyl84b0Ii0o3UCFI3Dg8eHbGCj/1y4
WE31aCbzdhtGmX6H1O+WzHbdJQq4XSYaimLYNA1BXvUffcDg3lreokXpMs75muGW
7vuIxnn4MdgpBcbZPCgorurRQDMseQRm96S7yhRMJtlawpkRIokevNXuA3hTt1n1
77dyKW7VcOpWt8+Hlvh7rZKdWO8Vpfsd2MzpB5l5DhGVKjAp1A2eOcnM7C63rBMW
arNosdHMhSfGvzM0OTAnFk5nvGVTQOQYMjwReHSOvVZfhbSBvp2dYhyD5sIJmAGo
05IYRdph18UkH3MuPSxdMrk678IgOobkwlsbRsSDbAtxGdbaAFl2jyxyXvfMDz1P
JW1sw0G3ddyqXRYyLBlVlB/x8H2xa0SyI19PJfjJGe6PvCDypGqr14iyhf9bvjTI
V5j/Yqe2ngFp7gdhRf71qKoNtyap5EcpT33e7OIVjcw5FIuQSEAKRjz3iaRjrbN8
oekXdxS3fGtaHsywmNJZ+IX+EMeRwH1BP8YseuS3+Epv9NF4PVT8QehzI4l5/cnR
LLdG5UNr1/4Z+8aeNYFsqGGY4/Y54PEmyD/LsXv5Wc6QWS/eaVtO3igEokvKJZdK
C0PZA0hHooqkfkjit2W2wfQyea/Qv8whp+MJccO1sQD/roXT3WlLSHhzhm35Al60
JKxHLjOxFbdFHfUcGxF6gZYqRF/em8teO/Aex0nU7xwGMEf20N2gQ7t/Hqd+jvgk
/6HqoQwAb0a9qr2m8dfahAnVybBxtHiXtfRgH2SSJkrCrGGK8z/Bsx9mpUnLWGCf
/bbBIAmFV00bSO7d8c0WG/5Pw3gX8V68mZ5E+PbnEqzcyE6pxv87WFUzfGi9EpwX
DE2PEZcItxwgEEMw0CcQeniAXwwE7rIK8Ur6R+VenHpfJ9YGytYl+jE1AtEARLXh
MeturP/19N7CTwAPVvxWohd4hyT4Jw3MNGIqZG5f+WSqj/lCP7N28RwPtVsqZItA
1+bYT+cGtdUwO9/saj/jw8DCnHFvvw/2INxZfR1LVkbNr7CB778hkpZ2p2U+8uBz
7xgK4svGTwx44zNTgfyo4axDdKqwpEoDysPnsdvWOM5nmhN0MpG141kgErUM1W6W
3iZvWBBQ50gIJfVuUaEjxJsGGXyhmxQ1znIsDgOnu+kePoTsDnMGiAi/IhcaGa3L
1Y5zU4kNSLEJfGKBkldDTX9D7/AmuU8zx3+1htZiUFgKsdPCwJgtXOECwhAz4clp
xTYFxS3rU55Qtx8X/ULg5vTlJzyfsrwQg7gkhTEPrv5aPy0+85hTynYuK9dCq0U4
HyOFuiEVzkZfANXdfKtERgbw4kEW4eQW5cKZc5LGM6EHpghT1JeK/CpDy9oJ1lyZ
WwymZRNL9WJ2p/zFxq0oT4JIDg3GNeYy8vHwTirt7niNEtQB1RtIMf4zgp4WP2E2
X+v7/M5M4+E6mO64vEPHoZPvy74QGwgp/Pu7dYfASvYCMMHKMp0FqSagcLPmIcGx
XTbC80iPnNoC8C4yxvy7tBMFStjzD8h+BtY2/4u1eciwrEkbgAOMVwGk5iUxVm8K
DuV1v2rlVIUiTealkeLHiQK0KRVdg0V/2OmPO83fNMoPLFkHV7wkq5kpy7Ibt517
BXpIHYRJ8raL1c2pL8PIQmgOiN0wlwFDaTJQlGY1FsS1Ki6VO+IsYXCBFtRTG+4W
wa5bkr5dHvIxz0sgLAwYPee3J/SsLPezG0etxDtcXvDz2wQwyibDdtMK4Nd8abmh
oQssTlTxXgu3BYd00wwmm0loW+gAdTYyIBKlQEr5S65fVD0e1lgqiFQQ5r5//S6+
TyRvLc9XUz5ycJmMbcibLsBGSVlev6/DU0JHwN1wjc9HW84v+vSBKYcvqDbdFOgk
yH6o6IBIL0Y9veQs4q1SjlO6oDAlsgnWa7UfpbNd+vDotaRvlLcbWZA0qJnZw5SJ
HKhv/YZ56pfN9mM6p+/yJKqvhaAPB9ynzpJgzsMoIJ4WTEwVrI77tLsx5KpiLLF1
XUarza3K31BnfWih38eDLU4FgBGnXyVKLrolTYhyHjnpJAHnsigVReqcMKBP1LxN
t/y0TrJd4zc4HXd8cW2CmQEgOW2+7T+CXRfjMLexqG2FAO553m0wdREd7ZwTkYTF
qT5QZIXqdSi2Z5YLkQ4aa6ncz8HdrL3ZQyRmmycU3FpHfCvpOGoyHXBKc6oudDGC
x7qsMOjx9P+dnGVrPuUltWoouuhVF4GlyfoCf7auv0uEzLjJnSfS8eqjHqIINuHA
J3wcOCHRGAK5qjDImBBMw+CeWD9k/+b1/ppMrQaXnlh9rB8eDHcopwSh59PQPnn/
1hI+6rZT49zKiSbT22l9c7Ttg0tQYblIXRj4Wv/fvxlJRTmi3MwJAgNNIllZgDnk
8tH1d2d2qnc/yPqJiMDSMpq8xkWNzki/rJPaMhPcUcR+OEbTsSGUBoMtrfmKiK4N
uIyq3pdz0NQ/XvX8CfJ03TRC9gogBfNKGgDcJMIMuP4owUZksoVmnkz7bQbHFZiR
eFyyy6z3zRfbKyPB5NUVvnJlNTo6aZtdgixQssRkllDALt7kSnJ6wAYYQFsfRIbZ
hyRwA1RQkCIjptdOFxeNl/+ojrMsGTADhC9OU7lHJRlyT20qW/zCJJFXRk84cn9+
w0PoeR541ueyJAdQJnCkVe22+iA2yYA/BKR60U4ou2t6V0zfToOPO2ylvbku/Gj0
xW5afu6H3V3QAVZyHQr8sm/sFVVLYzsXRZML5d/tShDzZfVsNwUGlMM80izYKioM
iGs0Wh62UleC7mQ7hfptBtvq7xpsWYypZDMod+2L4YKDeH5a5tbn2z+bdSqwJUuj
hmvMR6nLJhoAGuP9E28jGoPWfTJJWsoj03IlsoWyLcU0DymV3W7bu2UPU9oxD2Ut
xI+/Yv8tXbnjuNKSA2w4Ijr5jjSmVPgNKmlbXoCFGs3wcHskUXkDP36cBPiD9VMp
CMIhTr0AP3lZKAheJOBT1WjSppp1fle3P3QSDWCeBQ+urgUn61IGQa8poxVEc5RR
0NNVdtm2P31+mvoL361/xW0PKRu0PfmGdMuNEnOXLOX4BZQnTqK9XVrOQYbnGaS8
QeF8sONIXoxzJWskIxMTBm7f2hbz5Hm3RZU+DHYc9eOUhfar2flpxg3cB7enjAt+
YCwziVYlwYQP/oR/WMhtENGteaCOR+xOfdQKH37XxMUY3heYm9mGNIf4FNiUOfkA
tg2HG/zDZHO3uZysnT7TUBepSytmf0l24rhC8FLbs4sGDUW6LIWstHAg1ukxuoym
UUAGsoOx9yLDbShmx2C9RUWWVm1dlGBOXxcuE13L/VVMe2NbXJap/2jKE4gtKUER
eufE6xyCiQFtqTfnGmeHtcOYvbKyza4r/1k6w9gOlAIoecWqwp+T7e76NRWCRhtE
+u8hvDP2vYlmnmrxdDYl7RphsHACh9gL49eReUhDvRXWtdkpytvMDpabOyw61mLw
mO+1kuEuINyVUPQn6fjzoZSs2PrqsxHUV3gg5fSPGxTtj6+4vMGXyLCQiegk1Vvr
+im8mVlaMZ9JlRDeVtMHNuBEz2o19f5FD4u1P239VQu6iHN/dXQvfT6sZxSCfY9Z
ERAZfHItthU0jKdGHbj+W9pho51S2OWjmmRpVLvO+40gKxUDZaxkmUob1/QP9hLa
vOCbTGux3fosDvddrLhL0TAqVc5gRRGxYlZBItj/5QOgRw9fmJ2pqHAu/BOJjw5p
d66Ah45rw9aJwrbtzjnElz4HRqYITJmzEskCVW9dcNuZduvVsVsNbNLiKAYkQlxR
zhUfU+OwzFoDjLnxfE1jMy35lqL1KwO4sNCH9k/PkvBpPIhLtXAW/QOF7f6BXFX0
aF7BUxZXpNyYvHu1l6S2PYiQfSqMW43BtvKasLEedsM0IJMI5/qdRVSojt74rDl9
dlzPiEF0fmKhYPvuOgKKxikKS+B0OHEn0/yGJIGM3KSPgGYf/4RPJnM86qmoX7kZ
vxg3qo+uJjhzIFR9q0GCZMq/J50OJN+gh+IrMa+DV0fqLCNOe5Cjws1Da0Z9KuCY
hcPRbTW23gJyktg3Mnhd4DuUgEx43Z4jTvlBXRVKZycxAsR4dznLXzAmv98n/nWH
+MBRM1+kD64gUTLNbcD/Cwtf+RuoPnf4rJr3ExNGaZtkK897vd93lWVL+tsiXt2z
ug3ZqAPKsZNftOFvHQsK4yv8YV2y2kw210tCH/oZLNDnGMlZboQKaTqPFLu3xDxn
Yaf2tkP9DfsEt5gxW2UboEjE0zbDsBZU/4213jXFIM7lvXwR6S1aiIhcM11IRrEl
oWCmvTOfPudVJYQ2ZJInM0a+Po/Z6hYL9HB269R+kefG/aWBVZ8wTzcp4HrR8Glv
JJwYdpQ9tsqwIAilTC0S5rCNFT0cYKRAec805phWq1INmLH7QAvhKeulO8NjulCz
G8jzePuvQFPcPCbFaxR0XImfEhaLoTaHw5F724xkoQqSkP4JmfjMQIHoDMlk8MC5
X7wSxjpiI20kBteUYoqNmwb4x8uARtqqLRf+Cp8NAXQFIeUNK87PvAkEpW5LnNId
qEo20xtfeHslvko3TaPzRlGqi8DdF2JMvUO+LyVA96ctlAZddiaGT9UouMPvIC8X
OLLi+eAmQ26slmkZXP7RiM3fdjcDzJhb3vavL0yTOKn4iM/MJQklQX1RJvOKfssI
1c3Eqxys9XllYELzbC1AZGKnTgI4a2SuHYdeze3efhlx/s3iIRYX7xnbdbe7IUDY
1026Sv64QmNe+N3PNeZltgd29X3PoPt1lCjbMIvCm51JigzTHBIPovc2QEvNQUDo
BYCgzXqU6IrCQ9SNSVe03CvuM7Ynx4bO16S6O4DoJQZcn+R3i+4le99G3BZDlhsw
zE7M8qPmG+f05RISkYbxZb5kZfPE0PSM1WSdNd9Zzb2mkYlwjI/4yGFQLk589taS
0c8LTvkbMZxWK0RUuzD+KopCOIh0EYH/8L1pJ2RTDgZ1O0lFixiMbNfjVIYj/l1+
kEKtvkN7UDXOAvYXvI6ouvMYDiVk7l6C9gcD5YazSiidi4vG5h9gt5Skd6lPRbbs
8TT0bCyM0e3kknm4mGG7cp8WGf6QkCzc5UTJYuZC4IIR0EWQQw4waaFZ72xAcXpJ
WfhvAZw1gFkUJHp8+8N+86i8tti62QHNVcFfVKmJX43kY04kgKS6YKT9YrfM6ZZ4
MKSi9S84MTNdkl1t3PV5AZxR8qlpgTzSSKFirxuopQikEXrekxL1tJQ7PO2sSxJa
8zn3TNby3kv7JuvAlN/yTgK2hfvU+vd0Bl+HEzSKFciFq44VhEMHDZl9Kqv2Pgv7
V6e9YKktpvgyDvZVK60qch9JUN9csbBK6HvszamsWCbjrmoXBsQNuQ13OZgHOKXK
9f1Lm85+2P+gmMbGnav3rIpTfm5DfByiBeH2yn76uQ3GzeQiCvIyMNPXpEbXW1Fo
ZZDwmfnH25VYcUulRW4liiKYJbl/RaGXRxILKjTuBY/KOBgvfw3uhm5vVWjiWYjH
+QQ6+zsLLjpFSMxz/frq2xyn6cXA/2QfzpO+STPUD5DYoDMS61zu/2DWyyNeB5LI
GnOmcgwiOzU43HgF52JY0EtwOtc9Sks/ZsSo/ykC2CWAuB7tVEZj8JYyAjztOxGr
enb/84lzRh0e2fpMwfVWtiMtSlmfjiz4fr3SU/KAL2AMKrpbtabwFWeJ+ozi+9zZ
nt8Ghnrc46gtKaWnHuzNgfyIPuPtD9EO119hPNfnybRstpQB0wGlck1OI1XCMCMi
9mW6rEirBfqxNMA6tf0UldGZjsxo3MVO0sQejFFCu4c+JxwHFWMih9z6rZU6iEp3
+wH+3AA7t0z7KOMQRzckUo//RLgYKRm4TlDD8Fhdy2Q/gq70mAn9LkA+LhafIcpj
AgDRMWnE51oI6Y2GqyLQoEhenaSDjTzxZcW5FNz22FI/cJHkYwm5SySnAAT6bJ9P
KYXWw/PZcf97lz0KdAyyhy0Op8a2pN8nnXTsiuxxwWTBy8Vx6idTrVeh0Gp8reK3
4wTBv7MJ5ED/GHiImI1lkGtkp9S513aieZ73aoBd7qcqLYrg3jS0kBTn4miK0VN9
YrrMISySahdwkHZgSYEz1awCX5is/huSEcqV2pnTiZgmyALsdrednzAcVJh/hmWj
S0E2g7x/ZOshlDe983Cq1DU+hPSluchlGw6zpGc/A4k11GCSktz7SNxdfPz642Ox
vh7Qk26fL8g54zHh2ZwEX/yyumW3AEXUAYu8o+rFh/cgbFQVlGrowIYE+9jvnMvN
AlGdzenSyOpx8wI6WD9z6b2aGrhtP/q9HEnZrT68zscP8iDmIlGyEbpCQZmSS2y2
qXPWaO5PyR5D/W0du4lRUe8kxL008vm7ai4M0ZwEqmzPkCjASLOhWXgwkr4sU6pl
4Fj9S5xgcIUTCqKL3s7BZDlujCb+nLEhhmzNAvYlvd+NH3LxUy+h0HLSBmYJyW9l
XKAibJur8L5e5BNUjy0gqULAQcQgca5RcmE/hBN0gQipoBlfG4QQseQGXuPxr9vK
zT0R/3QbhxRA5sSDgIr3eLYVW6Tm/jE1hbMqIJTX4Nl10ja36ZP/x1DlYf9v/vBt
zJNiDSnLv9ZW7ZGvOden1vJWR1/5Lyx1D8kBlS4sPpdDGVWgjmWvc9gvMuXv3nxY
KYNG9TIPr5gaAgMN/OKtHCTMRpqnwAzmyT/U19bjpIzFGkzcu+pLQDhlY5dK215k
OKPqSH9DDx9cltYyYOkp3Rdp41qNfMEjE2dqkRDYPJGFpNLYv/gy3g0zm+Iw4JDg
nN9pWCMv4E8US/qzx37yKPJD6OQZ0iQKTYDDp9q8uiNUY38lMxdcMgMehrMZYDdc
ZaEPz0xKGyl7SYmgqT5JxlzOE0UWpl+8IxosqhOHv/kf/U07Yf0s+2DMF3K41kPh
5iuUrpwaTCn6XXy/j6J8zek+Y2liWeeC6u8Ugl4DdzpbBT7BBCETcxH/sAa/pONI
pQNx/SBlIPU03iPa1y5ew21tgZHq9k4T/bhJ1pKWZlr3DJ1aEQJHTwdhMo/ox4v+
jSpn7rzrYRgaQ6tEViVwSB6TuafE2k6WKq4GhTceX3vTqs0o12o8Azq5r06jtowT
kA6t+kZj57QOUVewEY/KQPK51tY/RR+m0bHGisL+fQX5nTcE4iTAbM6g6sRWDJOI
+soKZmAGJRzCw2y6d4Uix9VSHSyo2iNzTJf8qVd+d3QXL5/XzgRFVDrZHBAiEB7r
SDe7yW4nKdPZDEV71czkbYuSN21uQpvpUL5+8qvauZEgFK9y/SwSqh6LNaafKI7A
BA2fZqygMBC8UEvCnviKTfljb1OYJT4XJ/pdI/CMOMjeVr3SMtdtVlkha3deg/tb
f2lxRhvNEos9Ov/7slU6YufrjxeJW550paE9lKKYikoJAUK59NP7JPgkmP7DnDmy
LIlXZCSQ8O9Zf65eJaFVfu1+xnJsg48AB9fTY56dqlwCA6jXZ4/CF9oNLo3oe+Gp
8sflxfcGvFw9+jWUfo9RLbBxbOuuS6VsOmkVsehFX8c+wuY3bjWaWQsftIc0+PCp
uDtsaWfHA0Hz8OWCDlZh6jD3EvB8dypKnBBWhUscpw/DPlB3HkIQHMlurrB2eoau
VF1fs9a7xed5sezBzyFYkhOuGclO9Px1D9ouUo5yCLzyZL9XVzLAw9evHKUqmkg/
o9Me1kbuavCtvzV2kUMQDgncobu0bDEMb+cTzjwdj++SbvdnacC0xDAs1FwaZMDM
69nfzuNH5H0IO7H4AcU+mvZczey/AGc61o4FiYe8wMMm3q8EDNtz9f32mAnZrWYc
1Cfs0/2BSg7ZekIhv+Zy3DtXLploc6q8UNF6Ns52ghsw8o95oDx5DrO+mxln/w7y
1K9ONTvAid1GfNplxDumef3/wQiaFQhS3fWVT5/wxBKhxeLcFDisYMcwyVPWvrGm
ahqx4bA1mViVOpQZHpmMqWR4luQfDVPrG20MGjolC/ZLtd3/WBTYYBD/vKfbg2Ip
0wKVYu7Q6UFyNbAuFViMdK/G5T4+mep7SzsflD3T47Olj3E9tx2163z+IlFj28rx
SRFhKjAsYE9idbE8Xwg0NdP8FsCEKAlo1eYvaC0mkULOiEOYZQSe1WhHtycNMxSq
dvYtWRJcYRLahIa3u49EuALzSM0hIaxk79RWdv6EvNaC/zR5N6PPCA0wqqKNBPXy
jtsq4PHj7UwJZwGKgVKXjT5utZRhRCIylPEbuPHJIv1Z7Lp0kVdp/HM1Kg88t8QG
IkXPVp1tOD+7jalNIdoc1aF9oPCKD5dNYf7q7o+TVYwzGs98MP7UcQ8M/UGRQEPd
oWo/bAYIq+VMUwBwuemCY+FLdvK/fovutAGeZjJFRH+JOQhBkOh+/OlBHxDT0Lft
V3pIvTTdqOUI0MS20fYeom6zfoTOxOBP/zZKYc1sOh+iUVjxxKuJnn4MxkJKG0TJ
3vBgjQ89aF46R6wEkGAz4R00zBEHLi2gdKbdco2DP2IeA1wS/luGdro3Dd77rtL4
cDszbniGhNQ+rYABegDonrAcM8dx5uLwsOjnIVqGfweAg/y0sH558hKYvHsNvfvJ
O6oKopXHtia8qauv6r1QTnHPnvoH9go29YOH3GUMRo+gvmmtD5SmPO6iWYqEn63V
r8OOlG5xblXlZYHiR0rEOSPFJBqORmhUI9Rahe0jFEEUCdbx2zO749DRSqtyEHCj
BT7uX8ObOzP4rr2WyIREb7apfSGatq3FjKUBN2d4Ziy3VK49tqQnl4Wl4fy5Oa4Y
o8GikLkGLSPLTMtBgUV1bREV2gN6RDnt5Ijl+Jj1QJBBayc1Wp9El5NENfIcAKBw
HAVSW12QprqWZyhYqY6TWrelGmt0RYaJGi0iB8hq224lYMZ2wdqBdYhZ5xXK2WTG
fvR+WixHmHYM/Rkigdh7mfkVVCiSZQM/KZDfhNBs0pC7SNDdozulvqVntzi67qKU
c4sXQMXUeKcU3kiwT1bWZAeJDeMJYGUem4kBxzmFTFN2x2RvcgHKiNhcBOuylfRx
KIuEt4T+kuysFCGRpoBIsFnBiFUtYgFvXmCpyRXQfK+2/e0SMV0+z6iMur8LRD9S
iDd5LBedLEOsMvNdFjR07UicjzQVejdz6mb3tY1pNbpwitN+zDGKUQwSsnPoxuZR
nVrvh41dOgG7TA8u0MfaY4NK9f40DM1JcF1p45/RVpmThWsy/K9Ax3Caz1rJBuqC
nVPIlYo/hE+WbXq2mjJAzVJN8pgJn5M3GF4E9YIXdq/QGYdCd5AVOoE0VMBsQZHs
Jtuz1TWzxJKLia5OtPOOBOWzLk0G3ie7ZBkkU4Fyb1f/O8Xto4h7B7Q5EOsBcO8b
fdU73Em5jl8LzpX3mttzSCw9YBBd5kJyv7Vp4bk2EdkF+k3cLdjV195U/1F1HQ6J
e3iow2PwI+xX79VpuuDuIkAsbqPONic43ibpGVZVjWul5n1lZKkYyD1Ln1yMBNmL
AxZgmAiC984aQ/UeKuywEgYHlX5rq59rdJwG328SA72U3bMwqhKSIyurk88Vmdyt
`pragma protect end_protected
