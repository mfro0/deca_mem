// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:51 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kwadz7arrnlwSdATEOyBTZA1WISwH22wh/Fj/aGwGZGnR7H5JiVIdR/VSjo5gCyg
mkJ06rmtYl9flWpvPQJFZ8nZ8elxMpWHntzeH0s6w034vQgG+sbz0fG1eXgOUG8u
KDycwMDEYML/26USfvP60HHzdAe2iGuv/rjJqr8kiek=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21088)
2imMTkx5jVqqb/Egvfo1qf4CD/XtufAvtwaGEU5+yMhQ0Npg1qjZ175FFRiW3Buq
8+Wk0vlkhHv717+7Y9j4s5V8tKG204Fuiew3WVVkvnN3xdkLwTE4CAXtjS2QD2u7
u8TG36CBnOrsEVqteupb6MpYEHwR4bJ0vjI04PimQNeMcWwqazDlCJCyxdL8sbuE
Xtj+Qwdb6/JeqqEicwaOljvCiYLj6Bj4q/nxBPH588qs5u10zEURzN3o0zxLEolh
lADPniO2f95a9kn6LbFxYY36U1FJIjXMB0zIfB5VFcsukG9v65nos24V47xO2nHD
cliOYq4fyU+x08dTZQRqDfvLIr9TNUUzy/3YlEape5wZzAN1rHYDxi8Aivw/NQl8
aHd20uo9j7QhKJKoxUjKoTnktyHp0zFOLhOU1a6C5J8ADRCQVNUix7qS/E+/MIBV
B7EDNEuqGlK9J9HK3v5qyDyVaYDtzPUtpkIpvsOcoqPOA7Njs2enIsP+BcJNZOi5
/J/YosbW/oe8e/rJOfEUW98HtEOCCTUxpysy1l2RRTwqun1ci4asKRb4VsTR0do/
mlVwSTSp7jo+5lLufe2rIn0zC61iP34UOoXplBFThYnTjIV6AErM5rNpsuZUgdjU
Uzhn5jHZUCUFB4gSNIEb4srv4E+B7rK40ybatd6XQhbRwBB9a46fCO7bthuYOK5e
PZxBpetdsXKhLOistyAmPULdiDbeMq8cTGqbeeRLYTMWypVe1wHGvU0/C19pQbYY
DkZbEGnTyMquymh2ZXjSrjIP1K7EQSw9uezZCF9T3WSH+jcF+pF3ka3WlK41Me8L
+Ws7dDAvx132SlSJqhqgJhPG0KAEF2Z2EwcnmzD3Fffcps7Xxvo6+GSCXYCAWSdA
0tXlviDBdN7scohYVIjsa/i5TWaEyzAK1ocH37vR8sE0c7fYxG5CnW3MAEtWnFOd
zizwgrnvp+4jccdfvrYS76slP3JVETxW0oFI+v6lggUyHQc06mrytki2aQ34+qfq
9j44kOztasg+VgU3MJbP2mZuT5yhmpHyPyRvfw7YZAaj+aebcdXZDKFxI8zX92u9
CaHonF09zzzxIsbbaI5LVTJoo0+mWAyGf+xdUq3lqZcd6UouYLXbRwR+B9jRXY9o
eHSyv7pVh0QvC04XUcEM0dN96ykMGp7rIn3Ihew0ItRPrib3mYlWGeHfrPLkITL3
wfsHoDq/8mK7B58lWL0WOHsuHzn0OW4lpdzwtHSCg0sTFc1lq8iA9ZER4wBfva4p
rbtAc33uZugbxffV/cJMVKQFsu3kz1Xd1jgotmWRbirIAXouoF7oSlJYRWVP7b+A
x4fNgia/X2oOUp32PpfBpR+Anv5B1HecrtgXn2C6oLIqgYWBSpN/WECx1ic/hU3a
BFvBJh/XMghM5rnQEpXu/QJ9KPyLk+2S6x30EqNUpffgpjAT2AyZuHZrQ5y34OaF
CEVTHKDBs7iBCMFAqQVX8/2DY1Bt+TZoh40Pl8m1+JOmvES9eGTtTPc4xAnILZH7
GTJoqP5iYCu23QZE7pDgecXPRiU6ko0wNpBStH6SirZAANwyokXNBYg8ll3wvH1z
dgZhwnceIx3cP7M/fZ7PAQylSPp7Of1YcUaz3mflTIIozljMEVpWo2J9gFOFpOF4
Me/Dx9tftNPZHThMMyIfXzkkt2jWVPK369QUATmsNe6mz2BLCjZg5DausNsMOM8P
cbAQjpvnREIb9483L+AD12jT3q/I/D855/3ZU7/TzodTfdsD8LJuiAPETG2VNT7z
NpQFmv14qLUb4wxcPtQuWWavFTh8UdlZsK625w4WcWBDbIExVDJOBclQQHRezLWa
Z65w2GufXCc8n5lXx0XfX7R5SUOHsqqlD7l8djpSZUh8Z/rNT8ksIv9iO2n1G6pQ
YD9Z5MmfMoKH3nPAj5eJededO6L3a2jDPMrLs5GRH1HoQgE7ieQJHwjTe28vQW34
g5nbqXcRSS4Hiurd6s2GODOHe6VbI/Hp0NySfRpyozQ5cPaBRGbyB9dgYat9VBcH
XYAhkBjWs0CZSQlsUmIl7AuGLKAK2ufeUIaWE5pXc9RsIs/bVoFLXFh6wGpO14NU
BO/A34V3cFUQt7bqOC6YvlHFcv27ilXGsB+JeNduR9OX8hHTwe6dd92/7OnJ/fz9
7RUrOE6BnertKkK+lMf3Mw1Uzaed553OYAPYCifF+RtJZnEArzJ5jTPI3Kh7FTne
DtFDg308cFOGlYMerzSYNY2kv8Ewp10lIp3vkSEqJPa02poRDjxgzxO2ABQFk19e
9nUY22aC07LeVVxEt+ayF4q1wDiS/J8YtgXHN9ihafyd7HsNWvWw52q2UTh79JCA
bLg/0r998dO9NV6M9BaSq/Jj0s1cMihGby1b3CZOXiu+5kST8HODTkp5DmlnqtD8
2jKpzG+oERp1zw5mCUFZ9ItKVNA6cHclxgt+RbyarCIfHDPB9VCGVDlpiihNHdHV
6rF6ugIG43kuzngvpjJOYh9dT8igUrmLp8NRZvfrYYUapgFo6n/xf1XFsvSqv/uJ
mA0ovibH7lk9Tt9wD2V+0fiwwzlpWafESoce8KjAjlXme+P43Gb7xmZ4rwVAUciQ
/qZRtv8wEXyJ2sPf5sFdvGdILylH6zQuYYbLidvTMWHvOeEW0NmNISyj2+uaLQMx
HIc5Q17nr8Tw+5yB2Md1CDChl9K/yXW59q3oywlKepq/Ktuper3zxDLVktQP3ra0
Lh6ynmADQ64o88mZZV7lUipd3Ij2d6x05+zsZ0xzvIw9PrN8wjC18kf0SfwvOZoG
xxL2A5LmZwmoJ73PFCjPJHcV8Ry5IVFacf1hg8eYuZGqtcZRWLl5GH05r/BhYOHu
+XjSV2M3+rcpt1XmM9imeO5vBR+/Om6gSEcRHSE1x3QXHnen5veLXUA8OuUTALtI
q4yMitHAhZwlRQWFMhE0WGRri9iesD3AgZQ2WfbAXaFqBXS+wjgtH/ribazd89wm
QwYEsyMuqeKyolU38jITulZg7Mcfr/V046Kf6WQFPZXi0PH+BJ12JTm5ERmhbV/b
PA2sodPTDD8tHxT8ZhM+uXxXD+zTg5BioQRh0yl0mVLszIR6Vo1fI1uA8sWOCgto
SMsZe5eZONkSpYFg7gm8Mxvz8tz3QqKXFQsQ0dvFzUk7OtC4EP7FxjMWG1oFYK9C
MwQkTkTXnY6rEd2NCx5nMb+Hy8grTDYBrVKXoap5PSUjQrebnw8dzLlojGmfpcCa
Q28TqteMzFB1AlXOvlZQI+RF2NRr+bD+cyBC4l+CyqwsHEKHlnNEyK17xJwB7o0x
/cM4F6ZidKmdvizbUlruyOCwRR8aXpmq7CnAxvMdaICeEtkCUXiATwLeP2unzhxQ
sWf04lX73B5DzLs+iDt2FOtswz72TL4XE1M2HkeFmZA/3tIe5YA3Nhx4uMRSs7HY
YbqGqmhASworapquR3v3LwAzzhyx1hlXAxNNMAH3me45pDQbJMNuLdCAZQpzTH9D
MmK+oViR6GCXloME6eb81dTkyYsTGt+/8slLRCp1vQA51r5SI6F20oX/Snn9Vtpg
nPwFp+9CO97Hrdnlm58IRhmkqvQ9MFRMGQrjhh2UbOTKghObNP0TgjWCNeR7BY1j
6pyck2usf7Y1LHgm+D8yxkFa0p7gEU6UyMwsH5iwo6Ycrv44fRGy3lGFOEacRa+v
efvNDZUyKVniVIZeY76ay3ND28cS9WBEkpvHqeQz8y04g/gTEegJtFb2blqaatXg
zDUozrc9fhHwv+79pd1ePze9RA828KVKj1IZgy+Lj9AHCWwcFUNDQ/UPPKAypRzU
imgpcil2UWJg+w9Y442SFWC1PMf3kb4sq1roVVkaEzpWF6K21e12Paddhn1nE2VG
9dDwjX3usW6B59CHYOeETKLYL4xs0RYOPw9fVhA9MYEYPnPPzFLEgFRkCupG3sSq
QJgDXFMTfL7DZF54yoEmtluxwb/Tz4d1m/LH+tacWY7ShXQ2NfK8eYddsEqE0K2Q
JSVHCqvIO8AuT3Skz1Y86NmaRGyGNQneBVsGBtr1A7er83zwoy42JUiU4zZiLGVX
k5CJ4Z/CgaBku7dA6KpzVNufXHfdv7CN2YoZsG3mHlMnnlu+66YYfUBnE585gJ9d
X5idb+gJ7Bhl6pbqjnFYLFjpWkLXkAOnBn/yuEsLO5rROeRv+Qc9HJo5Fx1gftn0
DZ1Mw6Ylty2xv/ZXHiqQoGqNuudVhf/RJ4WqODxVC6E8lyxEuoBgkfghRD22C5Q2
phVu7cVRpT+kT1Dxa5SrKk/SBlDp+t0IY6JPDWiuIi581ocHl7mG5TTCD2OWeHCc
wVeMbzpE3PndaTmalW0KXg37LW+Np7TtBsx/G9xy2KvJCdRDj9SLMYKrMJVQewmb
P2QjjFpBqIlUmw1YM8ZSDnhLPi3wkhAbwuIgKofQ19Ws4ayBVr4ITMW1WhwU6gXq
yY2PY9wFFfr2Uh2yKJ7UupvKGkrQvp4qoz6akelGjFuHV/6Zt3PAmjnMClJovOem
iwo04NiYJYscRBhH7SZJ+S70FT7wQnxDXTH/sTYuvbttp7DRKHBurHdChzuXz3t/
qiTWjRdNDaWw4eAv/LmXeAU3+x28lepFWLUY/ZRfmJtE5C+4/tr0/Gqo1BQB4U9w
5rl0Fxe9BJRcditdgZhIh09TOV1JOQMey6AycenesHGVI2mRInr6MGukHF2MFMib
X62iALA+OebowtwXq9WWQzW88SClZou9y9+N9MhQvMsuiaM5xQXwk/YBhv9Exczx
wnEpiZLlR/aWZQi0l9AaEBlAtYkNU2FRu6TqInApegwfiq5PrRQbAhGEdiShp6SK
Qs2IR9Xagkre5L4UVNgSIfOpeW4gVXOqaqepoQIXf1PyBOTryr0DIUKR0ZV6r1jd
OvQHyly3Nw2dIozLMDNAqQV8FqMnjugVsrWX4JuMFv2zFIywtIcCkCcwCmBSW/j8
8TM6IpDNChalJnBkYWO8b/+M6d27O00m0zP4r9MyBoZFF7YnuWkImegraU8rVv7R
utG/+K0N6YXcg/HG8Sj8SbsbKFwm7dWn7s28hC46XQEc4jWaS+cqPj9u/RkygrFu
WjLdQX5r0EQPnCyMjrExawUgztwylX+EfKGSJBmhlvPoh1AHRMBsW5cGibHIask8
29ouQ+pu53yVUIwrYhGMd4jqeo3zB7vy29LvfpKIZPozv6hX+eHs8SQEsPBIjNRz
DqDOQABjIDlGciCO8ryHkiObFOZC/68zxmg7umUY1Np0giB7m3VKo1kCTrlB4i91
OMZR63APxopmytUhYcudWPIo+HB+nVyob+co35W1EuKYsqtbJIPhOufJPQR7mf2z
uP49G8rXaXGd7X7Paoq16SzIJnbkl8r+4vwGeE6MUcLtmvUiYf88oE1KqsR+AC7+
I1orVqN5PTBQJXh+5/xAGNUyonoJIM2PHgWoQ+sljPPUOGTwKr9mXUDblpogx6AG
uuMjnZSXhpeCPOZTcnS7YVV9EK/x3RkVVfIgePLtXvblFGwH9kIzhOlWljEbCiVt
zJ4HmsAxr3UzcTtlOrtKbGJN/6GjPTnMQXlBsvoen4KuqMX4XqsLWrDie6URGzCu
YhOobPMF+xuedjxOSIOM7i5E7dmJ5H5vhgUldDjB9qky5UJ7rGNTKWQ7gH9klz3u
ekx/yGdTpPwiyj1MoS9HZK+FgsvuswmkOVZ2VL3+AkaXNDRBgrAMAU9TruaVwGfW
DwOQVglOkpm0iDbO66wg5pBcXdsPJK+0rRmxZcaKY/vwbOLYL2qy2qEQJ6/PSZmc
7wesUWfMfxnhPKHDzDZlC8YNQ9HbylT+OdkkEMrfv4rL8MixDFwkj0KMxbrx4f8a
9EbS1A3c3jBda8mNBFoJ78S9wqqhLKCHTCWMYotN4aS/KC5Qi3Zd/X5JRrmfKZM+
Sw7IJ1CiLTIlPtalafKkXetpTsXAFfarL5JygtqZ1hYunfMCeb8uYUOFW8vvqSMv
YC7Ie33yrjOPJIcRRmLFR7RlRQPdzvEDK897W/FY+zOuF8rEOlnst1xNzExiG4kW
BI3Kr9bunAgSRZafocoiMgv34jfwnGQktnxR1lPib/j963+1QsGBI+LBz3+EP8OC
BCZUkmHCPvU/KvisaxHSWVDP82wYjW6gNibiWu5DPp/VULKc7ImWm2nUSFo0Tqjz
Gyyn44D/OTcLzVksTeAx2EmgjhhTXhNC5hkML1SUX/XtUevTLOAPNKFcYtCqJXCL
9rPqSjXrMWoFK1X/F5tdz37bEVzQ5pIZmmG4EzHujGxuqSs2nvrWS5Un+6irCLMN
P0OU3669F5KM1CMualPdU96MpxWFezoFhYh3q5xggGpIcpXChAEmHVYF60X8aoeG
bNVVySgaoAQeyFPeyi/Qm3dYNgfmE4ASeimTdN6kil8x3n1mFIHuzNh+7JXFqnFA
SUQTtytxLeHUJo1y3s0W/rMroSeWp9NNQcMM8RBUT5jSHhSQwFYtQG0Aj7+FYsKm
/QMBAfPsRNV9mqt073ZyFR36x0eAp2OhrxOUlrPbwVHB5SKRIKYmpZn6e+zrG/hK
kIGltXV3OdZlHwrEcMoWWxbzlVgEYpzUxP+FTyuj1NEvXe53DmSYnK27soel6ikH
2XU6d2QSZ+Alt12RBiQ1i6vpJTh2eQJd6bACSdpsJGzUrttOFfKp4K79Ow4qDQm/
EAYaIhAkX9x/q2KLTHt9yyQx9MaiNQaLmMVUTCMvRo2KGkEY7sJmlzmyNpW1FD+o
c1yqs9VfM3NOSHaRlxbCyhYdyM7hG3NSMJ3WMbS2S4soFPaZEzcQ+CbObF7Vb+Dp
VFJIobu3OXVpjpmujZZVzIAaHO4eikVxlQFdM4736SJbr++AqsN4W6yx94Hdit7G
rpmSFTy4mVxJfqZojmtDr01HsSPZ+b/ZMZQrngWy83rmIU1sn2or6/z13kJf3TEr
nwmJQ+QEtpIu7yWNtDj9RpPJ/1QhivIflwVnps7JLc0urqcxECvgtGFXuDPe+PDM
HqynY8vsrziOYUWzFkgBwm3IT7h9dmM49Pk7T2Jd0zQHZMasVzCi5Gg9mlwYZwYZ
VeRkR4f3FOgW5Q92cZjNdvUTLpkyajEdJnlwz2weXAQzbrsp+s0vd3DY6Adcs9wG
SF+mxs9qr/2MOIgtUjLUdcPyHwSvjBeORW/Cl/+/5/DEmLLi9JULispPM0MiMwuz
AbHPiu03cfOasBQRaItdYln3PPmz2qpep77o7zQj3u4OnuiaM8XmyDQzo44Rt9KD
eLQMtAgqSD2VFbyDoUJqLstgdLh89pbSBNdvwyjjY5i9/dj1vamfEVViEAxJDpUM
mrSciQ5ndTOpgJkm1EpGHBh/CTnqica0ed/4TKFUpFlPJ4Ptyz9d3H18Le5PBTg7
cxRIOgGXDvIV79feaOIeMelcwk6DXW5oaXzlYAdDIVLVGOCJ1FhEpTpNfPaExOCH
Fs0KzDbrhhKugFWGQEV8Pq2NoevjrGjtYylAeL+ToBV9/hX8/DZg3vF3i0yo2jBm
qkuReETsRTbfTAn9v6luFr+9j9swHPjWDtRN0gX95slqQVUx44NHF2ZzWOP9zksQ
fLtuUD2OBeJadQ2IIrotaw858ZZPFPQskebMn8yAyRRJCi0sV85vmXQq4vKD8iCc
XPN54C764YlQhJkI4m3mOWRwglcbrZu/BUGuTIV/W1g0gddrPJ0pcT11K1a60BfL
AeIfMk11PsLhLqwJ3v1btGbrSvKxqZdIIWb89sunvx7Xhc0yS//y61tLQi0x2GfR
baEEfavAc/vooOlEseoBSGBf7SeqV7MuhXj1CmP4acg/z8NLRY2fEFVVoAt8uK47
BMTvrcMWqe6JFMtB1B4kfNbYeYe2+20+jOYx1lg22Ynui0WJqXc/KBs+62CQPU3O
uPf4Px0Mvmh07yaMn+ewSZ2ABEONyVo2Q3kJVF/8hV4VGvHXHIN4i1HZm5W+rYng
yuTffF6vAd5nJ6dr6y1UB2tnYrIH4DBD5GJQFPUqfzDXk/vj7R2F0wFMIaC9Y+Vz
QBbQCk+FHW7OZIzUnvoheDT1RyPFsABxVuhxja5T2LjbRFTaxeIMxxPIi6z0EMNF
cNRjCxBlHY3lXho1tc6FqAjtnHhKKV7U1yez3kG8A2so4Z5SM/uDOtqRcjxwWiK1
KJydZFl7oDY/Sg5HzFO3cbbOgkKGsZqOjmyFOVlldfPrbQ1IlG9J4RggYL5EaqMQ
l6uni27a29VQsyspghooIIk2kxQtq6aGsyJz4Oewb5NVCdp7PH3SHeaY0qj5XtZE
nnTHDzGzZudT6GDdz0+jD2+ZqhV1S/7mQNmiQjb0+tXplY4RZ/w9c3MkT6a2Fqi/
Px6fSpFKE1fm5nwm4vdboNZNCi9z/EMYvSZWK3ZBx4hBwEnpaTNORR2vBxCh2FOc
cwYngyxzMFvFhasqaq3ydS/jls6sGNqbqsXE0a9XRMsBczUufIaZSHJYzXpB4Jzi
fx9792VctvRzu/k8ecIrDzh2LdXIPkgVKzEwJbmh4JQDXr+QMOMO/yZd6a5yQVBa
7Tf8A3uSob9ZdwQukNjl+hP19pVE0ENrRTx16g4f82UdMiLGF3xjQxXe4b980dt6
LHC2y6tfPz+oqwG68iZZ3UeBdi4w5wPeAJl+vFdo3SnzztUHlV7oxlTdqERTiXOc
LciYEBVKh6WVand4SRARunvoJoPU8Fvj5PgFqhWTrdw+RR35W9dMcTm5N+AzxKRW
I0EJ+8ZEgp1TO7I61Tmz9OjIIhxGsRD/F2Tkhz1eV87S/8eyD4+qOjcsfVrPwgvx
tlKWEjT4fDJjffkC6LVtyEMGAQw6duRfxWAXBPotz9yrM7kIE7RakYNbYhH3Mqet
lXTJg9TfaB9KsCDi85Q3giq+ARy1e4eiafV3UZkvgE591jN5WapuK1EuM3XZt4pa
FYhHAqjo5DrCS1qnl5Wv3EIXlJhB3gJ7pdgwfIh1g8StnqTk4pJQggtADFEEAWjH
NEX8dX31jGg5dz7PgzvbDLs8om47g/IwHGei7hMwxlNsMsVofUGyOLeuQNHuVLub
mKHN9x2tf6fizHrSezIg/rj39AFHriDW8/FJrdXPatfXFYO4Ks58uWRVbPa6UENT
8UQI1PqXDyBd3hMJwnCBJytR4l+EoJm3H69gqlg1wpFr2630hDcbTSQ7Q5ArZIcv
BZh8mE1IHu8FnLgdeX9iNuaxV7xUOq3BDWAPnKsV3evCMwUeEtTraCIj63uWLQj+
UhsPnSX+vBKwjjI16mzeLsAiDHUlv2J5jN4Ecu3ZWsTXlySDrdhXevctpfgio2yH
/E8hU7xM847esd1ENxxTK7L1Nns7pdnt4wlYCv1L9ettSVUzvRrDrUsPB0JBaXxe
T5z2ByOBRc/uBboS0IMuTVbQysEl+T55ZS4ifnf+n4fnwXaCKTBFBewmLpvpaOBK
LyTa2mTYnPm1udZZ278NQnOWqcAdEvnL5LvPmXie32lIJ7T/EUrNg5mr7EzWazAQ
2V9mhIqUA3U/KtC3nfJ6bmmKdD1kHP3loqGKmF2oc1IcTS/5hoxrjXVEofK5NGcU
BYPgeQAnZ7a2+N9hGzrlv9hPcBepalFLHrAYeqQbW99B4JNWBdaxRE3pDYJVrpZi
SiraWHf0CxDcVa4hyr67deaXBcUU21F2Nd54DKBWoKOsYM4fqtWJO319+4LxLoEr
TjK0b46KmW9Wr6l4CCE7qn6mX2xegiZO7qO7H0VJiQnZs44SjGeX30oP6X0u5jXM
fW2t+IC+DfquqMEB/u1j//kx2o2IWcMCSqp059qRhsPStrrlB1ENcoHEtO+q7zhx
DJiNm2sktjP7fYRHlT9DrhYkgqk16IZY41zFHUvIIRE/nnREYatIay6MQEIxF88S
IoFS5a30JBKBbEhYHDXdQ7WdYHcBqrm5hE0NQ3Wodew2JNWOXr5IaLzeD9dzINOD
Amh5/f7/mEQW7V064ElX9hIgxge3pgtZ7fX/XRcIbg5zW8Y+GGsat82zljaUHJYO
e8VOzysxqvJsj+8fOdbiUaDQM7EEEvn1fFn2xYilWV6dE4qS6FttiAN3EWD4Lhmd
wE6fuXG3TUbCg373ZyV65Tqsb8TRUPMzLatZV6NO+AB7bW6e5WqXzG5AkYkE2xF6
zBgCKCd5JcmWiD09WrvkFT0kX5HC6SYKGh1od4tVPtGFtXjQ5q3c2K1lbthlicF/
8NMSYfLE1JdVZEcRpehn92i0mcAI/ln4SJJLSGD7k4VVYTT3X8CKJGSsd+8ojDOY
tJyMh4tfexCLEWqRcMNKXTfFjPQfqRE0PtMHMNAiM9BiDEZvCSmOAKTUCeKpbokK
GBRTIkooRmcwFonE8n5l1OLYS0ELliipEBl6YJzRDL0MJWBW4DJWoPoWKKbuAgu0
wwurSTTdtgJfojrTw3B0U5C2wMEy3P6CLh8XpcGsrunqwrZS0wOpZmPOmAlu7cUO
nGolsvGcUWwCf0S135EniQqpnCzhiMNSG9pnvbm06Edo1OdSsT5vAyG8Y87Hxj75
dSWOD+KdYCjpuj7WRkGcA5EqWsvEHidP0ZvHANtw4lMphBUiuYNYDfOF2X/310Ns
JuWpRWS2XldEdrrFsSyD/97jEDVyh0BkYvjSvXHSg8t1PpuI7iITEH9SJJn7/n97
ATQHwtkiWN8cqdmpPlkOcjuQtvysdRD64A+mtSO9FvSSpUZEl1ctjgth4XZW/HKq
d7/iAhGImcKD7zK1ydElUlqlptrHiLG+gWGMdIJ1ErLDaPFJwFXVnTjlWyoJkuFs
yT9uzhesxQvZMxatwy3f3fVP4xwCHefCzwnKbf/HOOpJMlpotlp3NWnIHUbapLl5
wW4U3WSakbcz5D+k9kuyBwysBnqUyzHY/C3kGYQdnfY+VBjWIle6PVUKimWjy6kb
OPYEJjNQfq5f4Ijqfm8cm+mNGz4GpNAKfHYAILG/h1H5wLMBQRcowCWH/+SJGHS0
iDVamn1cBwI9D7PEcxOYZNQZG+vucLTZ7+02VnbWSb8wHcDEyqfjSv2ge0aw4spb
qOZumxB92Bv1YIFIgxYVgIP6V64sGVF8d35ikO+5zNb0ZGo2Ok04NKdl782MYPoe
c2YN1+zHnF1YRiGZSH8OU+ZkAjkWDbIhNLAXZbgJSvkBOJsdHSSSntiy3EwT0z6a
Xct83KZ1E6kiweQIODBRNBywELQROYHdL+0wFC4HBSffohSe2sqlxr1yfbR4fqsH
vTUoznW8dL4aJPmI3Ex6zcawo4tnQeghfQU/NQSeC742hnzSrL/s3WR+j+HHRbW4
L/HjnTsvMi62vzjEdx6wkrzoMw5uprYA04YR+7XoOze7zsbtXTeY+1ycaTnoxXS8
eLriJDcym+71ovV+IushuymxlczazGMlzRVkA0R+6F90O8yOIO/JYI8MGNrK3roT
fGLQm3Bxbx5iHW0MDcCRq3Rq1q+3HWDcbL6Kb+SN6bvWJ9acnfLYf+xYTxYSw+H6
dn1ODv7iY1tsVfX9YePhWwsn5KaaGqmfe1ZbcuToNYneaGR68iLxyCNz4NjUp7rA
vUGdZ3iq7Gp0G4RUWP+du3IipTmZ+Z0jivUl7/H0gCohcqbKhWYzb1xSUqYArL4o
3Xz9H7aaRdXrviDGiK+6BwODGwlonVac8nqNvWLJU1q+x9A4vgfA0DzrGKwUjULc
WPdoYc4iRG23vFNDHOGvm+v47PAzgcjZvVWdvQNM+l9KHFBo6op37fr9Vhj2vJUq
axuJaj/FsP4W6FOCHP4yILW+e8EsfOU9shyMk8uFBMxPbFL7gf2u30L4DjzWAZPO
6OKzrVFUW0SmS7SAyyXynvZ1nYKKlH1kiXLq12Fm+5huYybIch1N3DPbFNuIlEjz
1LecydHrlD7gBnB/ES7qXJ3u4vY3dUVZFebKANt9qWgW1hT2xMBjqa5nZhQSLFTf
jLAzY+/ip7hV41mXIRg8IXSMJNkw1Lfqhcni0aCqCIfnclhaPXJxT/ve7ZxMEysu
23GQemJy2UkB/sQ//bCU1WWbNArY8h2ImTwkezo45xIybOUhT+AzlklUHcXOhErk
h9U1APoea9TimiidlpiKIcT15AR5JTfmfRTlW8aibr6kUIuMpTpObV5uM+GtX1oX
MdxCBli1oFXO/n8XqmH52qnmw9jipap+b6mOUE1ofh8q5Rbgjq1E/FBaPaO4KEW4
w/1b1JODXlTzpTOxpylTz6/Yv+KbYdCANLXGA8wgzhJlIk/c4wXKVK2FOWaPWl73
A5YhyAUf9nX1WCf7X4XkaHpULSkElFjCLBFobQFsfWNzcq6KiJ7xjxnNXiZ1hrYG
qLAHSZPmm6RH02xgrtmn0aZ1VTImhQEWSn+MHpr3c46baEH3W/AOzIongu0tvG8s
P427Q6nQxzh8hx3BAL018OoFwsPsD+Zq16Gl3qf3YhDswnho/m/ErNuNr5SghhBu
oAcZulyIOIx4wivdDlvlQjh9Ytz9JRXQEeaesulOFXyp5ljV8dTasBeTxtgmGwqu
8UIK1mvR3h9ugPVsLvIxKV0fgEWoqHb0pPq9xnKEh9xaQF7XvA+bo8JCToKmIa67
A6kBhk6GW5CrE3sJOO4MnozCM9fkWthc42f4X9/NoV3M9AcUrdenjUGFuK6+5ySP
n5eSfObQW2wxnX9Ph7Gv6ozDAPrvS5z7L+u0rb1l8qZ5syTOOWeMSxD6qyXstMwn
XtAWioPAy8IAEBpFJlkFLEV8rnkC4JZehxZbmGf9qoy6DdybbG3KlAnamUVv+xZr
RkC8Ethg5INPrDNS7iy7JrhMBdW94Sd/VfDS7OiBlGUGPQdFs6beWFTyPRfgCN3q
nWILOJSA1yutarMpWxMCYyKyEKe8n52g64Mb5H9Y9JxzCQEstIPeTtiy5x8QBIIz
e/o9uziJLBr7WRj5zy5AJucBCJV4FaMXj8jm02DI5ogFfl8nEi6E0/sMYS2+Xx9m
L1LKUknZ6/jTgOHOslvDfeH3saCTfDXqK1xK2uYLI9e6T83R5Ul2GJULQinAg3qB
iITlxr2DZ6xfuCenqDc/rsHNp7qk9h2/5hjUg3KzQb25H0USk4lhaJR6TKngEjpG
RqVTJ3yx3z38xblJI5X4GOdA83mXpOaqbsCa4hK72wgnl0D7Uw03E8FvZjfzDM6K
MQNLjjvwijSlWn/DebvHP3bVX1FacCPigoJorkZJ/pLIGrw6uHa2h9R5zk+eWKpM
jF6RoA/A58t20lG4oZa42D5HlTGTQsp+zlCVddPfizHpf+kQJEBueKvwej6l4z6t
kEBFfDF7VxggTceb/RjOHgR0YOCfAD40zwG5jdgnZdV+1Vho00++BDKVxFJCJUVP
CFK8+LsP0vAPlETv8xhtS4k1g84w+oGIpGCPJjqBEDaS3FTAecZfla1nrPwtf5GC
ZMN/LvNbRI34wOYMtV7thyDempZ5TUXAi4lm0cNUyldgiw5Qu0uBVLcinME65kyG
Yrx6vmIm0F7fgXQU0lqCDC6hV+oXwDuP/RP71uPzPWCHbxpvkF7OEgBAxtIlyikt
87Da8eMqH4PkTiQSIAOFj982crXRRKDcrR785TcxzWaxhYSuK3Y0CYXDLbwZkBoC
6augEJvJx0CY61wZiq4+KL4/5AbcOz+cRNFgUDT0pNF2SKZ8Lafb1/GPjZC/ZxS3
oRIbwNGHVR8KjAouhff3228yY18Q3lf4QwCGUMgSkBiRuNE/f0MhWV9u1hTCptQJ
jHXq57+dxTv5DyWCKGWYOMZZFVRRlSUF1G3ZXgUaJ1Vl71TVd+Kb2sbk6aW7fsc8
7HbzbjSGZ45Bam3bf2mmr0VDh8BKG9KavFyZmpZX0kiShKj9KOy22O6A8j31iI5i
rHn1M22eOwPN1YbEPXsRgWClHO1nEZt9ltCOwJ3z89JlcrNGb/xrpsJomGYrvizZ
huOJr2oW+hJAr11nDSQWTB6/PKGtNrGVa1+93qs2CYPC1lx/ycBqo9U5v9Rmthuv
0anBkBjN8pKPbj7UXbixxPpwMKVKoDD+I+GjM2ZRpIzp1EC39u1nwJckOSskoy2V
9WAXrzDz6xR1kSyIp55e2Tk4qYDkWhgveixPFpdHd9THsiJhmJOCt49OMppo+Cuc
xoD6k/CMHJ1FFQRhIXOzYS2crdUjaw7IH0WQgxXRH9vls2+4dk7Nz6S5gjNAAQeq
r7Vrm74ntZ+pJ/7OjbUm1dipVFuWGqzjbHUBrJV9grDqfTT5xzlm69Otgtsp+Ydb
FWRYjvSlbQHYSn2CTIHnKl2nhs5ZtT7v23X2kX1LjaLFGp11oOwQlDBRzsELSADp
u3EubQlB1XOJ2Szf+J1HQb21vCIpJFmF9G/7CukBRd+OiuyPTMKuEHcsInrfXeXb
6Sfyv9HVreiLwJKqecdSGBsob9Il14t0RcbWc3lRULXDzK7xqfqcCV0/7JV5JNpJ
9WDcui4m+NwTmJsALNG5+PIR2Xj5NvA3sYHrQESPrXMND0GmWx212WT7s6XNpWr7
yKdS3MF30JAKHRgUkYYR2+ZBrR5eQr/md8ifal5onKCM951IPDLgI3CY9c5HrLj1
4NgYN8dZ5FpkpqS31K/IK8fpSi25rZnlWyrxcJfxOQ5vkMEKdCziLyY0KpB9CFRU
GHV8IxqEC6IcIxZADW4bFFFPVyzNAn1z6H3NIer+5AvFQZcZe972+lCntPqCqZjg
djz9Bpp1DbmRCJOOBCMQzrO7zBJfG9d4csd/yXjobcTsRdXY5wtoBvRMvBQxjjZa
j0D9vLpUHpda2K8lv8olUhz5BylBfiEHXSDIA8hDjey8vJhvKtHKortnpqBEve0X
KJqljHOvGqJbyj1VQmNLV3wHjZFAmQzYBtlcrhp8gEIO4aHmaRo1kYbVuDTo94XT
HCfD9anp5GhuMio1qC40hqm+1NEVyq48zeits5K9HOrskdYGpo87iNZKj5+4o+I0
zLDXwfyWgXErD7P4hFCGhiHsjRhN1gSwxZu+pIS+fjtOMdr5yAuDzhrdT/s6VVPP
clE182OQqRpDACk/vdacFQs5TvFaazfRQwI5wmWgUc0KuJlYzFilLwK+17tShLgM
4EICkv/8ctw686xEzW5c2N43P88XPqvOOxTu3N0u9KzuOHz8sgLydYEmU//CYc6z
dN9Orj1qrrafrxcHddWaHfmdhofY+PnpAySxCsAOZ/2yJjFBdIv6uDmWJkg3DpuT
raiEnbmttYC4+VXKEXQ5+gV63klmpPTTfryl7BQDvFePsEz59kQfEk8kOSNEudoI
arJUsStHTS7/UrtdHwZEqWJIDm6kCka8WPq1PlYCKWI1BIOq97Sj6eSqvZ2hdyYy
GztNccd1gxZZIjZUDjzByex0Qgl78fdhDSYKOC8iARI9bUFhCpqcgVJFy0R/Yn0r
1c3iuuiyiCbtnNbQrLhHJymO669byNg8vgfxziptEZpOVBkrmVhC73h5jGAnVBId
qEA5wqr6cx38F4CsT58hW+/hJeqI+dq+bq5f9gE9DmVnuTfZ2nWo88OHo6jRdgnV
3x7c20P17XCZchH2fZ4m5Gv1kbKA6ObJ3ESIftbWYFX7wOkQE6yDnSnSIWmBivzv
kpJyLwqxpdqnRV2ZXdTZypvxjQrBkuxmsJH6NCGAYzZs2t1O0MrPsqTHfPR5POVw
Dt22P6E+W5UyeT+OL18HvLwAnfHOc8KjM+jQnnJu0jSiRISTxSMdXfrS5TQGEX06
N8mzK62gGsRY1oLKdsvzTL1bbUh4FgL7VDFgw5fTAqSWlkOSpqcXsOraYGfQ6bFk
ylYCuPa3Hdiwdhi320n59+eX1sWXH59CTVJTK+bnKYzwcouYVT+SLLToFr9wWYea
fEIHSYSIqV9rdirSooXsht3QbTb5A4MN4pZ9mDx9El14ScBMRp1ZVds3P8wzlsK/
pXTEhp+r6eTtPVpmFm7IskhZh4yMRXtQV82P6DXI97JFApgLHl+2sMbRwGQoVPjC
P21UtLw9IzQeGkgj1U/IhnBCYqyYDjuMbEsvBD4pyzAgxFAZPlmP7q1umWRTKMxg
TduRuVUZgmvaIytHmi0X63F6W40GqFiK61vH6Ws99Ydvyy8hViGtoAE11TbmXSD4
IbTm9qmyJycwQL0SfPjlctgTbVB3a3nBcN+8e4+biaZW/o/tmXrGfM9gX05YHUvb
LJ5hkbZPwEl0TZ5K1NiLQL9mAbReUsvEBrtdLqm82Ue3N5NLVvK346g7O3zR4wOJ
ipCOx20vFcVG/chnhUzRBLHVPA5Tv8cP08V8viB4xY4YRnkE7qlwp94nfmS93jVx
ENNaSkLMDZIG67xnOGlpMxJUXUyx81hIHffvHTjALQ8oXdN9fMIglsctKeId/eEo
G3Y9xORpicKR82spsned/Ys4TfUe6mJxBz8QxYx3LRERsoUlVj9vwi0TuEGkvIxQ
QmLfmI+AnEYzGK4ICYSkfnsKKYyjOS+PWu7TcnMUMQUVP2IvT5t0Yr2mECToNws3
bnc4eLzR5RAFrpLz+4C33xgoVFAU6iVEZXBsqbolt0lBju21yFLWBMHlbjZFQh5q
dkwkC+RAZTZzBnol4jdEdu/LM+q+JyBBbHfWY8HqKsyMRMha/tO9PfTtrJch9sMa
U+gJgWikQBiEPShd3N3/o2HLJ5hAlGvBWoiRftx5GyAsHjP0ifTQd/9Glyd/OwT2
+0cp+QGcCqOO4aOrJC7R3NoFxHJyWXxj9SEBh5Letc5ItS4CjC1ofdI+DV6ELS0k
JyHSveg4us7018pp9oBK1wwHUTr6gn72D4FM2XVA2ZQvIWt4InpUhIF2t8TCfcSK
wu0Z+5uJXXEAQ8jegw0iR1rDaMV0LQIS67zBavVYreTZVTxvejMuqFyFzJm3TzlQ
tmpkhV2tlVbAx0wUHt6jxOZkdM8s8IZ6arnYaOS7l0ZW6E1a4PRsZfA33USu/fQa
Til4nABSSA/DLUcknSemeDs8g+VB/uFp7VRFyDXlGeg0Igk0cjAwMiGmWy24+T1c
tQBQM91K1i1roXW6Hm00/uE/piiDrCMscJkRpeKy1Clle4w2uHt1hSYWKEno5KBy
vEpXFmNi0qFeKog5itf0/7ccfauhwsZDk6ejOSK4Hr+Bi2XXftd2IOKm35AjHvvw
R3hVMS5t7JUBFXi6L7keU9W3fzautv4qPNj8rxXr6EHkyyFf3mNevT9iW0f1NwH3
VmacDExHeP9eSxKzjmXzhGIKvV4P6mycbCyrPcptF5/6opcDxOAkLLMafzMG6PAH
jjAjO79WHb+WryuXeqtdSHNTteMwRfiCHpUb1fW/4tU0tBdWW8mJl2Jk8HgVmCb3
DvARBgquIf6NWRZYahHjIQOmJV5w9FhPHRyS4yUeB47gh6vw0KjViU8YrMTMBLIw
QvIyPi/brytckJx6rSgea5whic3BWnYmCqz2KA5OJZUIS8+zMfXvLn9cSy6jrWvh
t52EVGA/AruRv0Q69N6mu90XrbVGDLdMtHm/YAyyClFmQt4fG/j1upkWjqQP5GFZ
5R4KyILVd0CjDoY0CKeKAEkpKlWOtdiWkbHjTsqm87bki5w4r1fQYc2Gt2yYkO53
MPYUTy15xKynUzpISk3MR62Bs+vwxCW4Xc8Ebl8W/3FW16zWv9eImbiC8ts/g+n9
RRMHMRUmtw5KGbqU3MDGQwH72Xu7H/yfzPafufiMtVTzxfzNsv6du3ERW9Aw0pXw
29sTe6rWVdNVQyxD7/ZI5Z3SA0qE+4AtAwpLA1OwOoMUwNHqHE+w5Y2Y1ZI9NSjC
uEeAq4CgCNPQt/2vc6JSRZDTitIlG7Dph/Bcu6QfAZPB8o45fXWfHI6PiJq1lOqv
pB5ywIK3haro93Ps6B2H3utD3/6gkgqsi3xg8scdJCUJrdZwALvGvJx2Yb53lrKJ
YnPZuYwyOPzRM7rlB8xNc93JlFqaa9d0UFDS9FBhELo0goS/2dn1Rqg+bvDEw0I9
zwFssn4Nv8UACIZBgh9pqUU/qJDmVgE9uKW8XSiHXdc02kC+Gz4KCzptjlAqA/xv
Ohc6mjqN+x/QayQSPkP3L1uo2/q36cxxtUsJ3EBfkVj1StM431tI8r605Mopr7CE
shUwlYoWchfiY88OZv7Y4gO7Z62EV7BUKwT+tym6KyPPCsBIR6Pq1mDJQSJhhBfr
vsk8TNtkyqQNORE96dtOE63p8sPzb9MN6kR00+OmefQZ5aTWEl4kfP6GuepVD3GF
sQmda58kL/K6ZDnpiBxe3x7sMjmrCABbwvypZsLnzyfhKWQAJVREjT08L1qG/u06
8i59wcfkJBmt3LlUbM+WvLmVKN++KEZRjANDMxoq2rGZjDd2UkOD4ucbay/DSpXk
AcQXAGC9Yky53z2cvvspCx382BoZzVmF8xTTN3J762d6IU1mVS1p5QY7DNEyKEkW
3nQfwpStc5vBH9vUtduRxQM5aqD8NVbCD4hbpMZH2LioxgIreCbTwufkbnJ5/29o
/zSpTZwQHu/FaWb2Hkr0TrPF07lfbOYdRD7tLUcB3LtB7AJU+E/E5pMs/2/6KQEX
RJOjYeyQ1skOuhh1pypUaDA863rBSt/PMqUez/zusRHEQOB4VvWHEp++TvYjDbaR
1Vh9hnbl6hfXk4tmXXe+yFtznmvUCWmpkchaO79rDuv1hLi/1h1/aCy6BBrhM9N5
xBGlHI3LE8R2T2Y0c6Q2637eSfwsK7ic50QW2Pq4sDOHIKvbfuEYDyFfGnns3DOs
r1gewG6725TEGAnoUSuj21DKh1F/+ErfMd/g47j9RAYpDEIwkfdehKNf10EDVpjS
95kNfXgPDO1646VlNUCy7wZwX307ac6x56Nx1wTRh3Miyw/gfMYMy52SGbsCd9L0
u9om96Og52OIQ4DXcilB0GSxJPdn41Eq4Bm9TEKFFGG8HoXdBv8E2QufxCovUDYO
Vtz691PcJE60suaWlHiQbScwFOpWE8bQrrOZhuMCGV+fuNdgzSfoPe5yyaGIsuBQ
IlKLX7NJ7UzesS2la1NgLanUhGGiwqqVUSPRopPGTjX6Y7bF3cudkPnXwuyEiSKO
TJIequSuLCaTtSRNWcc/bxaH1CZz7oeCauw5E5hT142MISuEdwK/+mczEqLZurmj
kUi4a4strmxCN1SQ2NW2KlTHBCdn3Uks+5C82s5t1NmHJ7Zvk75bNF6rAgTIAtmy
CJE/kBFfhDmPRu3BPBoKO+ylQp7cAqV4bMG+g0/II70uuQygvtv4ZaTmrl1QctSQ
1YO7eDo3czEYFoBTuwioZuQM2Z90BrMrDrT0upkfvElm2Xwn+K2HkUNWPoSTnb9w
Ee45LDMBGd4xSq2a4dW1HqZ+1DROcYQ4gB8j+XKJAPI7x8wCvPTt1VBeXs6bR+6v
d1ecfkPR5oa+ebXE3RxxrSbnHILOdHnLoWpwx4JoQbg+FEcMsXmonejleMJzwGlr
DiSx2xbSNlzUYdZsYTMYBjvLHQpHpp33ElyPxh3Ug44NmxSB9gq95l9++I/cZ6Qv
S7AJzi4mPgAJ9bO5BHt/EF8yYf1MVALIM5r0g/dKjcqRu5MlXRW4rjVCvLwDrWvD
6o0cFEE44rqi+6zonxg9NnfMB8bIL16Q/CYuUKxFqs8UAwgUZZjjsuoOqHPijmKs
WMBqsKTKThDxluuZvj/NHH6Q4CX9aiH6RogVl8Mj/HaKh4XSCW35PX3d1cW6DMNA
v37gqL/hc2rYAPFvGeazH3F0PZ7q+xtww8rXQ5HUEhstGgJxS9FItGOpgMbHRNy5
5RR+dqZbDo8vlvultRT2cinYeTzSOb4wIlKGjB5G/HH5kbDC05EHMPi8OZTgEg/a
KmQ1VGSuQ/2eVAdUIsEIqHPHWYvYHgDcKYrji0K2m0O83/dUenoGbX2RKKcRfni9
PI2CB/uydJDnTYv2+tNXeggqic5GLeIbue/0l/656A/9Pip90cn0NUPe8DswDwnx
vhdqw3N0ZhQcl09elaEXfwcTK1wkfnHeJZ9KLRHUBlR6Tj+rI5W4/P2F5kwwtReP
4IpQ9GJ3NEaLv4PKiabCwRfiJhm35CMksYlbjlZPJGwW3XUmwXhTlZexUVYKXjv3
L3F3Qlx1lxAjvfw7ft3ACb8zDLRpZA7Dt02C6Cwfq8JqpmhgREgbSepzFROo4eZF
q2TQYo6mrlE07SeNknxUOAHl+LnoLFZLJIUAqT4zz56uj1Xayd58pCORhiZ+CYxT
glGBT+3N/jzb31uZtGhXEs7m8YtaXKWRcIfmlH5TIo3jR0tKdx5+HSHq0EZk7qqm
lvVPBjZ/yW+crsIwnGB2Bnzpc4PiGt2YZERYRH4cha76lUcnXXQ/EvkOZvLQgmCt
/d+Tq9yHBksNitC6ikbT7L7/bQCFtsADouKatkElSNVVBumQX79/4sKydT9/RE3V
2zK2vIBc1p5Gv4sswA4nXnLQA3fYW4liisktOn0WBsVTaLaDE1UK4D4vP9gkzH4b
/SGlS/qNhsankL5018MQthwK7o2vLvVE8f5EuegVJqf6mq/7zjRnw374KGmYwf9x
7Y0MeDZ7tl9C3Th/STnoMlkdAadESgUyrwarooLZSEEq17oZR5jfXtZ9FySfayVU
9tRS6Db6OwqGnxqOqwPYR2giZYRLP5Kk9KBSr34vfcowW2iGRwlFHC8yv/832yNJ
oyBLo4iqurEmuCjxvIVGHfw/FosYxxVpY7qX+klQVypua+V6TopXQpjdnXNgYpY9
Vxf791dBtbM6xrX0l+3pqH56SIFsU0CRCB/SQTSo2ZGNQu1t3ORUvfC5cs3IvFOR
8iMGFt1LNq45aAf/aYx4dTxlF+Sp4SNrKm+B0nQn2JfndoiDYy46lpG+e85z3REr
ir44RGuRXg7GWFkrYZFOQYZ0Fr4vxsKzj7iACmyXPac7xQMz3vdqKXAwzD4q8Lbu
8gNiBvwdu7czn545pEBt3lnwCAH3i+TNKQK9zjR11loSFcgTYlJlGFpdaZQThzHV
FDhSVebAIXTbRkaUCsOme0bWpxy67qOWbJc4UuB3HTVeZFQ2ryWlFD+irHvVkn2U
JoJ9np6pb9/MhwV3R6Ncv81LzdZNzy1G2FHRSlt4mMTsaIylbylJsDMyRFSQGatu
TVaFgUHW/pVpMpXXZVTlnIEXzGV3+tjYDLYGaFYUb/RNwzguCv1KC1+hCNzMm5/Z
DDhgkUnhsCyxIWA6T7p9rboO8F8OAiU5JkElUrN5/bBSZZDBxdSH9S9sMCgvgflf
JWVjxkyJ12n3IclWIrEvqmyxa37/qN7NTIEGBf0OS9UkotAajK79Pp9Y+Y8EyPvs
04Q3QPxjZh4z2vNOoC8Bzinz16LxfzW9lRRTMYxp/9+L+azbknclCjwcqf90ID5+
i+3n8KK8kFL8ftHDAQXYUhpwMNy5en4uOn5eq0vW60jOkEUnUkuhly8dkE6fZ5LF
PERFL1+4oSU9HnmSORJaWhmdaAUWrTCtnBWHhCo+d7Bb6BR7z/+ErvdmjlIjXsM2
GRqW8a4D7SYkTtY0TmbCb7Asj/aDNip7c+piDwyloyNb6kIDLsWvudRrmKGEhpNn
aodWlgtcdGgcTHHhLJJrWoUg/n/ZYwkDttR5ssQgRTQrVdNXPlrMke++M78rb4rY
nxGuod4mythVisrJupHf8dZLNJauygNv3JUNjZiacVsWgc7XEMg2OxdU6wmWVFsx
luf3daO03TzV9em0iRyCST20fTNqfOInbuPtXhA6tUuseZBeqEENIfVazMQr+kPr
4EC5Sl+QzynzT+WBdG98PcFtSG0O3QsJz5+ZMRhrsozqmp0zLq+hSGbS/grXMBre
fYIUJd1gl8qq8fgmFMsrMNFQ5z8LUeNvG8OCOD0a0PfALHMFZ7daTJKMontZ864B
OgTjxT18hKICWnjpY8yF8ZfJ4ur2Xb43cCqvrLi9CFOPQUk8GCvMlVZH3S7g9KyI
y05ymCiQVYNbNCLOesCwxxpF6rNtiZKbCNWZy3mOGnUb6Am1LUU7pQG7tMdLdqA1
Hx0BVxKpWOsxYXs9+dQngkZWIBzX98Y9xDC23N/agH9/jQpTxh17rTz/DcgzysPE
tdHKSryvTOZgZZQfLH8gNykDm9B5xcARwgMI3qTmqAzfaxFFVof6yYV76HYT3mVh
qrpVhBxTeKeyD5Rfi4WJlg88bk2tTruYTSP6E69pY6shRH9peMbyiCqsnJk2EVnt
psAn9eV3Uuhk3vQOigxJcTKIoVYKs6kY6QKNJXQk4MeZz36HHiY/tyDyQte3X1GV
z7WlRYMZEbobfkHT6Spwdqy6fIpUdgvSHBOnGpoZuWlbmdOJYSYmzsWBG7eaoGrn
ut2kIERqIlAwwf3qVDafZC00VNS/bxybLpeu04LPFLWqkuDihcL4rxoAyptXpNj0
AaX8d6DkKXVoICD0LtILHuh9P4gOFixUyEj5PLEwgKZmdqA40x8S3qEKZVYXErgi
OtCAoIeOdDyR03U1ZPHo6RBPa2aHaYRPE9+3uNyt2a8M8ReyMqeNic5qPsh30wsI
75R0hB/C5DJTEyd+oDJDEDjpJE5ToqH4r7AcN9QVVgIwpf8F3JgPboF0VQdxaLdg
7prFbfGsOfVxVlqgXJQl2YyQ4xQmoJuA/NoH58frQ4wT0g2eLEDQpqw1zbe8i97o
Gml+z0DymVcaG6byygQqSC40Kg2ImcaQkEpR3I+EBfv8II3F45IilmmsZeChKKGE
sQEwb4yUVfiKO0T62G06dKtJuTeNRwJWhN+0bfOuZImxp8ePvpS2DViHEZACrU+9
UvqeAEQlJGlBpj7pbJVVf6RRYXygISOdkvlXIJ6HaV/w80X8HU+l5R7m7w6REhyA
hrf0U3t6ng653CHZhOWERKplVNmt0aA/LhkENC7liyE6vZ9/tplR0TPoAQ/yGsg6
IbNdGjvSob5BAMTa1KovP9y3i5gL7rbyAHyaob166AyBTPxggehvQSCgyhehoSGW
IiiqTi8NGts+kx/oU8bMs9cmvmNknrmr7DhYeXzb6KBwJqCidrsR17Q2AVIgHt6g
8HJT/Q+QfCrKLIabJA4fcli3xfY6P4HvfKHI1d7Co+aADTw5FQuMBlziFhhZGsnc
meuFviVbo0RdUmFRGJNK9HNmqKZboUxJG+CVbsvY94mn7lH43WT05uhsL4PWAI0F
6tvECJiggOpFGKOhhuIQkytlzqt9G7bziCdfdWRTTOY7zLhHY7Ju34wvzPG/cAtJ
s0ifvHrvcf9KZKfu2mTV8CLd9shK/uOHmrvnfaQq+rflmDJ2KMNtKxL2J6IWTQZX
2mD2g7UZ9aCb90/CdqUUU1gol46k+cwEPwyH9BTymGqDzEt3TKSnS6V6OegOBsJJ
CskeHo/oiQ9RhgxANdj/dLPpMZBNTc02zk7JAd5qaHpyDUI+EXCfuuml1GAxCvJf
940ih8rNCouGM3icg1+XeS2R2qmSKxAxzLaJgwSDJesGhQ13U7rKvzD0/gDeIFOD
9w/qMnjmu60jKqditcccgx/KVbW4lzMeSuIz+6DggGeEIBPN0kCAzaVZpMqJml8c
MOt67VnkVdrX3LkEcncPZYavn0Hd0fbToynbJeAA26DOLTcXq9N47CDRe4CuUYGn
wFa1SaaOuCpRBpjn4dbwkHiHYO69VCw3zzN0akGW1gxIZdvqGU0RqiGvB/tsWZLq
8PFCxx+TQk5HPDWsU5vkiENMeTfUPW1a2uOGiFJl9MMSDejkGYj2fiCU87TTqlYf
5gm++RCADqCkdrb52e9uYSTJUWSz7NRiNcRRx2o41m9+HYUFe0qQDhaxjmMU9PTO
rCMxw/EC+5qVpIsmf6R+5AwjAQtiwhHh+AyKVyXp0KYXV9l/W8FTuRlnx4Vi4wSl
g1ep2IdpkK7boc2F2ZuU3d5+iTbRPDna2tUbqzbXTFeGSF5+lybJbv2+98QDdTKC
nNsW9K2mevAjkL8fKfPKx6VbsyTBJzBOvne0E04WjLahFuawrP49rDt4mS6nMOMs
GAx85WgGkpUfR+/7+FIwtm/Lj+hxj4ENc1NY3VGZ1KVpcApBPuTe2Y4IibGDfqO+
WP6jHR+Jd794YdfZzrbX58/sUBKt9DadCUl265UAThqW13h5BAZ0qq47b29Pyve3
CNbC6f4OaD8fnxWRqHNAt/8sjd+DTqhRKUnNOuP9ZQlMHDtr4T/QIuq7R5Y9Vu5m
zSP2lHUQc8zhjcHJiGnTX8nFoL1+h2cLrtB6dsIvaF0AyTUElhESqifVltSoFyQ4
T9kq64vkelXZsnwdB0M8PqpQGSVhkLnyHL4KDbDfpW06G1/m8DJCgoIjiNnOd43D
MVCOAgmUfQ3p3uC1alk4IBE2xGlyRaOU9MO9POUyx9K8MhUH0dkPoNQW2TyYDhFB
TynVskyTOXN3IN42xTMZZNmzVimWA1k3rz43DixX/XfvKNqoyfb1JjkeIXS3E0vc
i83PkbM0A7eP+XThzviZwkJfMGJmshOQvgtK6Ox9y3V+4JC1DatDXo80Affnk0/I
QHJ+qX9eLoYdJo7GL0v3fO/fvxLZSodfBFvTL+TIitMjsnkoKsx8YESWY/aiqa3l
ur9SZp0ZMzfYUp3ClRZOgRV5A6eOOuDSrSyNLo3GUWaKRz0KP2pLrpMWAxqxOF3E
mMDDmWdSCowg/cR9HG8A26zAyBYjM2xWsYcbEPXPKXJ0SaO6Q7QUZxeDXdQMrBzU
maf+kkRWorf0IQpZM0PgA2esl3TEKqTrZ8UoSYst0qKtFMrhrG+VpX+pTDQTjM9J
tKomkiBaHHpZy/bVB1JEPmaPcYd1u0EuXQXtvNjq7UkvU6I1dPHSY64ytrbKRSbL
4/2x2wuqmP+PgOikk9mUx0eGm9rykPm0ZskS+o+2hR+wVpkDIWHfAUzPVhGe65mN
YD0LVZ9w+Yg9Dd6TiQCe/VyS8ILMOg1fEUettfJ8aw0SaW14xo6qp6L6nbiSE4gQ
fuJTFDqpiIIr/guhw/+sQMKtQhwgsnCYFUwwHR4UXI5cV419QgB26wtsjaF4bA1V
DbIM7YuH34glC8czWOedpTPGX/RLb01awjIHlVY3sd9yOP6N4PGLi8kU5dXTe2dg
Y0mxEg2ikUxc6KQJJEIdTxaEfBmf0ZvxjFrIM35PiUDIhEAk9eA99ON4fvKBR8JC
gW3tqoOXzD5qmFZu/tr6JnQZnappN3uAwRtK1dI81qs5eUugHtQehBNVm1ZvUjOD
fYZm5t2LcrY9ahaX4L2BuqdU6+e4S92SxFQVVKftAf1fPtnpsdSt5G9i/jCbQO06
8XyI6bbYEc1ap5v9npdHBh8l1+0+u8nGGo7W7nT3FHwTisUWHJK+/LMpmD8tizO5
g8z6aqJ4c+fKgX7ktZuMxoqgzOl2dfp7cNXTLdxX+H7W7vOtkqG8wnrZ5bPA3fFi
43HjroOkYHP6jxu0Vf0afTJVdDtIFfAFYMuh6rRf3IK+/0+8rFwjnbbjrzchN+/F
si3ihwcFq2LbsqP0FiuKNSRIS0lfYs4UkcsQ0jlPKcf44WHMGD8IBtD5eSYoJXnI
40eNFYfwI2ekF6vY/Z9/VntrYsd8y4diffjV1E6W+GXzDPoAFVwy52OzNrUtzuTS
TeUchpe/sixjp3Z4G0ygKW6Wpn217LLKFt36awRdnIRQhvOyfC3ZHcpVzvqm8RMd
VTaWuJzi3Lz16ZNAY3iCpI1MHn5JyN6IbpnCG3r2BWKEGmmQwEZCrTckKXra2RHf
GEPWqvu8qKLCAN+lyAm5BglnISJrVKlRiEsHArjiwQh/RTg2BcjitmnsXgiLGwQ0
PrDZ6JJasQQ8BxvZPzMURLEvBi4+1GbZ8wbkXLPPixhAaHPEdk2zBbzeXUZd5akH
LX8aAbNSrwyxWwHr70cI9UkMq2zRtmSKWsXIc+FbTFk8LJaNkGNXef3L2ZjJsiYX
voGP9rebiqSQ6+5KEGhUN1TqHyFmIXfTBZg9T+uoY6rZ5urpmpqiyVqj8aqaw/ad
KYjtHABwhOYer2Li5BFcASEmyNYT9aqzZGXW2lre9uR9BaryKBCzQFATpvQ4/gYO
HO0GNZRRZDDRGSIus7cGKpDX+Mf9BBHqnrQq9JXQJ9V/M49Df0Q+YeXvV2Hnay+4
2z2igapg6lKdGq/4BFpnkSIBDGe1kfoYAqla7rcPVI1u7yfgL2x37+nhwc5gbUOA
roiqLJCYUdaQ7VFZsbGUL7yNT6VrMlwhMc9A65972KfogqhzulBCIVs7Ryd8CksV
aFreeV5bqtKOOBSP47/FwjDu3OG0ZxbRBPlXHi3dIY9f2S6/07/80QvA8u2qQNc3
9pUnGFdZ1mBe05OmGbFaF3hbmau89503ZGLkbdV1eawqysNy3H7LU4yLDZN6gkKk
iD0ylALo+1w44lCoG38Vsknc7zySm8wIyg+rGX7LeBrIvkrnrAo1msRsot91oGLt
7ajTQX/Wz9sXlScay0B9F8NCRpsWVnm2dlKaqTuiBMOrqWsgIqN7U0ZOw7xns+zX
LP2Hu8YpyNEyeWVmlWMZMUIiYQ/IYHUKB3XmWeeOfFHMliMdU87XvUCy8jJjJIVe
tm+noYmmy/LxDBX9To3gZFkuFfFO9ZF9Ob12pCtxWAtbsTxGjWCvAdoCvwZq5In5
rfLyYxvwtSxvYCQO/g/pkz6D3RWfjKiUIaIiKlKsV4NHJFiyu8e/Vfh+y2kg7P+j
lG5j01IZKQbnlSwuKBWDkw2p9vRFtXnRIfSsNMXji2xOxeOuWKha5mzNDMySGxDF
uBT8OdnKw3otI9QdeHratg5U72rsInIyoGPDJui/b06KHMcGzgh+KwarkdVB2e94
QuD428ftO7M9lQf15dpMdtklkWjip67VO10oEC2lkrLMFTS+I+BoJpT05s9jy5b2
jNknK0Hi6YagTy9MdeXeJp8u0PuypkzNZoiVl9IFqrpERieiKLBYy2xJYLFPkeM5
fnyfjWKlucHax0zmtJIB3owDZDD2164RAHnbAac+UNVIP4AL/dqCArS4bCZXvm7i
ffoSLHNUyqTHN/dM9HwjLLD7vKkBzMoX+HCO8ZCC30lcGjgnJfaxYuHOyp4sa2UU
YNoS+7+SNMg82NMttgmudHavcD4OfnHBvBT4Q37FsCMGzliHHmT3M4RCgzonfqEe
8htEVMgS+5nRs7zOFENic5oTViXkiPJwzc0I5l8M2tjfCP9JDyNGO6gNVB+DSDHv
yhvpSNKcehgILBmxfYNoWpbJMPyCCdhvdKfNgCWXmBM6ICrw/xZCLnY9+6EwwoJ9
7/mr452e6p2TecGSsnqjIW9cO5O2SAEax6COx6ovxGvPDvn0rtelkNPJjhQtXVFL
RvLKGdRMQ1I9ujKvzErGN8kOrSYNxANvE+RuRm9PJ/DOZLytX7U5jkUpVlwAGAym
pvOirJvE9BwljIR9wU8IXJw4Fspb1vNrh6HXhtzG9Y0sNkHS6L0PL4E036x/E1Qg
7e9jp88L8/DdG9i4D+TA1+nmCARPUh+W8HLHEJVxgG8BPT27zxn/ysizGvJvSg0j
tLs5Z5ottdycQMtmB4SigeG9ZAQ5fHGR3xVqBBmO1wV57lficmM9eIpMV4bdwkvL
CRedxytDFswSQN6a/PgelvhNR3tBeLARKRRv75EEKUkzywHwtl0Mjste2Qs9Yi1V
F6Rj+rBYzh0wEIiKU/dxU5F53ahKdnZKeu0LWnSfiS5ENJiVysO55y8zeHcYQfVR
CN8L2rRRNENCrEAl5JtIwgJoasJgZhkUN73DC5uz1sOUKtRov7961tR8bxSd2bmN
Njz6XFsrdLlPtgQl0fxTDKvPrBi2MkGfH8ZbJKGvfJWGW6Ko8NCS9mJxFxQkqtT4
6PuwbcbaZbhC74T2NQ4NplMiG0teE2805tL+1mEEJTi2Nbsvcvg9YB0cUGOHO8dz
KVnLNj/sXhp6EtsEHZeoiR14I+BaXvZvlujhWMP7RuAr2rOrdstAp71oFC66iTq+
kgONcifYpl/ViH3tFPTLKW5GUEfuZKIT/YSrWee6+a1q10qalDO7dZKha6tR9xyt
K+IJk2XC0VndaXCJLLyzmHknx7t5jh+aM+WKX0RT3KZDY2q7yM1TSpVATWLt1daC
lnLgd1AEdLOyKlh/SyoncA==
`pragma protect end_protected
