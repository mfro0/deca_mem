// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gu0Zu7sGsc2EdQY8UDIv/0yPJ8cjihW4ke0jZxg34hqAK8TRZ6TXpRBWGTaycAdMRUcmAMAw9Zzl
AJ69sHt07ZgSlPNj2OpMus7EOF/406/JGOXsVbTf3AebnCRFWsEI1ea13JKSDpEWZo8XukpQtSEc
uHXzVd4eSCxYbVt5N+0BJkfcQzNANYluSXYFW2JvDN6bDVkDplnoN4kqcKjoOS4AwBupmortDAz3
jR0GrayCV5eA9DNBV5ag3iAYNcwqNdzdzKSqMDnpxm9CXLBufU3LmPjsh1ts5hFG9fmnxcj6/4l1
/YoeH+/Yh0OUOmn2gnXGnM2lqjzw6YWRZChJnQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16880)
fMycn6ijXe/sqzQnJEf2HF03PeEd9iQi32mZMvpx+4hAvxTUPKE3gW8ZCJVvgM63R6oBQGQRNK5Y
SyOnAX9vMlA7WwSUo0RIAv1kiS4FsTH+8HLVe3drFpN9xF7MJMIY5vPN6RCL+7ES0ZaEdPio3daE
eviRbKdv6YD5ERUO/Vsflul7Xm1vnE6QQVDjaai0q89Cvqfxjv+S8kSESC5XUV261rILQz0auf6b
zg3SAlfMS7b9pw+RBwKnU5VF+L6gX2gr6A2rlTMYIw+LBJ8zbphL+zMLmp21KO3qW0SdHVodwIJ4
SjgHfy3K6e0jwxh9UAE5YR2U4xWn4tLEd1CXAEpvUGgvGDSvtDF88/X2L0shX3uR4YzGW8iINJzV
RSJkgCxPK4ZbwPB68mwcd2prkbiHXRH1a448NXAWDVy6roMVG/PCmAJrF3nXIesWBJV6hoDrllbj
0gRUUqLS933LAhVnGBZfw7j1DnVosUWiGVEU9WqmbGh1r96esLxDkzh2woHndnWbrbSL+icTr9Kf
/z6xU43hQa7SPBDvHMBu+Y1JGYbzSpcCQ8JeeCSlUTnkR0/EYyuHGhsOEviae1EHv2wJu7NZ2eQt
PmuV/f8JZOCKBWfXDPCIvlGhtePJrFh4+q+vuIjkUK2iWZEmMeWsLbqL1TmCbiA6anPRDJBMOLf+
ImZX0Peuh83Y/oMRWM1PeJfeSJKE6GrHtn4Gq8pJqZoszzZAYiJDG3WqdJ8h6Je1vzn+G0WE3Yp5
WMcTZGk0YL1Mvt9fSWViZ3L0bsDe60QG5M15/YpvFo4rCbB6v1WGFOYkIyZSy/xVPvbeB49jhvEC
Rtiby+jD69HYZv1ZhMkVKsIIQc0ul4XbNmicAQ+lzxqlv68ctgpobb2kNO/TBJq6BioHHIcnQZai
zLiJfMwe5mBEw66ktltEp4aBZvAEIMsGUb6VesdkmDcInWMNaFEwxE+leijopO8kYWQ6FqAmrfpR
2Hl0V7iDd3GApRgnmM1nuArtSzoUiUwFJMyvMFHDPG/hGuwbjr6k/t4FTxN/JcreE0UUFQYSBhaj
xSSpIHsVrVrye2vNITdTA8XbJIKUM6cm6wP89gh3SyeQuMPm/KHzYlcgoWxadkgMeCWER7KonfMF
VckFp5umHWZnLUlVZOlNdU3bpBQe9GBkzYCvOWfsjYIKWA26riPly9nGxv7n95M6P+Sujb6X08er
/1NROLJuI8bMctdkwv1M2s6G2gtQlsPuL5qf+YCcbtf4GSGUDZOtmFUIJeRdDJ0h59TxspAD/wdd
iMRTBmAVfADu1mSKYIq/vg4SLMuufma+mGOl/+JmxmebN/ry9xPOd21Zwk+bCyrTQB0GT/TvUE4t
dgRJ9ewappLYHlTQ03Icc/u1omTxwiF4Dqp0jflC9msiKEs6Fnx2bHXhM0Vr3jm2448t2CMbKgBg
h2TyWHo3opEvHbhkR1Zk0mgggv8ZgQOGypACED0dPlrFe1Eq1CBKpRU+2TdSNyL+294gWP/JiwtE
bIcae1eEQvj+nBXXsC6e+aop2W7BTXGp5G62wkwrxslGNOmSsbfit2ptAvN2UKmSd0JgBwfyvm3F
8QmlxwhBRzML0RqJeBda1/7P/yvXksaKY4aHsHVK68G7D19y39lquDxZZkdLAJO+0MFFoOy27pyy
G2GujP/fAKRCxNI6r2qeGp6DWxxW1vuicy+yoP7C1verNVrLWF0p0SmQwlDI1+j6hVkvFxbStBKC
Tz5se1ShcxuSjf//gioURlMcS2GiFXeQUgSSy2V0woZV6jPFi7I/aDkTiVWf2phgRDS7cwL3Zgfx
z4jSEp81xQn/03Htj2QQ1hhdEX1kwscolnKvA+YkF3kCMN62IzKrYwAXfe9gDndWVLjc4igCqjqz
0oYWVkNFNk5+c/shWS/7dGpqbEbekFX51QAaL1OQzXGVllnXup7R4TDduwWDdmcQ3eznYtRd79zW
/XAHGreqmVxbJm97zgPiiveE40i6TD4RoO7ZMYEu71tyzfykApKTnsi5kEeFQ4Yd5iNvu7UCAhAp
6FGRBf6rkohfW/Ytw+vdERGuReK93/w5SVbbItw804nHPA3v9T9v2jSTSLZH5ges90A9blvgXf9G
5bOifiFboGQH8jzF2aozaa7Yx7N8A66kFn9krMGuI/nia1j9DdzieBxwvaa+ZIZYP2ugVWjXmZhs
L7D5U4uWXMFFf9S+OSmm3D3B/hvt7gTOjgxCbeGfTMIkI2JOGk6DlCg43BZhqZcYhrliMp6GYrx+
TL6reiHESHswJlRTGUjmcXoMVUC7oWOJ3g9ke3P2X/pzNhUyWq1ImqNzPVRVTi1Gvs6D1p7j805h
RnbLLfwfYbCpbYXXYnsFOhkaYQYjqmBQaVUTZZwUoIP2dr0tC0C2ORZSDId+dcBV9Eo3HSBeAg2Y
thayCoLZcIfM5KpG5akEXwysrBSc1wDhbyU95w2HduIg/9cirKCZVrA227ik56XDVU7icQpbaJxc
2fesF9EJMl0uA7wW23UGz5DB1z/0328hFLgca6WgZ5Qge1PxqZ3D6oV3EXR7gcfrjNkaMS4JuKx/
3Gkaxj0k8veiYyhZb+bn1G22lAdQiJ7jyn7ZsgClGjkY1U90ECmKbZIQVkzgppZ1TI1k1gP0vCc+
3qmYpvJgswErawHZYenRUPyUuiDjLngcJHNHtoR+s4qyzLCE4mCbp5LN1uwBsfHtzXWTOZ70jeoQ
8hQRWpigLnb7J9ai9KaFR0diNB/GK3M9uM/1SSITaJH+NkTSnOKXbQoBRCxLXWgE8SYSKVJIjVgP
TRstAUx/GYK+W7KrMV85xpJHQF/sUseQuIWph/srmi0VJPFEglnVxt5k9Kzjm41gXD4VTf75Ek76
FoLXyrOECaIwf9WnAGLJLloYJEoNbGOYli91zHWTnErU8z8tcZwl3V5WifTL1SoCgIjyaBFfcR0q
XapgdDpBzMbgvODb0ijH6IOcy+yNKcdKgW3SMuMa+I7W/NlgeZmCRB362LmHUai7G8fcZ+f4R2n6
0JGnkLBnJX/Uv/YOQcp3zEBdUeNFcn+X3j/IRtyxmrJCr0jFtZagIRzF8wx1PppCXyoo67vUsMIU
QDIMw0y9l8rYqfKpuS3FTHuqBny+LxPnY9BWBDjU5n2x8jCs5NUwz9a79lKeijr3VPa4iMdFkGyq
yqPgiOW2tnUC+4oxCag74Bi8BrCCCkIWPa25td20gVZcoqceaN1FRZ2mWO1BkNuSyUFp3J5TemUr
+sHUF+pz3gHJkXrtLxMeqcF1rRD9POnxpcVDgboxWVPYMw2xmHopqycFuHxyWQjJOTXkknpgnUKS
n48XPRtDsVMfvXbrujG8zLm17ZgQ6nEjy76ujH7+04PqIkNP4GZYuI7dB3yJ8KiyxwmumP6uYfh5
zPr3pnT+PNCh1YvXD5eaL8NRJVlukFmLcsfTF3a6JbXLMr5vvDjY7seCvzBvyVxBjyX2rTRVxR+q
QIxGH1Yz/e/RazLl8cUnhv9jepSatCg9tLbRDFOdpaX2C26bk45VPdJQY5Dix7ZWV7lIAb+SP9KZ
y8pEJGfYXDdB6hTUKIHNjQXwkntRP/nnH51M7h0L9mjXpAKFI5gZVdzPSAAXn1xBtHyO4AnIf0K2
aYAe1pByHqtMngYvzP+G2uTS+EqLZjTQKFSjoehzRR0+3MUHcTxG+52mFpYyEaqVtpdoNV1nkDR5
Uaj2zvopRdB8EyXBy5CsAcyJ17Xrb91+oOlpgbfw/Pgmn6MtdeeDze6aCam2svmAPq8YDmFtKyPX
CPubulhlk71hxPelSSJZKPY0odtsEDE748fyNp49VHuN6E49xhMfXMb2xjxoEqHw3ecwcw5cVjcJ
E2XY7MTDf+ameEZ+B0jt5mj6t4dF1UQZQ8P3H6emEUNs4PnBqxDcJj9A+OQ1R6BrzCQ6oZXb2Fa5
5CJrKJgM8rLe4FknkTCsC+erTbeRqDHT+4aPG7MJHGY5VZU1+PL1eu4WYNAvHbo4TLS6ERQ5trWT
9c+Zr9uwX9lmJ6HBcnqS+hMSMDevjw08VeOCFOq8xLoMgD33hTay8jAAVhZZxtZZ2ZPm2eWPAwak
9mXOtGOznwcLSS7keXoZyCA7WxOscautgu2acT1kKLd5IxW2ELz9gGf2nh3BwNoyvI7ORGCuxYlu
DECuNiYCF2ZGvOhPDSNvSDKhC8M1bFy4UvCmMbRy5clECZEN0fx2fZV9+ABz+SPETVcGVHaQrJCt
K6bD1/+J38XFcs26wbnTisdyaoRQylSYAWoMH6hd9VufIE+pVD0m7PRFJh4rYNLqtozfn32QFdCu
n146QXNhQ93WVlPkePolKgYKKbfEHK704IhLVAbJNyDMXK69cipdtdhN91fq0kOoX3Q29VWDtX4O
w2onOQG0hbkarH0gvGf1uPcWVq/T1YtlS3e7o3EqwCgn88tbTTeLZy1emJK99HIOe+OelKFCLdBm
8ArVK9HSAN1yPizQ9LalkOs6LTu4b9D6YRbrgKkT2HUR4dISsVffL3dpnfxAsFZrAACzvjpTPHDm
fhPToaGHRAzTr2tydEo4jB4p//cJ4vmwSPSoUeqOpCAoYJUddhOq4cFU+a4xmf4klbGn4rXtfirs
sP2Qw25LVVyYm1NORcxPL4pjn7mXLinnD76RqX+Z85a4GB2AN6OE+WPRXTDhn50NnOneTMK4+ZMS
FUIeaw6HRdswAD4aQZBF3PjZalvzoOenp+npgKmKFbyiJ9z8QdOyPH80aGBvO0AB0Iet8l7jyRlU
fgYyB0BlsPoeOGQIteBMakeIERb9Vrb7mLAGMXXRKIoPqrxWWns9UN/xsy07K7NDz9sc1zIIl9vm
L6EALk+jOamp5YgCC7G50oVJZDGx1Oikzjofs7YqRmv9IovK4N1V9kgqM/diMmEbUrvt6N2AqBl3
nhH09LuCCXpnPvwYBwrG9y08ryIAZ6AIFal9ShxqOwyDsqDIA2uXtlrghr0GRCU8JBjOaUZw6jSh
lCUzUU4pEm8WFld4X/RvvTdPB44WE7nkD7qfgaNFGxeOwr4D4z6mVPBuAoYB+3qEB6z4j/YTlfw2
R1YkAjAoEGBncXnJOFDypFFDKKe/OEtv2eGGMqg59ihmnayBGlIAt1rjWy0rHrl2y/C0F2UtCH8F
uQdYwIdM1Iv0KRnP4ihf4TU7PftxSrAaiZSfIANkphS1P+Hfa1yJLLjYwlF4+ei69JCCn9MMgVGj
8b+RIpuBhTLRdqm6xUc4BOWT9rtiC7FOVH6X6nWygZ9qwNqNek4usbq9e+ucqEAOON8u3FTe6syF
cR8tS+BR8jIBuzegwvGcDVbwseEfvYLnU3jjprNJ/BJcloZYIAcMnUtC57HGMBK2YctvqsuZ2I23
YEbTyDmbRqWkk1jFMW6tWlKru0Qzb0zCGA/zDGGZNJqUu8YOOFDj+SYGKk2yfPtpqO2KHzgEJIOm
obi0IEB3ybi4QUIzUT5gjv5mUbx1PJscQsmWOBZfXGP/nRTzYLmZr53Geh5AAIjsDYKhWorFkoFa
EqgTGePyB25GHF6O2BENPkXlcR0U299bCy19x0bJ2BGJPmAPbtKCVE6kSDS1BiwbJvPZeCRD8/jr
XvAZZG0g1uMB+0dpG8gEj+WBa9mTryUOQ/neYP4ogadr7vP8Cy6BA5O+QNCe/XM7UcHhKGYVQsOS
0XzsKqAfer+6/J/yObge+kcI/FvDLpZItmVoyQ+U2WF+IM8poQ2CPx2MSI4owlyTGAwioMzxOCif
TnvSqYE4hWTOkrGEdW4b5jaXxRr0TAhjDtw0+7ubCm25ZX6iNkq9HVEGSqjICS/8PgPLAF1Wat0X
Z4HQMcyR4OHVeKtSWSTkPyZ8QIsE99JaGaKS4NMZpaNGdsKy7VIMMRbX650xDSayQ80pb5Tce+Ck
8YLE07bnqXPgOJj08Xsj7y/CBAv+hYc2DGMJR12NasQdc/dPmcHbyvrykavV7rFedfEBADXgPdex
UwyTWjooLvWmJgV5hRk1ivRSjqpOigyadRwxge4iRhmj7CrHWwhwS/sBDvvnEc2SQ3CbpkS0Mh0W
gRCDrUkTX8x2vFY69quXTnPuihW0iiFg4zMzy4lU4OrJygrbaKTQVleKjeRycjCYTOU/uLbP+pzF
EB2GGR5TNIyhxby2CEF2Q20GGs9UDqKbHyIrIXvsGBt4P5DP6I/8mv7er2cqDABpZ5J3Y1JwxrYg
33tCdwY6HXfL4fWIrYgL5x8+ELIdOMfib30RR4YVneEXPlcBL0tQnu6oVsIomWCdLI0mIk17A5UJ
Bhuc0z+2/1FtPkGX28R3x5yNz0hqKIvHkFAOz12YG3JJ8LyD+oydNjwWHBC5DO+zcfbw2GxUX/2H
sTpK3EE+FbGYjKyAPyrn2xKpPFWgwlu0TpdjLjCabSDyXIU/N6mig4U47umr72otBfB8NsRkmMzk
K+ncF8CbIU1Uo0CpYPXPoV9I4A/jKTNyDtCKhxImtrTfO/DgfHBvIE05UW4qEHZo+mulqrugDwjs
6EYbXhG9J2kuTIddJ8TvXUHhxMa6h10x1AoB18IuRgh5tNAowz2Pw2EtOfRL4j9j/MuS9sPz12Nb
IiBVKozOHfu6+hDXoRFqGvw+1syAimUCHAZIxLs1KJauNbZgV5TNnN5xGKl6O2+vD9Z1CynE3KmB
udXed+XMhE3A2jGWcBDvCvYTJhlcKUePG+2sgOEh1NuDz4zcp1kn+jljoROrr21ReMFqT66hIxMz
nQPgJnIl//qBg6tuk6SKzQ0GJCIOunVEenwZP36Fq3LS3/IQ5Vra/ExoJ2at3G0cslP5fjtGMoVs
lj0dyZvMICfFLuK1kXZlCK26JESKScSg5i2ZYYQEjczxy7LVNY66UpXnefGDhN64nod5SCgQVrZ+
AYbgudqD+VeqLCmKjHYbx8aoSUkmqA2Njd+Xxfq7iG4PUpTSgf/CqHHdK/w9plXjXOQL7czjbN3Y
momA/OiSHQA8mzf5JmoIUucT2ZAOr9k7ebRGKrblKoWqatxxmQkbjruIeJcd8gyC/jhKTdbjmi4V
gCDv7VcPTk0IV4HeIbJO+0JRlxOqmULTswfeITbg5EWmQ5rnKg5sOo1M9YEV8ed4pcDnuf2MM/MJ
st4yupZzWIxM8OIy+vA75zdzxJs4bOmfOulUDwC519Mud5s5Rf2h+d8n7ewn78eG1exY113QKhnR
b2B6neMcov/B0l5X4pSnR0SD+bIXOrGh/f5rLGFrgwLd7jEUpJr0UgNR2KrrxXjTcKs7pwTYSsLL
lIi4kQiQFwkOIxAG/6jGFjUgvHfl/jRkToI+bXlXdfFuT5ZWv7sIxOZFj93IGNvA4WZ20fPmPt2U
kd2jSBUkthnWhd+ndAJ9s2xxar5Qe6lxi2bJLWZxQrAiUhStfTkH8PFPpRz9RJAkbg6LTzQsjAXS
xp3TDmbB/QWDdqYfzJcYW5fMW11lePjLEfhaBagX1rDSzPdy/ifF4hLNmsekJzqr2QeFo03N7pek
u8WThRHqjdmZkytzhwkYfoJhO+OkhE+ukyCAA7rO8eiX7swTWDPcymQ5E/gBxH0St4DpvFajPDrH
Ik5TJKY4EZlz5Gp2kjVYDm+42rwuQhac6T72mCQucZiYnNNY6XG8s2U+hYg71WDBmIUk5XKUHVpG
NIikXqrqDEG0DoicVilCn43ulJEb+dVL++nPEknYEthv5kG8EcTVBfS6GUJJniQsaEvN2WYxdbIf
Cp42amwo7KW3AggBg/PDCXLOecl/WOb3C4gGTTwBvKH7+XYXoGqb3E8UYkCGbQDFQ3o6JkgtcsMn
JHw0XgsaRU2XJmVw+ahMAk99hQvzn00JbeuQgteY5UnlSs/gfhW6MPCDL3267e4/S6Wl6+Gob4ma
ECr88mMfJSOQ+0vX6E/l58RcJq/PfUEFwFHLAh7azOL4xSSZ0hNp1JyrfO61bUgMeWUFzi7d2YOl
slPRDskmzQ6gdy4mvd3DCivU88uoHZLOYw+u5JT89m3pV2N4mtuQ4oi0G5E7L0PJ/XCrKXm3qMsa
GaigDzMk4iRn8adXWj30RFHlDs0YkKTvEgURIF96gBwTeeeUZbvmQJcdixaYdnPQi5DoEVlYhGbS
EmDjsGZ5QrNKxGYgGTzV4ETlKC7j4SQHKAOa6Xru8P3X6/au9qPzjOMffuJkYTgUpdAHamTR+XDP
agy1k8U7v+oQgs1Jyc2jGmYbTI6j+gXXQme3ZfvDneRUqjaRsDtS0Tq7vtwzkbtvk67TEkhLB66+
L2wRUQy62UL9udVHvcpwrlwNScDwJCqoXKLtuSkH1W0egpP5lDObtGW/fr2HrvlDGphK9oLVSXh1
K8mSXoy0hZK8cNEmXqYgk6upNtO9YPDxOVGwNVA9YlqCFF7xijywP+3XzXMw8kMXWvdli77cBrUT
Zgd8KXeoBQhgaPpTpy3rHuhlWjD3KXZLWeeTpgS7n08/qF8QorLHdBtxEs89NHTZ1gzkt+21Lueh
KuAtRyVn6pshmwVHcn5L9KunW5JJ7Fz8TfDKzRtJa+46ZQ+2QSPYCV8vCjtx0+Wb64kp/b5lHC+5
Psz41bSAVhbWt4nUvSARE4mpnr9fZ4p9WBgJnrxqgnwBBOCOXdzadVOCgGC3ch8XuLHO/rACdpdW
GpmmXixxDsTbp1OM4HJjBgrqeIMwiwV6yBYIXRWq0yD1PwEz7S9KXsQ03DnvqmAjLxi2IJi08SOB
t4JOLNHZfhu6R38d1SvzuRo5PtyHn7Yuzn6vdZ+fmUKBYv1erfws7SHnl/w7YeHKcnffkK0eQALC
XfdF0aEgvfqy/X6oLZO2zv3JZKuieluV213Q+nJffVy1mmROQtkLaia15KGS6k1Wx4QHkwai0Dzf
iH6H6GmZuN9NMcq/C2ls/2fH+7NPtZBBNWnp/8QIjC2mUDiJP8QNR4shcdWNyM4/bH4VLwwTYX9A
c6Z3jE7Cm/pmeHD+NTAvMpw6+6zCViwxA6ClKFFPluERV7g8Ku0o+boKe7EhQmO1NHsGO9Y9WdKZ
f4il2kCDsPDP6DOd2l1uD6dBlQrvIZuRdGUTDFj+KBJoSCukCvFXkwxU1QbsGT55XifBAEZ+6SKD
fkiZ0/052FyQn8PC6Mdw+7naTByY5eTHEoby/8T8UxPDR46LoJNu5YTZxP1OfLeTWBwsqqdyLkpd
m4PLT3i8ZMCqeZE1WGN+elIbCLfd3MQ4oeD1HqvBlpNcswT5teOSEZgSbpssv/7tM57ny4PeKcT2
CA/Mg6SuRBOPbiGpWFHsVqoe59TvK496qs4G/pSlY+2OJ6Xu5HH4Qa8FInrko8BwTZ/AoKY76hSt
rEsDGDJHXkljPkbRVGx0QxKeYCqD95OZCK6pJQZhHCoLkmd340uD+F6YMUchTq1FpDNriA1sboEs
jUxBGDXa/dBVtks8SGclwPN7A6PnSa4swLhqvtPFx4/DO+3QTwKO1A408tEahO6ltMWy++Kzp4fG
tcFY9GwqhL9QzmP6ebBDUUUu9SIQMa9qe+M12L8xLs8U/CO3/SxKYjF0QLuEBuVAbbjejB9JKmSQ
FEyZ1Xf8VPzT9DAQZ5YXa5S9jRh8eLNilZbnevPLBjMPRPQ/wQlnLVNNPnm+MC/jPdwW0IvRYZYr
X2/H81r8J+OffWiFt6fz4E2v5e8vKYYhGCuQ8ggzLT4TOZlRGpzSV5kfamlXTC+jhurPN8v6xNBc
tGfndr1zXSepAsG4Gu8ngJXuYJPpt5K6JkAAuUyvRJVbjv1MUHxmh9dGVoP4Q6iMevOkYPZ4zRWo
G9BAr3f2gh7Gv1TiTudExhskL+grGwrQAPn9GjHfsWWU48ffe5B0gEexYbu0PyE7xVzJSovhrvac
Cc0GvPbF2r+4XJVNGb+XKNVp6ziOsLNHZibVcrA7oGMekbvxy80VN+R4biJrmwEfSZlU+NUgybDg
yJxaS6Y/ZwIT8J70b9vDs9XE3y3wF90b3///onTVQEZDq8pCv1WZvr+jYY3kk3DMGPGwiT+lW1px
iB8eNvlkD7PhtEGZkYUFgMl5H/JPB40pnx3HFmZpK1/P2UouiezfmJHQ7o1C5kZyQRuDuhB0JAO/
WWGF3Lq9BDjgX41nWFO/0h6NAdhiUWsDVAXNCIzLmzle6g9fUkOakk7fvW5WwtxMdqJeo2kJjJzm
MabkehBDX+ePDGMe6VPFZBY96iQpfd0l+ITNu2W7DMeUAbSEtr/wgucDwLLiTb3ZcgL6HYtLmPV9
fzC2UlmLBzv9ecQb8JQlaHpwTGuAqdJgg8DUjT51Uw7JNGafJ+8QlItAxKtmSnZkn7GEK94ggcKh
3r+Dde8J1Fwpa51oS9Lr3pKGROZ5osq6zSxNue9yYijN3MVnnonaf0H0V4jFx1N/gSD3fQUf4oXP
SJAcZh4uKdazGCj1S4j2vf7u4yYY0G+wqJaVcC5s3OSWgto3n94DEOo07rt4yggtAT9EI5OBceiQ
tMQkUXupozwim9i40ypHpNIFKoj4M3Xx+75AlSRW2fW0PJhJJCDg7NctxRtPRrSTqJ4jAyxc4LmK
csjL6c++MYd6E0W4xkPjDkCBhr5AbiSsLd+59wE1wNFNbcHyWMGySIdvZzR8gnVcWbpC47fV8h2E
tr/s82F6ITns4FWW338XNqiJOTb9tJQPB7Lo3Gf8vEpwMM0Qg20gxopEY9PZHBnz8SdskmwKmrPN
7ry+hKcG191msvPvLuOMfXC4acQffpCqr3kjeJLOzxJex8FK/Fkots8c62mF+y+vMgWUM6Xq+7pI
Irh01elBP184VnvsQjcYVo30PQ3IiY8LhRlovWnJBW0T5J420ckbmre6ZNPK6IkEr8NRWNEoIhY0
V0/BchR/B9kM5JA22AHyZJ2rEpWv3fsx3oDQbMfzqMfsP4LZHZl7BQlCTPLfEjFfXsQdxnra92uY
1ukW/H4MPPmUusoq6lnMlNJicU13AMfbAPK5vS1Cat38gAukhhZIXtsivJJ5QaaeGZVbrNiyJb5S
9TC7G1fQAsDBsueBKj0kL5oHYQNHUmngvXzsZmxqPuUDyCkGZRyD6G6R9PKSR4WcRwTrhMfDbNQY
LJEKYeqzHr4JyQehtatgMe5VGrbfzd7HinGAG6S/mNJZgmQIgSAf6CoCk5zvI2gpfx+9iAeP+St2
Vv1ykYSXmwM+vprZPdoZ7vOHJ1EvB+AT6edtVLpA6GXQBgcwYzT3P6Oi7yRhFzRe4zhll6PN+J/T
bfHv5ICRX55kqEjpaILvdWkrUiWraH0KtGB3Tq7rhxiGaiBEqmlW8XeO6pEuhbjmzejTGxILmxuo
Dk5iwbW7o+b8u6aSE5vF5mT9iaIBzQBDsireSpLbwu8cs+pN9kT70WmaaHInr/mZm8MLHwFW/xEn
jQCTZHhyHUT/ZZdQwiQQEfNcIXRizceCDF3sD5N1iW3Mm7wK6J0LXvY3Kcr4FtO3ywPmWhbxUTBk
yPZ+rf77omkzaY2sHfN17eWVg52hrfyiYhbuEkhf8b4vKmZtFE2l4ZnvF+yOnrp2YzS2Zn8GK0YP
rbxcRqMcgr4jToshyDYLRqFbrgV0BU0R4pRAkI2MRkWFoFPt+m+1XR4p0T7BQ9nZ/Hdwq5KpiWsF
WPU0+3wwa022S5O9UMTbt614kjdr3PXVJUUCAxqOcyMc9crJf2Hm4f6QZV3bO4H5wtYEwg67WgjO
8eJQEOQMrXgAP6yt7xGa/QinNUtARxya9wBkr1V/3sQltj1FjXLgYhUIV193Ak7ikzqK2talOuQz
zRYzavcqh4lacYqepWIFZpHjgT4RIu675vv/iFQ4FXeVApzu3xkTqEkynkpeRQqWQgbjzWneVG/y
EmMOLIKfi2Usl08teJ0xtBNgmg/DZc1j09pCEdN96AzKarvTPoStrYEVy2ZlfMP8y6ZTyh8+vOc+
pVe1EKAnh5sY45VXusCEu7xxYfSAnpZMX0YmZjzIWFDyIQXIwcK80CuHh1k+qkgDliKVkgoPb0Y6
d+nuz/FJHW1JzYUq5toNVBl6ecpSOWO9V+U5oimKEcmTPJDno1/UxuTFHUNjfYphmiWL99z2QheL
Hczg0IJkbUxVgP5V5DNgyTxG6+41iWsHxYC6lEmuLH2P8KmU4cEHOdbwKdZtPI2UDBnEWYW+vNHE
b0fuvs9drqPCOjiptWpk77KP5yUWpzSfmXzZl8CCNY3AOuOU2+bJOZlJGBEOQJHV5VV36+JFB8al
muTWS6mU7G72p+Q99JWSAPwh7pE5tnMSD+MqScPZhdTCMR/3Kw1aZSoJst2k5QirmDZaCKkmxTpg
l2ua/89CZWR5McTkLbmWw9wnhrmhB98Sh32DnfMEYLz9pg6mcZWxf9Q1sd7Sumfe+oDMi+ENFtwV
0MmNBMtIXEZSjYHtLIMg2usQxb8q8osHGTU8B6lQroJl5glye0Nxzr0vxTzTci2ZSc2meez2GX5d
8xrzu7OXsyjo0DGNxMp6hJ81tYrh9h43zS9e4vTZDX1jgZx4qGbtUQTpO3DfiBjhnZusfopYESKU
YCVIGtTv8V+Hryc1mQiYbKI+b8ClWDfhoSBgVOKoCuw+1OI1hFiGNVY7/2+RLmjZ19Skra3U2fhf
wyQfXPWQ9O0YlsAwb3mDddjnYfXxrcZ5BUcYWO9NxjvPxPwBytNhpvTBygkOi7XzzieAH6Ey5vIW
bDnWfq9LLdKFCN5IdF7OFWwumq49/CG5Lg/CliNloG0y/IBIbTLbHJcmdRf3o5MB0BTiLeOUqHZw
gqJv5pPGGK0cuVtmrKQ15OrYgeW7cu6QfSXwyrBPguFU/jVEEn2wttoIOymI8A5K1H5YObVZprD8
WDwPTmpT5+Cp5C5VMLSI64SqdNZS2cRGQUnUSs5/TTfQLkL3l4mA5CNJJ7PTdnYNX2L7Ni2Jk5R9
8iPU3UltQ/FioJq+2I1luC48je2v1xxTnu0FU4QCmz9YocrqCkYn1lW0PNT04H7zb6ljCtdPPurM
BfUlptxAlYCE+Dknskl10peR8jHiNRkKb0R5EiDHzypCyH31LTg0PcQZLbLxEf/mXeO9eHx6UMGx
P8uCxLWcCzioCHIEoeH50j/3RmMDa7trwsNcF9+qGNm+B5tq1c4ZD+dtKE2+q7Q1bUs4gUdKpHZ6
VI/gM9y5Jl5Lxq5e9kw9WN3ohsuq3nlgtpWBqwNeaUhGNceuurt/coTwUtawq0J6CgOKi2NxjyqB
io3BCSGHq/pj3YRPI2zTHNiOBOXBF7bzxXxru5mEa5RiKL7V6zI6am1yRIT+PEQI9kiNKClV0iBL
SD/JecSvtUAWKJsqEYZ19Bk2oYh3dI3nTPUh8w7TClxZZs2/Wa4SWDxk6JAn8ZezLJQWLv8FHU3X
H74FJ7uPPo4JuAB2/4z7rSkCeRh59LIekEg08ugZOExQTNGNqSAVtL+7qBCfDPMuhhxMp/eTv/1N
w38FXDcEmGCpWxwWs1pFqUuIqr4sla7bcF8BTijHb7nD1g3V9pAoTDb5jXIEXdcIrtwJtkkqMfpO
PAaUk3EuZEqo9iuMEzf8RT2nAuhywweiQcDEalekDj4R+owHgJO+uB/KvIC7d35grAPKQUMgG+iI
oYkRTfykMf3yZkZEmVflMu7f19s/CAnfQXCah9LezvbmRvAVOE58wvbqpZedEspshoFOCSTTJngL
XLQ8xolKw8CrxnvtbX7QcbyuMKRK1Y4HItb3JPUWLn1pOmGUM8Y467hRyZTqz8ocfn6CSGQ1tP3Z
LZ2a2HeJ/eAT/w7OoXrnziECExohO2uRouFQArWxyBcTFUQNRetvnKBKDqH7hlbSzGatxVRoUbZ3
Ep63I0s2X2me7jaabVeAzIkJFykAVvtFlO1PuzMSSV02d5tj4h8tHfYuHWnhPHHWif/9t4lT+9p1
LbkHE90rNFU9/aKJdV6IfLzxGOCN+7LqZoClaNga9sk8m025am8YtIz6S7GL6fedefT/1kPxnyVY
fasOJ9E0UbcvkGtu8nZ6QwkQonQ9RHJt9E8euNdGSq1LMnqIxh6s/fJInlSRwCabn+y0VcTpD8NG
9QJFAY9m1mf+3SWbq0SZQygXj65In1FqtYQygWWfcWLPbCDXRsry0BHykMp+slp2WEHymKnlCdkZ
iSj0EcFqR7FQfInh4unW1mjh7d0yCyjGBrVpUGciyZHtSU0jEFJC7tu3+mWOvaOEAbUHKabdMIO0
9Z3jXsGxEb50U9KsicvXDpu6NjHZGKX9XsfYI50NDYCWPnsH2Nx179smkIk6xS85H3MYIzNBqvyS
S8EgHPPcp40uYgNGkjJN+6VZlBN+Id+Bpx+n/2OZysXQRzECUNRekXnaLtrAb3d2d6GhVh9Jgcl+
VAxV9X8D1fb2Fn2/1GCBCULzuJLPecA7qw0nR7Md9sIiPO8XTUY7+ZCPI4s1ga6l4yYAuvD5jqIr
TcQjaNdoMv8nGdu49djT27fEY5Op87UmJ1nZRl6bGrVGnyT0ZNBVcZS7w6p/xLXmYXLkMfERnFK1
CvA8Lqob3NEFjIzdBgcvw3BOS4l7C3d6xwI2Sr1VycWtiOvEXBTk6mQW10Di9p3+4z0y3yXRnKXC
Z3kqdtyIME5qO/kokdcKwp5gNmaZO2w8r8D565QCs2qPa4RF/2Qclzg2wt/idU41WK8vyJgheKKk
X1tQz8KRtWeRC3Rwkzt8kr2xxDwsU/R7ZHYNY1vVxkfpkXEOSwpvZcx0p3zP+sUdEEfPqTzNG1F9
xGvJRWxqqPykQNXS1WulzYLKcyvfduc4z9Uchlu93jSv6+M9VPppCpEwtzE6yvLax1GoXxHG72HY
3efR6pxytNXHCDWe2kKFTxL73K1VXHbl9coZMu7J2aSoq42yq1eFjix6TA6GRQ1YoX0mSrUJQRQd
9L7i0nu21iSP0tqLY4S713xD+q4Un0j500OF1tQR/PxOvLV/7Gw3lSt6CWnaxasgP5ucG/SBXm3P
iPrP75+H2GYu7B3khKWH3h7UH2uSm6WcJSgsUBZGg57195ZQCV22exWOgz4hw38jJyWYahB8Pmsm
J0RAi5Bm2QRFVk1rVZA58tSUGKDG1jkz9xgJXEwy3OA3Cu/Hhcz7MmGgKkQf5FOIsQ9Qn28BVvMI
/dbDYunPLOCvO/Y8lLHxRWarwDvelcPtuKLIxm7u7ijTPk0zK+AcOttOt9Nxm3T8vWNbAjkTnB5+
IBCPxUBjO/ON4lkDI1NTicRMZ5KNJJ0Q4PVhvYaTqHFbcxSv+nHlVHlosKm8uQ8T9iaLxJu13aMd
3JHkQrEI26aKo2pnvpgBW0PC4B8Oi5SdVNEmbfZa2UXAGrH51PKRi/qvXKscljpwc3QnEZvAqcaV
9tHY4ZdkrWegauxaeRz1TyZ7SoAgRf2iCGr69WGBtgG0uaq6nmbdp1hLIrdSvFUHnncsrZtfpgTQ
YpkjFmwBw0yPQ160Gok9KmsuJDW0wniNZQ8HDqHbkMV8IyoPH5f5Sl0UgUiraoXMhef2x2tNxzQx
oI86j8cmiQBZmoTL4SmvdZtBW6eSCW2K4JERvACbaH5B+5HnL/4JdTEYpveXf0rrTU9Wwp1ZZSYC
6yti8Bq5NEbDyBT/Shjiqha0sTZ/JQJHCtsPYEnmJIYsgyvxz6Xo2OCMtZ71VrqLu9t+Aty7p0Ob
MYzoyLcEzx+2fu9JqvFd5BeUBNO5bLjZifAxjz9KhbIW9eptmWGD1tiAuNJKD3CD7uNQad9PHAfS
uNov7+ENR/EK6cgnS+KNH955A2fR7xtuWgzZU1uSo14oikyHRSNvNMfYMDy60iq2KdHXHtyNd9dA
wa4BSZvI1FZn9G/Mct0r3ZArsEsBsna6sL8m8hENcK/PQMChizJbmaVozAElTVkHR3wHGdqA0pJN
ZfDUsXIr4Gg+wJF32wi/yNd0XHckk/+vgOGmgCc/hCldT/rJANQNFhrPBVoi/7XBLq7XnyrIYkwk
tSKwRS9gYSqxpTs76F7W6GkW+E9EVEZk9plJDtCnvChcxYN5iQi5dC/CuhIda4gQLHmk7h6Ejgko
Imk69i2PKheeLlfACv138DS6mbV4uLCWjVBdxYfIzQx4r1tcCMna88p4R38PW0VcHKBRiQKg0dpr
268TkF6kykrWF9mo6zurNrNoILTEkLsUGy0ppDSGrqw/kddl2LYxm5PkkFWdiZxbRfgsdx+SrqgF
L1EUASVdn04v1jLCJJpnofAEr59IDULEMBa9aF26K7dSMo0OUJ6B1vigCM6J50UStwS0XU5cXaWW
h8jNhemmQkTCB1dwlum9dYNYP53W0VPny1GlH3KHWm9y00sXLU2iG2T6/GpX6U4jHAhdMsd9vy8+
zuxDr5ij6y/4HjxpIs6KHluSLW1rb9xZIQJl5npHJ0Do16q51rdv9hmfXjTrf8YDMY08sCtnGP9W
KCxgSzjbBQTqxVh3pnkf4fxosdP/YPAaoHmNtCNGuo3vYz3iIrpzopJiMsaMiL4u2A0selq1/+QR
sDBPCCLeocsJh6CfeMG4dsPs6brVzQAfVRVio3TQRIEDVgHk9+fotIR4jaX17R5HL2mnWQpbMBxT
FG3x5rvqsban+hHuny+kvbfKKvMgm6hsJb87DzqmdN/T9iYU0pLUE1VCtRus+27iP+yv2L4N58NV
g3dLJF9LVl8kmy2fwHY3CknjynX6VZjRiXjwHQ6Aj0c0Z4cXjMfibeR9XjQ6Cdz0JjypTOKBBR5+
J8Av84cKRVUSXrrk/sOvC9Vy2EI7wXpLPltq0ei/XZg6Lw6r79V5IDpl5jvcZ95Bnk2MQmJLwtEt
w/JUqFvy3tLpWeZpBzL4ArGpI0tgzxSG+NfJm+30fjRTwKBeTPuqDwqnSxZInZ/zk9f6pVS+tdxI
qoUBcD7l3ctekJyhjbsZqol4D/xC0Ymkm66d+fe2bPgGvEsducb2ZhY9nBYKFXUmEM9F5p+2GXtr
fNdROHmzpTk1AT0dLOs9l2/ANki3UNMZF9Amd7NR4CRtKEdrET91nKqnkv/AA4uCwzWQLPClBsnK
AosZszDDN5iyrQYmeGs4ueO4U2ndqStFRLu88G0xHPsvXfGKilo6yGYMtYFleyE78RirtDPtRsTo
Od82Oy84wXSJq6ZQ6fGpyAzuEdYCIydI5NT7xws3f9egp0AgrvDnUZWaXwx7rtBx/ADQEa5udbG2
SPI93jo7jp2yu5CUT84vuQ3Uff93vrjNe15s3DSPSkVlJufcoTuErwGjh2Y8cWe2LDVD07qrLZjd
OHaimgTzDfKCOZjOsOig1mlA2I+FQR+jzuWh1/Je9OZ79XgH6LIPqyjzOKJ8ny/Qdf3mBMGMnUO1
XuTJDlCUnyViVLIsJ+r1MiUhkbI6d/HD56Sil7tN5V/5QrozLEf1TAk5GlJqW98PDJHh7b9Hk33Y
O2NIqb883/Gpx48WtzmXX/2O2M4hP3L2AY28uQH0mBxFl/KUtmcPkrsfK2bTG/1dHQIPGPf+3/Vs
gfvfW7djB6u1rzXhHejpw7MJlh2TPgRN2frk22R5qRYPC3zniZrvPRB8GRZKS2mrC/8jab0qodji
xLmAaOanv4Qu+Yb57jPEjYYCBzK+tWGEZr1emlV3NezWAPBlcHK5oy5Y+P5yJ9QhU2/J1jO8sLa/
GF3UpvAKiJv7FeZ6UQSDqFfW6yiVnokHiECPEysNWbhCo4AhMZuBD8nHaHDZT7qpeVDX7/Itg0C3
GRiXo1QOMoU7UuQTvUVsdnuZwvJ0cUoVcu5cFiY+T4QK5knb+WWjE9wwzdLrkMUtCprjsvGOUIFR
o3kofhcoWf9AWxslONkK0YW0+OcwVVyIO3P4YxsmX/y7iF0R3Qyhd54eVwk7Q1e1HMTghuKnl3vd
2vRiNgxi8ssIPFmvwhSSnkbtGKQ8R0O/XhQZThM4JFTzeYR5ngnSChUUwkSGJ3+/m6DKxNGxUw39
xcgtAtVSPepSvybIZCkJBLAtScMR8hXDuAWbArTCd8kwsnVj+QlG1rye5qVFbc3a9PeGZr1gARqc
s+4Io6smIIQT8k5MQQSOFYItSK5C4+fwDq1CDmIq4SgUfIptvKfd1HTX1xhB0L6UodTWaIWEXOOO
a5rVjdeE8NEZFmQVT15kXWGBw16FPSyoA8EUxHZbJs1IYOIwkUcl44/9C78cJJjLwmfPP42Rtk1V
9aQlz1EqosSjzEYDzidOCpZ1mJc18WCf3qMv2CtAISTyPkKs3A4oIjq96okOd3EdBFs9+QYB6yai
I8EIwtXe10Wz5vf1CYTZW5LcU12EKcS7WjMGBvQFVt0wxl01BHPHUi5JbbW4tI9v3xk7L18fpcGS
No7FhkyaZNG7LKkEwgipjuDFV01krQwJIeTVgpoknRYsIl3imheOZiZQarK+oHd/ID/eXqdNn+an
4DaFAB8XMky8vNVMUwIVw01sthJLFg4jNe/OWj3p0xWXQzqf4kXjns9bBlULl8gR6yB0PZdHRcox
MF0dnbHmXcOj0SZnv1sAyQmDXUPiz9ZOuasVSaySCunFBCggMjSC7iVhfVHdw9fbDH5q4EI+RNXF
26HLHnlVStjm7JdOJOpQYU8tYnkyD0QqDnkeujeClhspwfh5bEhqfpU3hDwN0e82BTTS7GDGgdHd
abRNO6HBvmQYEyC8aeBt4BcBwMqvlxvQdevF0WeB8YTI2DvrTFoF4lwoA4aI6rah7ZadHsbo29BM
+5d+fEUTru2KgkeO/MFj4pw5zej23KP/bdMdnNppih/UPhfZQ/ZjH7MIA2WSqemnDD+h9TAepnxA
APOvC1d5rCTlxCtS9f33VgWGYub+JpzQGzVaKxkviqB5X/QiGX8PwM5EeyAWbbls5xYX+cM6fP02
ZHcHiVUv4Xi3jKN3u1t4cdrJLqmR64heXpbcKbCYUOm8zSAWcfNgAuWdwbIR6WvXvF1qwOVR1Iva
rlfXQbzpJq0wyHwR/Vlz4mrS9PiuVhJnHpAQxA6QpHxFk7n1udWBkXS7O8sYoeyf/biw8AGE3ljb
n/1TzOhDHyp1Ry3xP9nerGTPmdNYCT2r7WtRgKyoxSd/lzx6r4W4FdiER2mDxnvBVafxUJAPrpT/
QwR4acEPh+4A/b2Wh7NCmyPBdD1ThKyOwv22T/Iwx14VqpSNQB0YHAAXdS3BmQ6LJJ4e9aznXWBb
3eNdKgbIfyzdx6D57pC/CwPyhBpWnKmjnBqTeosKvIYIlLD/jaZBbw1p2GyuxweP6F3VXooP4kgd
B7h5OlKynnRgJqWd4uVNIzZ/movKQo3wSa8VkDKgjjWRcRZ8bxCCk6+ktkBR107eDiNNUT7H5A0o
o7Xp1NAK7CAlXjEbP0ZmASJppg9gtabU6/ar7kA7xUdEA6i12Wkms7A+WmP2ssfRZgSyH8Yf+thf
IXiUFtCuNCmxSAGxOHwvxf1l95YcuzXn5NPyoh4/OnAiW263uZrcQjYMnvOj5QGLljiKbT9aEigz
9Wu5RLK4LY6Zv1UbBN6pUX/msvNRoUs8kydqwHRNHMga1hCV8ERdXH+tGLSqYn7rsXLavFKbWtmK
9K38XAj9uZhIFCG9e8VilIZjXHmOMN+/OfkVaw5ISMpjv/o3OaTOExe1wJlxNBR3rwniGBWYoMud
LuJBq6DC+egumoKEcKZ2AIKaohcHkliSggvwxHRY5VWc34hGRxxWs8ed6jU6QOcrrR8ompyvc7Qw
V356CYlogaIpCi3sbH/mJMR2NQRQT4mOB4eyACXdCKZ7qAGRPx9/ugDKw618YsdZktZBayaT7bEX
XHsY26BQFxS6BI17c8/8oZQbSUYSmeUkJltaj/qXelhOaT/B3jlo0JlEphfG0fBEEPu/GsQPlt3G
kAqV4eOnrcfipl4EM98gQADKGpDtXv1x/U1UNfW53qtc8eLjxKHmr8Jr96hOJ87sFhDNrBVfJFQD
94Y125OuLhLlSv5W+65su7CJpxZJdDz9Sx4/guL3RJNYXQBxwY3TJGlxwCHZkTW5bkuTJIw2dbxT
8lNr+QqM0eVo/UyVPakpWFm8fbkq41qcOpIYxlppaO/Yzp7hStNtgBh2mdu4iTfUX00BfAesskD3
x3svF2ITYuxHYC6wb4hkyWbkLhSPIsuJMKwt7DE/4/f4EzkALzZL2LI5jK4eCwdwp1maNRcI/gkL
9bFOv1zo3j2QF0zF/wYpX5349D+Fogfud/1hF+dIxaZyZJjUowQKtfHJz2lcU3eZ8qghIT92KDUV
KiOlwdC7P7nnu0hIUMhcM/oEMrIfzo1NztIZuR5aszSLjg6k0kR1XixSBilcERp2stSoqEGLPQoE
qoKgB/VpxSRIyepwJQXoMrIVNLk7jqefHETyB3gtnRFP0bRQbgwwWybZzMMklPX+/Ap6XvsVucnw
FEyPWlU3XURStc9rj8gdrkI8RrXzNqkBgdWYdGPFzUUqDHMD5Y91DZgJ9YJb3mqt23JnwEldf4GL
TLthcacDX2KF1FdoRkFegX0Emdh6OXeaVQ79/OPlHlJfW9GhpkITyunDNmxpBd0N4ZATwcU16CJC
9gk9sQu4WeU8K0jUAkmxE4J1H5HPc58taV3SFrf/GouSBhKlxyAloS3L16aJIqAy1AwrAV/2sRog
FcL1LWnGxEyhTnz01kuVVqlKEpZM99No7YBvunA3mASILGz/M9llbk+1lLdBHlabh+BPsLByBRQU
eT2BWm9TbooPLkG02XeC/P1ou35wGYmwCCBzCVaD1BzNevdtPxMTabmAbgVB3XMfS450qNJupRBP
N0W3ZhrOOmRtgriEIjXnNougCPvGxno7EgqLAyuvh0hsxf8pJZmwmcs7iF44YnY2Fcq2iP5CeNYb
CWlAOl0kq3NbXM2+mUe7NPUkl3U9Ftb4m/Eot8PT+oxz0os+aj9A09eqN1bm4wZiFc5p3TnZIYPm
lq8jeX0rTEHhQFHHpDd0Upok5xTD2CXB7S18aTpazgqdYeiMp8JAfkIPpvY+6Mjqw9tjdZEQYsSH
MHukFjKfsVwp7jCxsY33DXxVk9qk1so9bONAxRtRvYXRbWR/7SthYTdYJfs3pjhU5iaS+ySTC3de
8Bn8n/UIAGtlsKHlIkT9W4IoCKghB8MTMltLOSobBOyuNPCcy3ibKN3G1U/N6VX5nQCIjFxrQJ6+
obPDd8QaTgv+kMsxQ4XrqpIb/B36pe5RjboDfZXSbY9eeCRvIl+TWGtw7CNk4Ma+BL84ROzZOgy8
6h7F+e5/xEhkVnETK8l/0HXfz5ul9DdspO04DYr2Njyux03aH2Sj5X/zJ6gp0eL+bxfWw8oHXFFQ
P4DvyD8rvquZmp4ZMedlhgw5BQbPTFuuGItU8zXaaGjbXvvGi2ku4Z1dCTyMHLNAKceFEa7CC/CX
ckZR93joGvUJ820FlVEo47goUxHr450vEIrwj+RLxvNy1L3Ac2hmQ/q2VBXgzqhj0C/f8BEr/U45
nbH/bVha/eJeJAkERt52YWGQkOlWgfUE0on8dSVVbM/UfCQ6az9drsdcf1Tx2/KwoON847bBDOwS
O/TeMRHPdNESJ/6N1kGoEtl9ryHdxqpnSF0B6yxX6mwgRwIAToza7z7hFUPflU7tv3gFuzr+C6Pt
M0VmfIgSk4ahz+oFFoztFFG/Z/k604HchgPjktVoYFlGJuswiyaCg67AscGie+t+/jmFlfMJ1dTt
OpNARgkNTqfgojwZa72fpyTXv90xvbgYrzJ6DISLpag+9/if6ehIDNE1BD2fd897PNLrN9MHjI4j
5GgLLLQ0z1hlEikR1SqfC9WmnC+aSY+vG3HyZxST0a+12HBy/n1b8KRdX35Mhd+rS4na+V8abg5i
o/oWhMjFQQDLySHt5hScJK4WmU1etpYvPDWxuGf+bCf5vm1UF1fqkPsQXLXTfNG3JN/MPdv1eSRP
62p00OZXRSE6pKVHMmKCzHw5V1pt5P2inHX/bkWK7Dbgr30Wytqq27XXCoSlTGCRlqNOA2oBIbxK
qUwd+q+qkPOPfnRt7dFr0Hzv7VtRgWxQek2Ntwn+FmUmQIONZc8ZT2dQAAtehyTtxiIJdwrykp6B
ij7extnVIEpYm30O2l3Zn7+PvmpaCFUMJX9J9IdomYYgGoVbake1ozfY3atgK5QAjpTt73E3LUGz
xMhCbXGAhF3sKEhLd1hOS3odTWZbI/N5RvP7lbeFTTBdXi34ImTzW0xirVR0ChU5XXinFJPlWvgT
EXJ2kDQ6c3zgtc/nWvAQB7ESUI0B02sEC4gVE3rlOlBOrj2HVGBxK1vZku/GtUM5YsQAIXm3GArb
hUZagpDvaXLjmmEHrvjB8SaZSpBmL0rA5Rjtwrss+Fk77fTVj/69PJ756f7mggfHWuV3EfXMbigx
f4Pn9ewgAxgMgTMdAykRgeFWVK0JB4pROlNNdQWRikJdzwDJsaAZ/m3IJb8pmdkbmwIi9YM7p6nV
G+7LT+aeLwkp7N8jePDUqEz7z0zZkFYh2oe72hkFRheBMMLvNKMk7lMl1Xb0NozBE/5O5k0lRxPZ
v8III+hUe9Y=
`pragma protect end_protected
