// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8OTYLa/bbcEiqthCJzgxIgzJMb9gvkmc1DFhniyjb91f+wHN15eSkK5VqPTQZ8pD
7Z+d1WRGRsnLnCnuLBeuSDpMLItxizOC02WasmLs0eP/dK6+5irFi396MgyE+bm7
zC4VYsFs9MyPa5JwIRqeRmVaTCZLbXZjXDR7ryelztwcGIllYzepRg==
//pragma protect end_key_block
//pragma protect digest_block
5Gg1u0vGoKrAxbgt6T1vKiTNMLw=
//pragma protect end_digest_block
//pragma protect data_block
os57FjsURluu8dlc0Z80WFUDl8OpdI3JY5UORucXiaf+EYktWuTlAOS6YZGy/TpB
GMsyiqpJByOvHARcBhbPUo3pfyZs/vLlnu4WPpZU+aNqYS7xNFVuHZF33Ie4UX7I
cKlud464gCjTh3aaJV0I+IIh1YUN89E5NNNrECanjMRy7JbuLC6QqManVdFw5VQH
mMZEoxGMIIDdLZZXbN3fOCwa1vEHKVddoJlVXzPjon9+ev2mWv4ahZS1gilV6iCS
IDxFiDmNOT2KrFSW500D/uf/gtHM0e4hKjVP3Ler4XOcuT0oUmwqQh2wDWQ3DbiZ
BVBc9v14XRiYX8OYxdMmQ5oks4skLpoyCXr+pgJ0XfjgNXhqUSjH5Ppk2Vr3nnEF
e9klJSwxMkhpLVjkWlg1mTRlpb442jU9m++2hwEnMmGU/yVmv7MkACkhiiXhpjke
trsq16AHLYQQ8lEC44ckYHmR3gjUYvt+sVI8i9fqV6F8KAjjOCzDMsv8ucSuZXiy
/IMQxVhQslnfO8wEdbOOkpEUztpCy279JpWzbNi7SOn1FsFrH5QoPra5yrqhRKUK
vP4XecyzMk71Jx9JMhbj44rIonPNzxKrsp0KR18OyjtWumHlBh2HT8sZjPaJ87QK
ttQdqv2D7o9SueSIYgsSR35x4lpsyY9PMjIrqtWRcXn27AP90o6fFVpJ475n0K+o
bGQpZbiIcPX5oDMAmVBKBanOUh//rtdLPhEv0cnNee/tERuZj2gCBXgaxbd5Y1fN
/+ngXRCkqZVfUZWzxCwOfeZYj+2IwG0iK6/tifhPSyCTF5FFk1PCLKtjy+xYhGls
38MkmzRuD0z0LurW7S1XQI6M6K61Oa219tdyK5QeiauoW4DYDE7yhpd9nFc7RB9X
iytaTAmeIK1c0hXecV5uvegxS0U56rTHUJrdoGP1kViEF3vFdz4872KBTUY6WL/T
yk+wxOKQNRKDmEyY0fi0iSmgcfSCB/lBomcGkYumPxC8oTrE6XdAEcSA1+ssNvde
DRtSXWjEvilSVVNBUg6wCtw2eVfwp68hYWkzdLlJwF02nudcQ3HgCe9cmiVNVVkg
DV9ZAdHAirJM+BrIKllWoZjNLuOe4cHfbL311GH9TeKBKzeZBluBabNjt5hRWcaL
hrAydKH8V8HTSgj7vTb9HbckEoB9YPA40Ot+VdCgUGO9G0Hjal61cAIZmQagiyM3
9CBC8a/KAMpCOBMaWZhmyC+wG7gLvlEiqGYzTrUHe9wHIkzaLfwXj80hvXwKxwUG
oyAIL4dccieYDdvwl8irXioCOkPCeI1arTDO09XCR4s4BWdW7RymTXDC8FES8ChH
s5raGapvXDPDb0dwLIUELdpri16nwoX6xL9siSdBSowR+BgVSL9B0d24DEjeIUdn
X0DMGPbFdrxmioxfACr1sIGmBi4bpa3fGGal4zjs+vno3LYiNWw7Hej7+ExKyQO6
2HDJyGNrv+ZoaXnWRgeWYLKmO2ZFOGMQQA1LDMG5C58vLAJ0dRDgkJnXHC7kYbR2
5kXvrCh+lrGoivD2a/87AAlpIyE9sWI8R93Y2P233IqaHUilGCzQu7/4ON7U6nRO
piIiPPuICedJ77at8mSE0nEI1p94JVTEiOtA31VIKJHXEU0B83yRd239fgXxaRmu
YqmZvA0Wku5e3345tbj1Hh1t9VJVhfDvRXXpL9xRxwAN8JF5rM7+GFPoCnxj6YYj
mPlOtdAXG9X8pbDejn+HSqwdBPtGWiC6rJHKgbnpWpXqxF8lbQOCFfYVqV4l+Khy
LlglC/lCVfgyt85xSDc+SIE6H7baHOdQyasSKkBrlnsvjzHumkMVCRvArep+iV39
+I6a/af8j8XP+gFCTM4gI1KjBc4Dued47gnqJTYcyfvsqbW5O33S+u6rHnM1z078
tya7O1BSOfpR1TgNqcUjnnWqLRdawP3VoCiaUgUosDfb0fxMb/hmMBw9SrFk6pnG
nRgsqQdsib4TkmcBYb5LgzBUColuDZ8dqd1IDM9fQUrkfD1+8EMAAUlNjne7HbBb
GQA7hGIyg8hjOv21Q9kfDKm5in65gDr/ZAbS5pgxacmeR6HpWMHkWVVEzmyduHzK
RyyPx7b9vH9UpmGOyboM0/kNCyTk6sE7StYEJZF4gpFNXWzJM/upTF+T9i6/pzCP
LlA23T0BL6clnw+843GEe1bQgExTsF6WFoFTZpZf2Mhuly81XtOJF2Rk/4PWniop
eq5RAWfwSNLl1+OsyXrB4F37xn4V5rj2vf0G1CsWEiw7Zrue86IuZHAoOM6dzHt1
aWwYF8U0d5m0H5BKNWiOKzBcEEXnrIgiX/X7Y1z9BqUKMsb1D/sqy4gSD9A1RmMa
gM9EBfQ66+fD79MKtzKmBYQrXLG7v/txDPdl5t8RL+PCLwgrqvXTktuOs6N4SOqQ
ito0l0s3BF3yw9A6tFdxMEPtSFSjV1BAkzIFP2PrXtgOZnyjI44OqTo6ikMN2AuZ
bD9aQZ+AkHwwszl9hJbd4dtZj0Dd4trwQ1NBM7cgvVOKIJDA9+xYUuIm/r52LkBS
Otpbv6VNzB3sXz5UyMQCCbDPkClO8qn93/b3o/HxQ2tEcimmuKgeQ2LqjZEofDN8
sUpeCf9jhl2s7bczAbzy08d4zN+SVCA3SUPsxC7SAnGbiGq8LsRUUPTcqzIejVL/
LsnhilCCwsZzuowjTiuXVgks22C+T1wrvP8I7dxtr/sSlk+C5u/En7Mq1p7bTN8Y
fc3cSyX1cQ+xX3OcAoSNiVnkpaSJ01q8qyZgbgA5wX7p6a6J2uG7yFfCNC3xEAzN
IYXnWuEWn2fZZR/9FFO9QFsacwbyOmYr0RAM/S3/uQ20tqz5Wdt06PsU3IFvfLLR
YEhxHSyCBUWCn85R1tBGmF2/R5vwTWtdfnQYE4rbUVjcxmN6NgiynMb3Uz/X1hOw
TBRy7jdsXZaP57qHQwQxRUgF+p8IhUuRmZ5b5j2C2XbLekUA20miKsyyKYtbZwOg
SNR51zRf12OHWbIFxbPBPKYNdh1AVTmOtlzvaSyK3wKp5QPghOoT057OCrGY9jLh
BFNRyuqeeB1BU4SbG/uyX4bfg/4gf3TBrUXNxvhobv/1Fu6aC+V0SQ8aMBYVeXSZ
pTVx04Uy/dgZeKM+aMMQEgO+u1NswoUj6qmk2HeHuAXDvgMKczsMgz37eERHLeGC
xTyVA7H9Wl1UUlxk2d8lERO9uukzLamWDysMHhP/MoeshFpcjYWj+C7fLvI7c+kW
ElWcNyk0nf1eyybiqG+/bCxV18EjEM+HK99Jov3EZNaDnmxQRIav07rpPfhMmaW2
KdS/ndgozolRjT9k8nZCs1f4bhw7XXdXnpcl8cGEt2T/Q9/cNijt9zvP2alut+uP
fkvJRChFyPFEy4S0Z9oCA6vM70KdYuZyw7lNIX3iOSbacQ/pbUyLMAaxfDT2LocE
69EBugDhOb6fB02qx8ydy5+GGGAkVgTxiLvX01lwxa846C+0moyjJ2bDFQYEZAMH
7LrW3BNL5B7oFGRJa4HhYjr+6UzVVBBC01dpf1mb0/8UJVmAvuALCjggC6fvKkBr
XWz377EiMdfxonfkN+M+zrDrLW7iCz0nHYuR/fbdn5U8KC/tzf2td8AzruPI9+jh
PjtOopqO/ILGDW+AH5tqZtBi9drrcZY2Fw6fyIlRc12bhGAokc/rb348HfAq7eS+
O3VVW/oxKYW/epMguGYDBLNX89hh35hphsk7Qd3PQ4Fk0hMapyqUtZcfEUZeUNNy
P6ndZ/WZb8YSzeNJwglRNROXGBvQEA3UQTa2rIfLmOhr++nEAF2jBLslK2CwSmHV
HbCxvDfC90RKL/jr1wFDTyHb6C2WrVewost4STLqUQ9YJI4gbEj1bJ0sKIvOZlwa
QKJgXI8ukPc7G794nyimS2P3+SfOF1l+sBrv4/t21SG91be13KHj9wdtxwgDdbq4
8YGDT5SujT9cuirk+fk4eFwjmZQOITsFwPespVL6jZfntV4DZYFrjpTBTVJYTEHB
2S9FLnsQaV7VZ3ui3/b3dzfuE8YziUDzezlBm9QjVI9tJLJIpwCGouyKANB4Dix+
7pE4Qj/QOThw5UJUYEyfMko9ANek3vK0OzE/EUL8yBocoQKThNPmwvS68J1mFicp
OAp0mtVuR75mH5hwgVNSwaFaY+fn8gIzfP1tan6I+M/6LdLqxNIN/3SgZPsdIv9H
BVFZGnaqCz6qeNr/8k7UDi0QCTDJ+IrAY7fpKeasEhV9kYeyjU5dRb/a3uDNPaCb
Eh9oum2hKMw0NyviqQ9hNP0GeWjFy4Mqo5y6eOkUs8atEtqyJKGdtPDF1AASKz3T
q4DEXjfvpTQz5Z9+Fx30YNLWHOFeWw/RiMVmgWh92feD2zJ13wWuj/RtKRBcP4HE
Ot/naiZmrQKN6mFyfSTJWviBdYZsvJm22vS12cvf/6lFkkxR8G4qcnSID9QT8i37
2asmQr7/qvlOm2zdMcDzgapdJIRo6i7fR6PxtFzH0NjG5oTXEZJd7D4EeLeThLek
zhP1uGsucgzHBKwznABE+Dtiedt8hCbptbejAVnuDwajsAeZcZ4jAUFtu5RHaRcG
HBgLYvs68eX1kkcBoBewK4B4e33hM8jUwM5BBhr5Ud4xHodIqgcjNXxkTaJFwfcF
nYqoUmhbiiQe0Zp/4e5u86K3+wd3uG4jVMjm9Fo0txSRcwJipWsKaTZc0I9uUKdv
XZHaSxquKrRxh5fpQQzpYHQdbrjrhVBU5sFpyYWK62cYO5nzrp5HNtdkizdSHpgS
6NmzbKEsiApWipgfhaPERKie5xm9kLfHUtKIEMS9H/0AK8TfK/9FHdR+UXPOABsm
e+G+pT6UWR+fLVmCt5R7HorVsnF4C3ec/rTC9PdF+Cc8aKq/ObOAsyu5SyGHRgRI
f0HwZ9S6HFbHF5j9a/ehiVu6ex9upZo1wnXwTwcnjpiU8XJlJP327jIDZSdni8Zt
axuuu4UDihc4wrqu9GCfcGrMpbOK2GHk2kgyCRCz0WToa8NfJa94NF1+yvPRKoim
CxERYfDWldXZJIDhlEW545gpp+5gw7/FLjhmnBCPk2Q8wSU6+bwRRoi+VRry4Sqz
EFfAQfgo+lmPKSLZXb4I2D+l8J+EkbKOhPCFPfsc93MSx00p4RFMoNYH9k0Cyvbs
NX7XYr/ByN6HXLb0/i+Bb/i+kOo/lFOHgZJklmUOSxhVjzYJ2SadSvIbMDMK+jFh
ka2xt2XgI4G3gZr3PwyMBnQXWgQUa8pY1We2qJSxsTmXNfu5X/YHjPhAvH6F7P+K
eYXaq9hqDvjIVFnRSJd3QLxjS2ideWjvD+ynZ/XPHwFx9I7L37omWcuJs08Y+VOs
Jk1R5NpVguSwlnYF+TbhHLfrDr3px/rMyxXL2TB4mnJGVBFOT0b1wPqs4F+vne70
UxybNGqnrMOtZkLDJU3NMB9ayncwP2vQgJcyMU83sgW5hYHKuKltAjDAnwEIzOt2
1g/Cn4Rj7vTn3q7X6YW4iNuKtYU5Bp7fIglqNbvRp9JTJ47b9NHBmfeJNS+s8l/0
3lQm+L6ry9dhd8lVLk8YcGuokw5R9vx23xItv1Y/alEM/IcrTWIvZJOpiCMyFY4l
NHRGwm43Z0XFED2X/xH3v1KDy4InSlSqD7BRcepHCTwJ2fgvlt4khTrino4aORSN
KAObg2rEEh4fO6Ta7s93zVPXQ5LLyflKAlG69/T3fjnhCfOd+RmvMcnooxIZu9mP
83RrdKdJIn6WgQU8K2LCOzvB2/7PAjeQ4o4227o4Un2LaTHvS8AQvZ/5Pq9rY+m5
tdxhFLlq2VGUoIvGoFAOUewTppZGm+uPFr9VfYNf4AkhFPRUpFw0HSVxbluBMa/G
fboBo06HGvdlRNFZGxVgnDLII1iUNTjgKDWDvE3pfV/ygOU35aYhxTUj7qs2qriC
glLY65DpTObF5KLuqhycvm+Qjl+G4FZY0UgtHL7n25A/+Y0E1kYaioi/RPsUDaGF
TqeRjPXxKHMuMNoAIzKuSWe1bdLlOe9irRv5yszVXaQ9YWjGgVNTgPqKf/5lBxPN
Kk9leozhNXYoXgzzygyXXNUDjLd8qUnT9kIs7ErFQWcKMCm3sv4B6FCIJBw+aEwe
o4cvoY/Bi+NyP+AImxAIEAqdivRhE08YGPaL9SbkrOcFdQhGh8LKqzViHiGEujrf
hlgZDwjDNkSLE6HR+E3lnqTHFH6k++61ZdILI8Y6j1VFnhBDNV5AM7yJWwfcEH90
r0ctJVB1RYpwtx0HtK6OXOAs4Bj6LgVxAkPE01+mjKKVJ7LCTeGdzfU3LpI3hja+
FoJIMT3QJNFRbueUOyKS0r5Fkm5tRvrKwOtJXQq9Pse9lyMjJaSfklsZ/JQyfc/E
HD3eRmn+dhfWzDOZCeRQvjs/RHGQwZBlJXxq/PzYOMsbCYPcTYx//IIEs+Tb+4bH
a0tdiNfejBixCWz9A1A6XmqqJlfp+s5/OtxbFM2W9vBZo5sWTHfH7VZEY50V0Te6
AwJx/Ey8yYzi8S9YnbmG3lDClVw/ePliMyUuoa17Z6EY1iZYZmxt3KT5Ve9CjBdW
mtsAX5+4IxxGgm1Ysd5/M+/Njy55hJQq5wB3lhmot28nXv5Z/9EzNIdD2z1y/8E5
UhoMantsNQsIcnfY2liJabMQCeka21zE6Bb8RioXsy9ufmymEy095E1zCNu0pzKU
3wvJpUdzH4Q5vH5tyf9zn2USVkDJlvU50yF/w7gPHa3lFabZ6dnzCuLOikAx7/z/
LGG8EK7GiDg0Hl9i4D8tXNSeB6BrETuewdAWxK56iyEsedomMSQlZkpqiv1voqhR
v/D9nlrLTmF/n0S4Rc6PRyeZEc1EDiz3+taou0hEUhmaNN6AkEVRt67iCO6vXbqV
bvc/x35W+gB6X8lHQjNWkPLsvNTIk72Jf7kcB4Ft+Y8yirrXX0CvFBTou7Hw94ly
KbQThni1lIzo1donOLVo6+b38plEIKxuAkCHTHSTZb55yuDKYJ1mEjuLcidntm09
C/b+a3jadYJu2/xu30/aK/RBkhGUtMSsjc9g07Eu81hN2/LJZX3jbd/VNo/sywTP
NJ9k2B1SK15bQ5/F7p5Im5O7zF/bCdcfMwQbKovJoGPAXS1OkVCdxLm38MK0nWTx
UqIqyqaIAtj+qKxua/k52BOauAHMlioOJkCYAyFVK0l1X/Smhm62Q3McgZwikcgS
+DL7jrmUy/sApwoowx4VbJzQ9lrgVBZ7E4wVoMmxV96oh3YUIaSCIqovGj2+ctCg
kwNYnU5hC4C7bt2cY+BXjG6vw0yNpoQ4EKRAxRmbjdycM4F7jcO8B5J9idjbXqW3
1/dg3yUtASBygvNjQH8jrN3DsO9jHGwZSib6EsktpHW39s+Ij31VqL8aVim/2H/4
BrRXFKiE/hWc/UfahBoFs43CzVWl6yoxSP3JvCrlmV1NGw5phFu2Qt5Eah5EEhGm
IsNkAYryVQkl3Y+/J3rpirYmUIDGRi3KP8H/5RiBviely7ChjItBuYWsGj2FkCjj
Db2tr3ARIS4uONds0Oknq2oRxqkNDxlIvZxy0Fx5qXeviRUAwtZmkresPYC6oYYy
fGWl9xi3tJQVrikBqfxJf1wwm0WbuZWRr00deWi0CPbM7TYExBMKpAvbNJr6t5Mh
AKMlPFWg8TcKyKKzQa1irytvxPZhjrTb7kuLbbqln8hbelSbXz1+Lkru5eneXJc5
yCqt5TWfYdQG6GBTho+u6pTuIZ//qqJIwab9T6P+CQBmgKGLPBnCP5R2Nv4x453w
0b+3Ph/CtHxGAkXHmknlw28+b7oP6THLbng9NKrHjg22wTk/AWy5vKBeKVa1MN4g
SpOixCgLWpKwuzoVx50YE6wdCQ/ARgW2ICJi5I6PO30WMcIqgXSkMQMyBaI0IdMD
qJB4DK9AhATHxDf3Fh5O/bhNkDBnN9irX1UtMTylDpUJecLBNe6ok9zMTN64GWVG
5MoV4cMD7cM4lfTBa/QMs8Ch8bW7yUJbdIqRGTeYOqH7fqCdN4URc/sdaakXw9QB
xFyGug4wJ8SBN6UdnRkOtV6G48hkxe06vBJeTQDMdD2HNyRZ4IzJ0edwFQwd8JkI
a53E3nGMnqSsmRkSPZ6ilF7JaoOwEV9Sut7pvE1bD9GQAoqzD+Mq3zmD3UqYnrUm
FMGMuFIpiKvUj3Yc3m39+fzOJpEwlPd2DzeQQYk8heyf/n+CnFPe4/Qt+4U1tGUL
H5tWyBygdy7vJPExVW/vdbIrFE6jK4b8knusAyrW5Wd2/gktDrBYSmopgYkdAM4A
E/IGp914yrv5/81g/uDqaJvTszaAcy6lPsV2nYQ5BHtthfNKpKRC/fJoy1kgqEMV
Y1IRSIsJVJMxyYTQYDolSaTV4y5mfeA5ibBxat9XmBg9vExahzLQK7iMa5DXWTON
jPZkN2o5pG7NmBBcnBwokbn1zLjkreapbqVtmDmW8YCQfSGHHa9yo2N440wtG46/
OTRpw3KFfZlHa/3r7tfV6tUhgkLdTNBTbbFNJGgMbI+yhsvCLn85oxsRJFGCdeW5
vUcy1EK/keB17xL3HFghbSbP2284GlXkvKNo5K3p8rJN4lsuQmft/iqS+6/CUsIe
Ot88Avp0soohVFdJR9rzJwenAeZFEuq2duDfjXIVUDZ+3uFotfMgCiKQBBiu6iAf
bjT4Eudt+B4ArRD3ixf805r1HiEnaC8R3iZuxN0eNwUx8LG2+x+sgLI165/GO+QX
0qzFSODyxvtkSPJ/J54j0o0elkRhkJYv5jwnW5pGPQ4C3vaIPBL0ckrr8oJv2mPJ
0aYwdpG3Q42f21afbLDwEo47R3D4vLTjbg3X+uXSKdqQWmwyjx0R+xeg2XKzCH7A
GCajHQbSS/80uFeTyjMQ1jCKP/7tO0AZlahYBU1y/i8fZ5EApzjL6LsWXtrVL6bI
JZ2H4lnV1UAdGvnYkQksBLazqtL1ia8RRofVrrze3b5deaRVWLTSF+nnW5n7xcW3
JYOP8plir4shivKcQU895HwQJceCjcnZqtaIjLtwxIF+Rff17d5mT2Iu46CoRs/d
tI5KQUh9RnvihnN3rJgCf5QhB6k49CbGH0Z1sWkuhpsBfTN0XoZWDQUnQpu7jLBs
/c/lprnMGg9SRWn9sxb84ABoRWbQj8lFt/OzdwXrbnxSIzpZLErJNpVPtajZ67N5
A0BU8+k5lmlJOtcdyRumdBwPDZAO8dJk5sJNnn9+Xn0Mt9Wce5GCbvmykE5Bg70p
y5AP1ZYHmtkGMelGkcXybtrHOP32T4g9OS6mKzY0aZ26eaEn6tFsFj0rG07oGCfQ
IpxYN5QnO/JZpAxFj3kvZlZwlp/JNbxMRsxwHw2lVIGO8yzZF56GV/FmYlnwOZVr
3wGx2dau8hl+/V5H4TEYrgZXkqsDu36B5EnRS9izQpxKc0OIt99oLmrrS65wJ1Xx
p62XVdLjG/FzacLKDhJVLk/JQL/ayMuLO/rvBbKEE6EmYjRBOGEKQoRSI5vU8iZG
cHCwdWjFciNwPLjBZ2Bgb2xSpiDgFMkbjTJlDsnxpJ15IOdtuglD6CF/eTil0U2T
6TmNBoruZkD+zXOQHab3FH3t4KMjZh05a4sDtUoIaZFzk8z1vOcfsxmOKTvkjp09
zej7bN9Uz5RTz2fHpzviskFjWzvf53H5k/gpGVTHNhyG8lPzQMMUkqkmLXHD3o37
q/L4orZbjk8uY6Aclt3v8SXNwo8QUHS7xzreu5RiIR8GMo4KWxYHMgh4PCA5YR4/
TSuWz7xOUE47OZ0CdZFUF65BulLq0hD8+pf0An6rCsPiAPyKou62lCfEn9VQp2ok
g1gfnr3yXdZx7khrdH1+TIL+svQxyNeiAc03zCOlE0so4/YhotjAMngFFPGFR4FR
uRlRH5uSMKZifh5Tgz0w63mmo5xHh2lPVFmzYwhc427sXWBLneqKq8pgl4ecKwXt
6Afln2UgXcU6ba7UEXXF9fwblljZEM3T2kfX8QVwHThJchYfTsiSAnTYev/GIRx2
7vEDAImeHfzNPc/6KhofWd7WBioJth73oNujjXLdYA6Rqrlr682aIxb+KMQcwqR6
D53/B62h+mlf7b3ezvmpEZRESkfamZYG21Jd1ZWQi2XDZprlXZsuDZ4/hivKbaMS
+tqMPCGYk6r9hqehV2liRltiVvr8PtAIx63iazytRRF/+qiXOZ+gj7E+8DEXzIi5
hrpveMMRZlcPaqI8xkdBxkn8kljV6UfOlkLk+vRO6bIDMoAcjk1WMaYyWO6wgEy1
nNSigzfCD+BciDUjCaMRsEJ/2huAbRVwZWk2n84Dv/6QxhunK+OhFgGMejOH0sAE
pOwFTYlX+HPh+yasMlvigYxGPAgwZch2kAYybFGmkcnJ1GVwl5mgcLQuQ7Ryexse
+QMosmui+uLjxOQiVAQp4iwtWm0cDCSRxgRTSFdT2+DscJzaFOSyaT2TM8SQADma
wc750UpyJgpuwE6RFDG/kLCUXWDSMUcp67pA573XMeU78SqeGNN9/uBjfBAcyfm1
aMOKp2X19pZf5/8bZ0li2u7YlMI9TebVBJzkQiqQc93M7Lvk4QB4a4vH+o19AtoP
eNHWzBJu3D1uLja4QocnIiWPKEx/fDJHkV5PyQKqfy2ExLekPEBDOmeHYwgR3Id7
Tw02VyTaZiHvSeZ4t0iWGxE1bPQrnNcMxvXPmBtzVN+dknx0Hga1CnOB/eFdoa2L
ogt0bD22MEj0hShywyf+QfzPleYpt71JzSgg0I4FFg+UThnc433242BzDi7rV0a3
lYxLi6gPxEcI/yWy0CfFWaKmpFLwdobKYKvHpfnpfTcHbUCQMWwo6nYvHfScH5yN
mvuY2R2fOIuz2T4foIqjJqc2bpcaAYzBzspIHBKKTX0NE0hIOGL/mx/7NAZM838q
5DaGrVPHc2cUBL+L8iVLT5HLYkZr4xo0lHBHrDWEs8O1IfKTeqoJp4kVYgHWVu61
GGpyhSsRh20OZyFi0aQnGxHxOh4bGeRHbHj0wjPedULCGyf5o//kkdMoXlrbSRpe
0CKAhdhy6+sLrnihcjqdQIrCx31eEIMcHNaKpsUPDzTWtl3d6JLce5NyLAzMYBXF
CCoryNx1KEPI48rbBr8gxUNT12enwa9XHTg/tIPqv+k9fBp6wgrou10O2tC1z+sL
U7j+pEXSDUGG68Uep/2IjGMpj/32/x/gQ+Pk7PzMYzZchkdTmKKsLNT1pf4vXGtN
Wdk/4DHq6s3Hl8b6tHM0PnOHL5Rb698geXEPGLOOkwRxsya7GwTAKZhovaQUSvkM
0HJCtOTBXEUnTlWpLo66WtNzVNh7QQyL5PDTmWaE+lAhzsDpRmsl+9vA5PQJZX+V
gobgJ1ZltgX3l6meElbe/NA3cSXS2XzeGWoGbsGuSqm/OEoT8rgJDIM+2eCllKGe
4O7ZMku9hEhoQExeMbStU65yXk9CPIB8nd+Ej8k2qa7M9WHjQlYxEhmP4m0UfnRL
EpGm6by+QLUMiRzFLjwaYCTW/wVYSMUSgt1rccBTkcisAbgbFAmHjmxBkj6DHtz3
+NwWSQmqCstfQIVzMPuU6ivvqTI4Z+e1J93w4quY2rhtBYtycF6QgbLmmLfBwDo4
9vtRtqMbX+tMnPJ1bFpDnVtkz1pZnJRC7tUStIoZwhCB4gHngmwvh/viYdjdnPNR
cZdepILyLVZ+Akr/4E8o//enxCHfsPw7MOuGu4DmmtRM3ngh7S/DGTHChNv8IcrC
IMiiQJNxeRxJSdK+n1q8jqHO81hUzD4moKa1VCA/tMjgp8xAtANdUbBKJ9BN2whI
IEGj6dZAJ3z8sWMOHBj9oEVwUOleWU+uHa+bblKYIrw4RQ/zFaHfUijn/EX6d9mD
/RqrHIdWH8Kdto8Fr6GGlCjbJ/xK1M+/nvunQgRL0BDI3cwldrMH6GZkeEwMbvAB
1O5/yt8ep9O0Na5A11vrKYAvcXmTnSPkAgMf6sR3Zq5Qb2M5J/gVNp6GNTNtmcz1
+hDvC7HnpD0UvHZ2i6OFHO2ScBv+0Jkqa1jlhjg7SwwqIx9V5DUaK90zOuHQZ/Zt
fhqPeqLVppq9cZ1WuPggn7/b3nxS94JE4xy/qOM9JyNzZM5XdFEsLckaSVYzs4xb
i0730ahFL2Qatz+QjfnEIzWKPoW0cEjliUa/IwxrTWndEX71ejD7VCggpwQu0LWP
MrE74e2zeQMgYh5MMHnWs4+oJ6nU9sCRLGO6+n5FqJK/jfCK5pmzG0Z9FAXQEll9
yTuEUlhmpEO019yxcQfS3CfsWddgDc1k03ayLycgSSKxAp01UvtLsQnwVmiH8D+6
hj3YsSrvSTmvQbZxkbg3IZVTecbxYGD9QtRIYHC/3yQbSirPi58Jbwg/SE3DAe0F
JVN0Elj1bRUdtzSKLkHeVHCrFS1XLxZB9sntnFcsfbgGDz2o54dvCFQK+XGwe0Za
2Jwji7VZCPn/VcmOXbnS/o/Y1P9dgObBG5e9IBPwiNtRbbYu8sd43IRPYJzPrMUe
zXsESq0FhMo1PpEiU+4GkjV0ErPPkmZbARsHgh5nRA3ImDurvlrFRd0Yp1mRsmiJ
T+ioHt48CuPbTrJ2mHx0qPTeSJe4lNrYggeCJ99rl09feqVyjcJ1bSAoYJo6VYJa
MZBPLF5BIiyUkWj5oyucgaJmEjq3nmSfaSTLbnN61pWJjDqaTMry3UVRTpK8uzl8
Rbe8wgRnj9K7LFb+qQ2iABIDaPJMMJuHqO4P4C6R+WNUTvz/UyXHviEPVhqq9buO
tWdEuzrPa1iJPYNKrRJFFwL81sGN1R37tI3Lj9Bv/FZ0/pBrZOKCOqg7M+h8Ty7i
+hjbTOiqojy5yxSrLNUNuleQPEMj3DWUa4Myh9zQAfA1ZKc/a+0eTxODQSEvuBkZ
Vr77Shl4bcp9k//vO++N8Xlvz6ukA4E9hAMorZ6se14AKKdUO8ejR1IBr3J0pSqL
McY0212EeEfCbL1aw8pzBw/ZX2zrd1SlEKGjubg676hkQsRH5ZFWGzwob3qjuRmJ
QBQqxqqlo439zGgOpa50WnoIk5Se8o2UByN+Cux6POsYAtrC+ToMsYP7U1/NDFR9
PRZeOE3ru0Hbe3eCezzXzBnH/QkH9rfHelJ2PCu/gmGFnzMBG6xQtukj6vQOjZc9
L7nBcCh76Wv6DZ2wA9yvlugptTeZbFdtO4t7hCJXuz9X/2QKFUjnTBKqRNYmg6eO
nuOphhBvYxTXfxyaevh8O9G/S9p6WbjlsNCAuRKS3Zf97bSMFcGHA5+nCL3jOEpX
eOLcpTN/P2zDWGmShcXD06OWJ17GXMbvjP9K6vSeqG0trDuqQoXHS7K8O3jTOYDM
fmFANiDoyyOgMirmHkK/vDRmxDAA+uwYJzOEoCoOPl69Cl8VNNkBQn4Ad/e/hydT
wtpLUSyn/CNRxhplrvuoqcdqRTlH0onONEddZV9a8VsLvBc6Jctfr6G/extdG67Z
rKtReGQ9Mh01dCMEGV7Cv7u+AfDNdZWyh85wv06HveykmfAsSvgv9nWoat9F/f4Z
JlU5vH3JJmeWBb9LWGWO0tvJhi+bNOciYclfzD42BQgPsGej2ebdXMjwLLDQXTrq
TekeYh6JOLRHI9131c2NqIdQTO+cCgwePC8gvBmWeW8YQNPkznUGo24lTV6iHHAE
iHCtmGfCXy6kicYKK9QD4qXwhwxRbedrWcYNfleeJv8LIPizPmy6xw1JVe1nPFaW
4jk8n3tNjiLWuJcw5RmyIUZFz+mRUiJY5uv2hTvJS/vvaliW1gpDaoz89BSWBFhU
JeHCTylGIxsQIBYPRp3GS4nWwKcWIR/V87UgiBXlkw6UYk/zIbQsfF/7ZUYNXRra
ozrnY4b0n5ZI+iqQVHZfTWTFmD7nSPWynqmzpQcBNmNC04mPF67M/SsMEKwiugq/
xwHONSW06hGP9IIuAo3Lw0X33nG3ZDBcXITrBm8F1VGv5OUP4+X2C7t25fu0dbZC
2hahdlpkkuZqI5bVjLEMvCeTi6u5tvc2eGaNUCSWavUr/x7DtTqkASjRoNxAiNE3
clpOUHbr9leseLSSwSEOrb4I/1GnzQg0HImdfkItSzWxLrS1SSLmssI3HOsPtRHI
xJEFqZA3qbmbX/nV90QGHoisPKFkX5M6Fc93ZWqbk8YLscgb/abIOHe7Copi79mQ
0lTdNTVRRGvZskhJv/TOSjfjVk5EmgMwUkLazr5xgOZN7sYB6L46PI9P3Nt6vWr8
r8AWy+/n1iFkuaaqLeUTK2U79w7Qu7Ji8udRQaxS/UMxepBCfrzWqpPxYsizRz32
jvRkW+EoXE35j6H3OTA1VsB1v9lHIe5d2I00vA7cBTikaNXq152s1RVL39OQzwcF
NH4IZ3ER+YSayTl35oUyBb/rNbHxTajPEgnlOps2pvpar39ZEX92CD8k9u7c+8Nt
/lZIEtFYLhvBZu4H1XBHocteB3/SvUDuZHVqF0ZoqFFDy9RN6gxlixd0IqXQ6ZL4
pSOup1BYM3wVNIL/XUQ5xlt3mreYr+KPFtsXvZ8WxFu08NchH/bMiXQ0BdHKArHq
Oy//B/GHgEWeUZhrnkgDB3iFKgMUMi9gwYk788t9o7DY3EtG7qa3UCvb0Cu5wknO
o3SldFl+AobDRn1B1T59f7sNwbWSr2OvBNVC7qpW37rS/nUKT4o4TU/hh8Ik4mbj
WjDQka7ctk8TiEgIuZkDtTIBUMQl+hNdbH0F4ptwsxg9Ic8jMqcYiSjvP5sUZhAF
/AAFlKUqZGw29GEc0O6rNg/z+eeNFwNxFzTdIuVwRqxdAMSUncxNY9vboFuUewpX
W9K3NChwvn9fNS4VvcYd6efbYDxG5cbw0aE0wY0NV75qjOWMNCrm0qKFCH89hQ1P
DvlTPQx7GTG9xBNWWNXR8jxgSKoDG30JvOVBU+UtL+g1l0hW0/Wbfwy11HsDR8Di
jLk0FAvniDfgjxRwdL0IzGFMDBz5YEKVuML18/6P/04EXFGygLDapZ3P9+Nn3DO9
xTAnqCX0Zedm+5f6E/gOhuwbChD06DudN0GT5WS3EuPhfMgEYA143lRGsYmyqFpY

//pragma protect end_data_block
//pragma protect digest_block
f/eXDcnUT9nkFLbWct7ltHuLhew=
//pragma protect end_digest_block
//pragma protect end_protected
