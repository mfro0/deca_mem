// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:45 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ILI1yzkCiBi6uj+hYRj0hDjvYgRc8nErI67dYFhQLMv+8A3kn2WmAW/LBAUcXzU5
SaPi5df3TKBNxhC1sOtWXEeSIBVsldloEJuDbT5rDY05TB85QFhrmanCpSTYS9J7
A4ZcRuXp1fzwHyuiiXUtfKGJfsJzT7YmtBeQTThA2zg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20416)
7z3myiujdekEUzdit+oz3NGIuSbg4+5NgAGozScNh+ETrYkbgONwATnFmcFObE/l
ShKluwjC/eJwsAg33EYMJHtDFBu6AWjGU4UVxLxHkjdjvfrgiIWp0cFoeOZbm7V/
LXyq7gN735+vD7YFWdfJ86HZokoq+EB31zrGrop+N/4+yEbW6RyAhA+BiZiFaH+3
bjBg1MxOE44Gn+3hPfLDjT9GPOVCVCObEAdKV7aobMaU50dXfA+NSv1dR8LJl2W9
S7Sd9paSy1aJJkKf7sKwSVNRYIGzWd229wDmfNHHZ68ZvS0XpklYz/EkiQTEwiP+
OhVAyzghhju2F8Zf3SfoL26Sp42khuSqnxbqg8o4bmibOsTaDhkMu4VEhom9cNlY
pCQ/1wfQTyo5asOId7mCU1+kpxPmgauUz/FRbIxyE3Z61velB8msKFPimBB6nsAQ
L7jBBXSMFiTtFMMp16S/87uc1caIiNHxZPp2B58BsMAJMI5gdSl+yv93WEMlWFUk
ec9y7jZd/1WzBOs0df9TSd7UbzRQHAVKtMUyr30Wy7Hmq1GNvpVabbouWvGFNytk
qFevzV50pLu8l3loJM1vg/D1wE+CRTrNRFVs4txQJ8UV3RLropwfkhEwuv9vofrY
IHkiOpeEU8DbEK2GGlisL+COv8tUE4fXl7eyzkaNluxFjarGs1jg7g8qD/iOQQpt
98ankIRI1ZKYBisJqjcWE7l/xJVP6ZVxX+qAv8yaNWPasm1tMwSmLCs4TDszEJQj
d/tpHjjQk5iCE4EmDqMtTJcDjjqSrd+GwHeA83CVlNWFhHbbjbt/v4YjwgJuafuo
g8N08HWesBNb3DiU88wyMtIluvwTJ+2DTfML3RFiGS4MnLaWzcCKIICWoUC202nQ
iVlhYjfFsgdIZ54NLd7sY0feKt+83oTWoOjDNx9e+o94MkvueaTEPUnnE15XRUCo
biOtKhvykKoTSYEx96JJ9qeezIsXHauFgpN1hWhAJNEwh8TNcP/sj5VTIRxfIX+4
XfGHFd/OLLAgkrfWQ5zHx3ZgR/Q2UFvwkPuCPVPBNo+/VK0v/O0XKNYeoqUpbreQ
weLjPhHKAlZ59ld2dqnZlKOgTsMnUprmXrvHCyQxeYxklU5vonc4EOwGrirlWJTA
zW70XLNWvMrFo3PlXnAM2v35l93/SSIhD2+GwpbvGJiBb2KjvODHyP2MJLso5xDx
Nrya2v+jEesVw//NJoDxuXetnYIxrUe7HQarRQJ55Pz/XJCBoIk8LFwxoHzTFYBa
1pv4cleUjsj6urFCSL/QDX+MzqrNAEqLIQom0XBHhwxhuf9aFVmN2iS0fReqIoEC
TTF8zIdiujTRGL9EzC0U7Xq6tkDgcSUaYKIZ2VMlmwsyQKyLRNEXaSXHq7lYfTLs
Hk7a53HIxh2/+aNaa2o90Q729FlSNx9Gjlp3MKwarqPwzLTJqh6ZaX4tcettdPMW
3dpLe8savYWlxC/1FB4DE5CrvNyOoikFC9VltmFCAvFABBPtx1G6O1uPi+rpxgs4
UUkr1q+LLSaqD01UA8QuVTuudZ7j4NpHcbgEUp/lF/AVIx1PmHtrEBkrzHTvZHWj
J7gDjS4YYKLu1fssQjLzs94rbpe/OE6ZKz94W95RwVrY1Npn8Q4hnuxQjKd0jhFL
6xjcYBjT+FmWzCUlqyacA+iYHhBhnkUiwK8LpFPKDZ63EbeRt4fQuUWLZ7kspQ9w
o2WzO2+FLOKLjkLR/DTUdkt22mzbPgdphmPpwpv4093SicZUVyURfO8MoppkdLAC
0vLxn7CAFgYyFKgBLaXtSR1+HG02tqIvgLohUG06yl9CTYFHwrE+V6kSqMc916Uw
soNCTT/jRuiKrfsPBI8hoe4hrluRjgAbSFHIKDbD2oo5xUi58Rih2LdNEaMT5Ev4
GD6X4b6PRDkScu2oZdfX67sQSBZYlFSbZmkfg7fxBDjtXh6+1JZuk9YE38ot701B
i+xTj4j7UWF/cZETRtGmMKoA00aRV2HL1b6UhRVGJLl+3yIx6DEKRaFPOVAWoW5M
poM4DTZJS2pugDh0X/Ge0Re7s3BT6jDFR4nx3gf0VgN7V0b94uqyoQ4u9TazKdR6
wwGjM7EdFldcXeJAGsRqTw4KenuN83rxvrSOaTbNDcl29aVjxaonciwJqkvKdUDe
vDpx7MpNeXZat6xGQD4FcGYRnNQHo4UpYtWXY70nzPOxRseAUk6T30U+hVpk6AJi
05cNT22YupLIJkMPj3uml0hnEcJ37tIhnnLqJN+oBM2ZTKi30icBOKmvCE9oK0eR
HzjgjIn1lTp1ErjXwen0j6IPsycDQDDXb7Gd9sYBpJUlkB6k8ohwxLonJUay8to9
uIwF7LlLuTeQXTVWIEJSxkK6C484Rzp/4xuhP5NXvZK2lAxJg00fsuDfyVLpuDWB
9nAjE1vTsODRit3v8KO53eUEmmqlJDI5TL/AeGJCDIdGYh5Gzs86fz+B2tDcHq0c
i2VziHgBzRAzak9sQHmsV6m5wcujavfB6DZfcmp3w0vI2iil+nusssNeC+J5w1Ex
28oTSuHSkXCSMrsfzpAlfgmTNlJJ5HFHKL0PdG8MVwc/epk6qY7GqML9QuJn/fjE
kmlMrZxtzmMnqx7zO3290nfO5Ds3aTGITu146NPjBwonz66z6bLCVMIrTdwTorG9
FjsaI8vdUirsA2ikOD32a+QE3hw51tBQscL3ZpV9ywWOXLAGmWsIUst1/TdPlNjQ
peEheAJJZ9wIQWiSZEZIobiiUJiAHJoHyX/4oSibuWYVcSYFzV38ItZDXvLZhei4
l2vBM5xoT98iMtN5R7aazwVy497cGdQULZYSETDTKeDSOVbsW5hLkwPOYABSTvhG
0PTdU7yY0niEn/F1zxqM0syLqfgVs4T0A67GCW3Pbwa3IvVT4v9yLPc+uJpLQP1U
L9opPMZNQKYSBN8Z83V6XCpsbZrJEFABLNQD7FG3n1fnzc7DM7IQWcwT5DnJ4Kf7
H8HjhYVD9n14fMvgXQhk89y2iDuX82zOIFxEHcmwTw/NooWUT3eSS+6o9SoH3RAp
4JLtV/RB1B1HvE/zp7F/DW99x1UgvXtKJLK4BlS+Qj+8veelkTF6oWSpdCck1SFh
w2DbdpO9YbWykITBDMTrixQTxJc2xqhNBbZzT+YIRyaw4mBV1ML2Auyiolg/qC4M
chwTO/EMZB/yKoZX18lUwXQC4Ae909b8XWpHHrgmfUx7k07yVO4Bj5yc6YeoZXkx
XxHDQco3h5N6dYM+s0a2pgTchBU6e1uIXiSY6UNYMT7D6rNedxqNGp17OjYowqUa
6A7qtBwfSiNeOwrSF0OVHPhgX+03w4nEW30NnTRFfEDARIWSz0D3HF8TJfGAMePB
bXGzo6on79P6LrNNlLboYgyXEkIWI5tASp519vSjERfFx7mCI+kzX+qMFcDqMSe8
Q3F/PvQ4v/34ekz64PDklUfGAcAMlXS3DNxry+iQhB9iiwLUQGynBY6f314BidnN
cM+L8rt8tEFgeTUGBL5dq4nmxaEZ2iLYV/+pJJx96SC90hhxX7P1kG12tAJuZ85W
TrTNNXsAcA5PA56jlt9WYTboUPS/7EY//RkKmMtROpoxV1bmG/sUniuv10lDZwgU
AhaCEjb8jxS1hwIfC3jvmjC+cb5fpcq6U2lnBwi4qxutt0q4GA/f/8ksE4tGZ/hh
WOvRRH6PM+R4swQkEDJ2Ycb5E2NPy9ziF91sUmQXOfoTeZ1PeW+l6sc4wXlIwGg0
7ecrcTLIdOoWz0IbAtjc9A/ZigEghDMmSZ9nbFeqen9thh0vKW/Ir+MlGFyFUqPX
xHwwKSsNWqBvcepbVp40GaSfE1xOTkVdc0VUC49K3BZz3coiMwcp8M9MofrHZdc/
s0+6ML4rfdXUaZ2joIleZ6YEtzI4ESTgwA+UA8Qz3libYg6ICRRAvZz2ieMN9NYT
DrDNGz94tFTxkPUlzFP6k1dUZKxCV3CN61oUY7Wxd6HAE+rf3spKGEFXQzPjc4VT
ZhyOzkMybPw+nLbef27qXi+Cv53qeCMqJ1G7jtS9PMAas64atgCNP6NE7YeB/r9u
39tf6m2J3bKgsF2uWnzg3QsTQulbDp4T8D8wZHlwpRy86uMBkeAnWz1n6P3pm6st
NW52MXiKaez2b5aX2bCJ4WjDw0Q6VtebisvmtANNUxMGZw7zP48qWLMHAv1rF3CK
GUMEfxoT/otpRC5eb/Y7r2Upbl4W7fbxMM+6PF3j2uryGun7guQUxqY2DMHXeRHR
PHV7kdQxGLBjYDbWHi3k2NzBdGHHZZk8Pv4wqdLU5wOy1Vw1t8qidZ5MafE7DEfJ
2TRNRkBsCrT5YCxX+oigtD93MMTrjXeTgbpoBNgQS3RvPA1oPQrb+7gDQVtLenUV
TZ0ZDsxqTauiVzCVYhV4aCUOVJiXFywhJs20bj5OYS72U2ZPkyFg2W2DyRQKlskw
wRwOSgOTqc1FGOKzLQjKnNDcLvWo66nkRwwOOYJ3QRLKSdQgnkuZBBOBhp3InFaV
5bSUCndZRqUxERWZpT22Sy4qokDvkduCjdfWFpYTUSCJtGj4F8uUZfVqvLb63BSU
RTzk/5oO/Skva+TIQ1wwO6cBbiEY6y5HcogRmsaM0b0zGcmnf/iYX4uxTWFeT+5I
zjoawJ2DABk+aXJ9P4/rNPAI3EP+d1F2ycxR8t/d0Snibdj+7C0L66iiBte/IeCK
AeU6j8n1m004a3CrjkVUfEccUpXkNXjDbTxWtHOWu0iaPMZDUWzP0S4F8jh0I7U4
iIy3Tw4rWEXEnhrclI95ZKKzhx1sxuhZZPDTNaT1rbbUZxFfeIaEjwwSIedeQY8o
WeJorvmQvIzhotDDGV9Dx4cPpp4RodSqADfhybuGLpPyhBGpkByWbvGDQfyzw8lo
eeMzc6ONW2cCJnTBGe8yRAo6odusTz1ZdWegf2rcibKTfZmnYUlhUr1etGnHx49M
70TaZy7Hbz1tKmj1tuIHEi4jQOfcXFjShx6wfuI/GaiGxTGQlkVNUXrWccBC1jqg
fIivEtW7NPXWFSj0tMG1RNzLa5T+g7t+SjMm1c35v0oLiSlkW7BZo+5L+k1J+vzA
jT3g2TZGNrDe/hJnilJOdhlw5dyBar0l8jMyOk52XTDwfgG6rPjou3zmZLWByZQ+
DEpZmp4qEu+YIHJY6eDDBCmrd5hn5IlZ32ExNDVzErZ0Sedolq2yFf1SophXj7Z/
z+8bn1Ou0DBGJAu+zl33c7A1oJhqjdTXyUH2ncHHUmueNCrPlr93/p2HbjpPjc8O
tD50jV02C+1ufb3K+EkCgQ3Qiq+Np3avRIHI5OzOWg+LLZjZMpLOOoRejmw6Q7ST
IdIlfl8IY8Xkteh1J0seKcZlpr7JZP+jzd55jsPIaiQKv/H9tWZ/RUKMS0GLTxzU
iPKD2Vp0Kh5Dedm+aKeyneKi02Blyin7WOalmreMTP+vk0etQhx17pILXvHb4gTv
YglUZ4EV31ix9NJNs8BcMJg74akLpzMRx6MCjuOczbFaGBOmXfycZTlyqVll8IWb
n8c2wJVfRNTggloYTLMI6qV3BsGwvNGO/b4WiasTBcYKRm+iq1QDeIf/ZK9HeqkC
j1kekG0/RrjG8wuny4Lr8uIbDsXYyZHxRYIS9YGEXu6VeYKqzzjFSBnNEijzBBuQ
XavNRC4ESD99Jsd+mYGbUKKdUzGg8I6dGh96rW6A3rPYjNectUWRSJyrq9KTXVF3
aPKrjzghDsTZ0/rVXlLqP8RRZ542srSfIgc629hcUeWgTdQSJFZR4sfzj5m0MyR1
XzfsjdlafZhPumw8wBWnTkqNyvClQFgHC027f5vdDvxh63M5SqtHHv7X43fHxU89
7FrLUizzvqpll1LLc2uJ4ozQ5lA2QzD8m1iJXSxdYTzl8fesshYwY31Ldd8u7gth
RFcivXZK/yowTftAw6WVb8pFJaRTxKGATTy84gGhhcV6WBnbX4HPSBAY3M7ML4/N
3XNj0Lm13qBpvDvYyxSowhDC2BKUU+eCe4aPKoph99+UzGiEj7DNyJcfpljVZkNd
gF5otYzWSdxtKYkqMq0hTOQrLp4Nm3AVY+cCH5WcV3RUvFl5GnaSPcDaFsPLIgv2
znpd8UIY+DqfMsFPUYa+0rnN4ST1igx7WHnATuZbEXDezwWo0mzbzqg9+xMO5W8a
geuMM3VsM1CU1KV2duyBITlU38J+H4KAYjUpqmRyiK2PdqWWVwE5e47xHlOJD5/q
OfjJrgljrInfJZSN7GBte2oC5TVBzvTPbkwOuwxkmNJwnm6a6rbpJzEfBw8zJ5s2
gVVaXwpxcF6kY3uZw4YHVw1zPumL5ObFdAlc9ut0LK9m+vO4NAsLfGNUo3trLQWG
eD+puHDQtwb3U5DLqd6RNZV6gPFosqRcVu6JA92WGkYD4beQyby0jy3LVhLudXZV
Jy12QDHfnC5AghOFzflVxuCGam6i9pHlot+gHAsmmibq/zTM4vwecATPOOxdH1wK
5r2CFRbRWVs9W7dnjhXrOXwQHQZC2mB9DkBI3aT/UK3eIRbXBXUU+qO2oAog0441
RG4B7LCqXOhz1Ef/g3wpM/p3SDGd7h0LyY/7ypvrSSekkokQKLLZGBQkI7GKP7Dz
CVluK3pbz/OQu3rbTfdUL88rs01BS4FJNlPbjT1BDGII/QwUC9y+Uw5g9NIuXSOs
y2otBfdei41XkCbscxPRZhdhMXlB7elLin5jZonm+JVmYKp1kq2vw5YfLOh382Kc
kl6UblbKETZSt12Idqtf9B7MzinrKDpnXLN8gdWHdDDXTTlFuz3iDSS2k25g6UIw
6Ph1F6ziwEWUs1jK2gWovg49syt/wk6lDhGudYgcMQR4j+cfhe4PzNbcZgStjzi2
fSAZjnZ816buk8I5ayOEduvZC0sX531qUoKOyYmooOgA+nndX6jmtG+XGlAQ9N4p
Rwc4kHrHFfJD9vxJlKZvuY3XNX8zfifzuwOSeh/00vnnjS5tVmE0SuCoNcv4bJNb
BhLLmUSwFZqu4e7K8ZLK6cLdt/6uVKjnYUDo/R5bOPSHO8QcJlRtR8478pCNM6tz
czj5hj5KDbGfN8cJ1+rMimpbyTOJSx3BoeQTaClND5olL9SQs9bDBtiRyJciH9u1
wWglfPaVGKLwsJCN4NnThCBK9wIdKNcSU1g6nbKps8VghDXPQPmjzoci86/wrq2V
cL5PspBUPJroGS0DdtGARe6/Eepyvh359mw/pxEibswmMcZ6vbYQACPzLxlbUmZS
bGPhV4kqAwgLa4tpvwiwtEOG2l/1PTXueffucGaT3Gr3IkmfdErkvByNDszgm/yN
Py4laEkH3gCvMHXk1KbZSjOhEmFQ+1gqdjV9vE2MlZRq3xIkv6r9O35E/1Z0VwJI
3/oR55IZkS7LJjIUyslZKQUvqFG+8wFlMzD0DocdrXz0hFgXdB2SR/ZgVT9WkQ1c
zeB1EVZaRfm+Wiw7g4gTqsH3hRf8BVzyo4X/h9/Evy0VYG6HTflImtnXeJnBuZ/w
1X8UDg5hCPzI93RZptwLtf1lEoo8NT/j3l9h9mNpFmgjevVaqbwEPUj40cy8rMYb
BL74EbQ8Q+NArXMFNALCpWIWcj7tipGuPdJwyQ7zwlMVwCalQVrb0SqQsgl+4323
mgDfvUThvdKRU/mnjWbpFDQWruonNa33FuG9dg9fxlrXRhSzy+3xBHSaPY9BSfCn
MNvr69t5aHaz3bxcnDUKmYl+D5uaY9DrYbLFYCnWO+f+4QJ2GSyzknx9FPqVw1bB
fmGPWq+mHyG+Hwx2m6YTJ3Lsw/9y61Hxo+iHOzaqMvajOvp1mIcUZYtTn0bFUmFw
lBCh8Q7IiGo4hzvi1FAkqbRK5TG+QRfp+yMshuqDKY04YsyOEEDnmHfp4x0cbAT3
Wp/31Yd81WCcDRHch8DzEGAWGXbR72KtSeFgmyaq0aIMH9AGypKCSkr4tK1tU3DT
rfZyelrlJvZVbpL0Nw1SqzDUSykU6f0zl7TOW6En8hmH8rBgFzNbInrLPoKmXZ83
79hnXE2hZk0r0G25MOWYI20HtJD0LxuXCvko/sDbb+EuF8Rf+qxs45CaHO4dOcn3
t0A9Pjmmo7VdMjahkXzOmNTWFafl8d3erm1DengEnrvnA8v9jNvOlcfMEsszCBwx
xzYeQBImdihHgF19X7onMQA3wOFWAK+2hkgr0yWk7yQlpBuIRLUAwPJPuAj1fLkt
86xqmPA1HPQ+tRmojszBjfNYl5TqtU7QaYDcy4N6kgJcWTyQRasWQ3UETHmKSxDP
i6+POFLO4Zrroe6rZQ86aBD6pVlnJuN3P+FnjulSq67+aaUKTW2bYJWshzlPelkk
OjOVOScaRgeCHeA3IzbpglZQnmt9yFRIOfYEzPnkshOGq47f+oNX68k/DTEhYFLS
dP34MM1nbTyZnciW6mnSGgLtd8joQYtaXKJnpEpaba/sAkYowJq6fglIqTuv6mcy
Q/NJxz/vXjyXaS6LzJarApjjebF1FyPLS6qeg09K2Y7tIfHObK4+4YIJBXmYTXM4
kAI723EJpFfy7C4xa6iY7Uw/LVDKbLb7OBBMyw3Nt+k1vnlR874fwU1Q7EoCwG1J
ZQ3X6fHfzpa5nCgA1fLd5XoVDeCX+NLAcHPnGeKS0iZB5W8H4Uw7lO+wIZTFlUVD
WSz5X8q+KysW5ufHbalykjPIFBLMn7t53cYbHgYxOh8SSgRPvue5B8i+Tlc2ySAY
5VhmTx/SUSNx1oQq/unmfhyDrBrZ0LHOeEWQx4JJ9A1bmWih7/aEWwB4dX6fFU0r
g9jjNs7DPFtOqXZL4ul9rP457bn8Dd1/Uu2eTxb8FakIPaMmhfsJJ0p71lhza2vB
g2dbZztJtnXXJnIuPMARsRILdSZQEyMGsTciEpGtbF5V4OiVexX+/v2EazN6sV8h
1ytnltP2WNupHdL2QsgiDNMPvxhZq9F3XqnHlMEMUjt+yWqdurBzJsaLI0GylDXr
ecKw4pYeSjU4sApo5I24SoxXgI/AnnujQeM1Iti2fknX25KBYCyfgEGiDo1dUnpJ
rT1F+PzjW+OE8N5ySbvX+bsfi64iEddn1SQQNOw0IVysjsFnM5OMdg6FT+wMTxzO
zeDn7iVoMPyyKLz5CJQCiHci2Yp+Ivoz4+WBMFDuSRVqBTHHoRetxhNspnHs5C79
wvuLLe8ucR4Yg+CSg/ydO2FUxzcwnMV+O/dYpwv1w62UUZMMvFhny2wCitikcmyp
6IdrucEhL9sFfdk12konZsxSTCLVshCzSVnnfu/8G55RL+qvWEZQyHqaS0jjS25I
YIjbOTmy1EKPnXtb/cX5jpL2HYQKBa2ZGXJ2Bq+jRnApE5Ec2JKapwVBUgJKzE3e
b2fG/xWYxc+ZZC4a9DcS2z555eMDaC2dHiyIf6jc12h1Ba73fnw9BEFbq+YLSQmi
96sZD+X5BIuqjLRXJRcdfaF5I2YjnHv3haXYaw1KVqwxOj9Fc7CuxyWA6buJmz/w
6P589G80OWaVv6GnalVhLjT0NtUxwMxD6+ICrh/rDmSzc1KIT5hMiXGkGCdOggIS
nZoLAY28hBdY5NgP1xw1/CH/EkrdpEQXRtQueuJuBM0TVVqQqssapCunODBYKkPT
splApAiXz/CaKIMEbGQUBSGC05SSX0OktbsTNUc5L4qMUE9A9QDiHjdrsnQYmzqU
a8AQSW1N0JfJGaKsLP5q68NhZl9+3rewcpRWgfOYTudUPf/WCIkynsv7eVf6kaUP
n+LzF+yGTKCh/tg6MdDOyRNbtmfWhqJMNw+VKhoaSvcAdfQ5CZI4P8cV+dY7DyOM
cZPBVPzSbU9DDdYcQ9CuSA40Unrxzc9/MgNjeGmHoPI6bti22rXchNoLj4Zxkxj5
Bw4319yEgZTdzh10btTJYDw/rNgH9DjTxIh1TIE4XNoIGH5sxj61t4K6olXeVzWV
lCSGDhNYpC7aEayplEZ2VZ9VBOerxtpLd7MeM+m7E81y21JlLLEfIfHmrvuypQ6d
HK1bIXdql6hxuRmo/zSW/sDaElEfMq5NVwa23vUdEkWqYav/Jo6biSFMPnjqb9id
Uq+4uIPM/jGK8mQ0XttOTAJqjxPmoFhT5Jy9B22IbqgpFUqxO9ygbjFzt8jWLdk2
nWyZxXjAy9RpxC5O6zxboqtxjIqBt3dvuV1ZLm8Fb49N2h3jD4i98vYHRlro5h3c
1SIA+czSfrsW3ORAV3DdsKsMjQkr41Aw/qmmtYABOZy7+oQLjmOhQsFVmDAHSjZF
N0cCK17gZFzo6tjkX0nN13rL4Q/pfkaFLJxPZs+kjIZdUNDwcSHsiYZ5vkMoh3Wp
CsB2i/Y7nz6F27BrWZvVwAt/s9VmpF3V2KKc7jfsQyAmyMg8j4uDrcRAXsj5yCEX
sU2wVJgbmzlUFalcbnqsS6rVPSd2DdGwnrIpw6i3rC072cVJa20EQvm1WqAaFpZz
F8WgQlM2RiSOatxoES2ccI4/as2WIVqrCjgBcEROjttWTxYjDecUuXbcvTUb8qnY
vGZsngDdWKtN8pIyNtsVyQ51ho+x3U6KQzoUTs6XB79f5IxoD4B/+eAWHhBeZKPq
WPRJdRUZ6Aop3/KUnqyD1Vs1K+8hGFWNrcq0KPtlhDQCz+L/GgM+9WyS+INutfhK
4gFbzVkoSEIiISi365ZoePm+xfU5NH+ObodVWtHkxT1jMcVGK8CSBGzPyPI4whtd
GjEZo0HSTQxl62v2dtfpqGDmYMTHbuRXzAkpDZ0wlZkaVvB3KoDnpqUCfdDei+GP
TR/pLsn/9vx+HDuQjooj6zy2z+g2DrrhUNcHuR8dIqJDqPi++Ye9lniL33mXMy7O
qq6IS6b9nYlcnzwaVg5KP/VNHxzuPif5ubTAc/m7LOZMnlJIdJ49S1Vl+xxdfRxG
6oKgpYKk2Xj8eo/J9/8j9ZiPrXincLmWw6pG/zxUgjNTVkJfGC2uwbBKs5td0vN0
TDmkkUYooCkRBI8K+LRk9ZtEoGlezS1/pmcZnpZPGKxCLDbfoN0aeNeF0GZkqHIn
Uy336ovlO39WwlTYfQX1oUPijD6jn1xmZ3YEwQ1g2+G99GeZ40qgRVI/N6oVXda1
iwpzu8nKErKFeUDZOiR7073xMq+rlOShAyXwrtQ+rfJdyFuzgR3C7/yLhhEDDJwO
JKkHw18+yJ6SUb8g/hBtClfPGqELD0qGhbwlQS9p9bGV+tad06g9vIM7382XgL2J
kgpwYX8mG1zbx16bWztGPcDZdhOhrTikEd6tXJQMbKbaxLDcpdctOjlwZcBsJfzF
YLoomy/b1sBWqkqVAklR8tRxdFAzjlIcaEKVp4tb+pdLTBIzjk/HrtAH9YcKZnx0
DF5QXyQ37BFsBdEz7bmpuFngzFQzw7RaH6hWRq3cRCTRVfX3HcsEXmr8kbxP293G
JeOaDDoRsYAkF+GKJTSQDg3j/6i3ax3zeiTsS44L9+M0MUGYgW8tc0rJZZ2PMTZm
NtsEJ7ZcL0zP53oD5LkPJ4W+iR96XIhd6vewJBQNOnD+DVNoNwVqoLwcoxmLTvuu
0IHli+JbLnCtz9RtYpKdxV6YfXiYPbverT3aVAlA/R22qHuOg+7Pugzj2QL0XD2I
pM9GnT0MP24mdqQ0TwBSzYvR1HOPUpmnMt1s4dWtnYo2E3Ubr8sf4dsIwJ123K8r
wMjVGF0S3OdXQ2ByHtTJqIZcwP7dqzTlX+D2CNmVCMijCqSXp4BAnkf5rkBB7aK/
v2+HHtgYGTAWjepCYan2kBzCpZdhdaOXo+WeZzq+fGpqixg+BD2Vz1ntXpeV5qGC
0P6LYVcAEIoZjGCN25cO4NUFJJT/gnL29sh+5vW73KUhdZN3VdrSXMl9sMUg6OU5
dZe7mxgAFvCnnx6uzh9IwyTn7hjbmlmyJWgZb8c8iFK584VqasQVoMsEc9ok8liJ
hYEtZyx4EA8Ge8FXO1K6obydxGIf14qayDfEfJ+R1LVdubJw6yinEdFWiGFLGk3O
Be5gqnxA+LQuxNQDiac+9h7m+Hu501RrAIaqxPhIJlcIEmF2M4qN918r600eABKO
ROQP0XrOd95HfCPKob9N/ATqI3Q23dvc0t7V8l7jYgykr5DP+Z8NrW9kBLseQN5T
PVaM6407jP/yeUM110TsOCyxeQrZLl/5RYNOatt5ze3hL/3l8LyXMWi6JTpi0sL2
Zh/r3yHUA5thd7fsjLCOzTUR4pbglfQpQVCq7atopHv5zMRJaLw9m++7hUvQ4Bwn
+Cc8Wbc1uPVxJMvrrD5ZSErNJL386mufd5/WYSpb7mv1injIsJyNAdIENFpqUL4b
BkuibeEFtYYh6Zh2UslV1mh24NBg8KqrD2BP4S89lJHadjUHT+Ni1a6uyVE5b2Xj
KeAIJU+qos+tDhx2ip5XG94a5W42YWgDt7bkfBL7+/Fax5fOiOshQKgSou5A2q/I
lUjoJI4acVTIDnyKcyAE36Eu3lYiqu7ssW6H5qy+A+3qpy1WZ0/sfrEvMTtvRlmq
B8uAE43m4OI2CDClG9EdRiXbuaQW/RtSW3BdEw5Lkz7BQ2TcIfEbrGlfS5XfI9jn
o/qQfKR1w7T5CFG5zrYpv0jxFxo+rjCEppoQbT8Z5QaE+FIoLfpE9ssgwV3+iIBN
AL8n4janQah9pOHBtd+QCgyJYTOL1KzI2HC1DELILPFfiZSm7pjvOnu/ys0mS6rA
Pxe4fTvv5sj5C4gMZf2mGrbCoSSIshK81+7J6vv3bos3DErL/68KjOlhjaD06CSV
uvQxERbhAk/Ndj89CkyA45AHUUYKr/2/DdRJz8ekQnMScXXZpRhKd1mDXJCcrPmN
eOmWxlWSelDDamT9+Kl1m51Xp4bXUk5bkr0OmKgKZbsAAcFqo7KBAiNtOeJpOaOF
lR6M3A6OF0I/IY/hHrGeDsYvo+RdjkahISSGjyUeXAkrk7c5Pijgb0pxm+3nuO6r
D5YLU6SjalLoKg7PAkffkkRjYQHxO9NfCbBMPnsqRmVknn/r4qU8nqPzdOU6VyUn
1Kbq3il5RMdaxzgffqMD+JwmJ5tRTd4FUHjfm9mgiaOtNYjKeHuRUikSxAJireQ3
Y7ShoShcrpIjWgh0hWOKcJehysRTsuNkQ1Yr3/ObwOi1lkbKHcWfSm2B7WEY7qDQ
fqRQdeU80FrGdr1uahWy3DzuhBylhRjXbiuZEsz31mokTO8Dmtn72bZmfF0ecIm1
4R/lGIwT4sPTNOTmkQZUEWUBgmYSrILBUjI0E0E1CotHIdpZoSjWEQ74+Exxghbn
lAHls9kGLWKEBWjGtGH7UyX3jsYead2mFgJTMwOmus+y+Rta2n/Sh+vhm+aLIBtC
6DeXRFlFDcLGl9SdOPNhJAI9m0B7t+zNIBU8wiWj7L1NYYzwvz0/O4lQPEofSsR8
9iwU5EuMrVxjCJVRN0gMrr6Aryl7lP4noghRkg9Nx3/8oERr1Wlp3/n1BsSk2euh
uRJ4p9F45Z251j1ChlrPphgjgKxJAzkGmxEK7mIoYnMdKIFMOJrYLwdufk5nKzHu
69HvigFQAmRE9KaB2nBi5gqJwEZgcAL5puvlFChZBFrqze3xhioBp5/HgkoglCVs
dONIUCsHonvZQ5uP79opInWUoxpvBWGcYZEeRW/UCPhj8a0QQOeza6O42yKMX+Lv
AQc+FFCFTRcSZqdhztkuW+2sXfjYCoasYrvjHOoxelnwIzjOClg4GQ+yjdt5Spde
UHmb4QOM5Bui13rwWJSkyk64DZ5WDKn0rrBq0M066mxGaVk/zQvWedLwws7xZpd4
QzGnH45Dnmf2P3TMW9kAc1wkLmYRqsBxbAYNGgk/FApHIHJrJKOSYtVMNhQyYP6j
RqKUa0y1UB9dtD3swNeGQ16dyzp0n4OOcJ58fJ6ITDyX8py5usiuJkcAetYUyV1j
rNXMrKUk10qbYn3+vyN3k6hJwri3bfGjE0A0QtlH2XuBwSyToF3QEMFs6kFQ+z2C
UxorftwY6HZyVjIZtnGUPKLXFqEZjtyqjt/Mf7SPTTgNvZzQ32GuKGXenmdev8Zm
4dYZXDcpSgHiyBbWj8hWM0qAGn00Q1zsdfUzu402H1q3s6a0R9OaEa6dOIWtDm6L
xhRFJQC9PVRTcFCBGsV4kbGU36ynlmvxytBuuPqJgFiS8ioNLAAYjZpTaPWFiCpT
9ewwX/NQ5t+3QPNC96GW8NuDHMMYM3QvQnc16hWOuL0DoF1VZhqkcYgOET140ahF
QKM0cgW37XJyFscuJLmU1FHTypzUwjSt4V4ZWimgNaFxjtNdJ+brIykYnFnlAQ98
n1jUG6elFKOZ2AeYUIFO9HLzIWhpzpmPpVg2kt/rdfYV39oahFs2zKxHl4RLcU1j
WQWPwicxZ3JeICmI5e4sA5m/z0FVE+bq9fa1FH0i6v1OL2wC26Ly5NVq2pdaVyUJ
UJbffj3w48HuSRweYEyo590dkeF9AsR5m30a+9+bAVFiVJUQ4p1OR5Gy5lVAdKO7
mIKcUi2gKa8E08q6lg5zDE0f5frNKfLB2OklU0ZxcN1AsygtZE2ILNizKL/v6xub
GtDpMDI8RyKWDX86Mt/Yw876x4evwwvm9V+q7jUrMVCGZx2KEW7olPgXR5gbpL3S
K0/ULxRq64UKhhvoftYlpmtPpWnmI7Wei9f5joV1VVp68M524brhKmTsWpwxePAB
u6Orork5fkjCwcW1d8kH/1M9qgrWMu0BI65boP16Klpwsvx/1fBe1RKijkX+hQO2
qyrmHargQcUSFYT44RZIsexpD4S5zGVLWgx2B+Wfs7UlQeyKr4l+Og28YfbtO8Q0
k1jg+yLAa5IAWyk7xW8YYnsESdoaGRKT9gNBYlcC26QtmKQUHDG+/0iLJ21/a/bR
uAgUVUMmon6SYa0Pvxa9lySm8cdQEf/pSBGFKcsLUjKlSwEPECdI+JuLtA/dj5/M
3wrqhyS9/pQKwUr7u2qicizvXBewdmIYQPqgCx6IsTvupLb2v4u3NHnT2Na6y9oe
VeMMdR5QpXKGt2aKRMMb0VI5YHGhXbIjLS+c3le3YVb8BfrdF7rFbLGJgDAvC46a
8XSSF9zZQUMzIUDPAxBB73RDGV2GCSEmlw/5WnJkS8wsp7BYb3tjZiGjhizMSGGH
kXrtjKMSYomSFE3Gr0nzm4v6+ne5waotReNFxJJ80tMlYhae2jUOlNZ2DmDEElmd
/Ee+/27I6ojNiKUG0SqDE3S/Rr6s0Es37hZMyeksVtOSDVecGtOYUcHJv7QZFBZg
w3yG4v4/V75nXKzQ6uOhu1FrS9T75wUtkNeX55dx4LK7tbBQrjfPTO7qhYNeeaoS
YTFNa4OfAqhHFYrhRYf+jdr3NQpdCoOZ3bqLQY9QfkbvRgPdq4gfzzQyKR/Aqlm1
YPrTfpVp7CCCLp5rLLNq/tzdm6bMk4cSeVD4ZhatCTW373cPIl0cvARm54NOpf8W
KgnURcYBqzEC8MX3fK1ZUCbEWyzOL5epsaSzLN5+Haz87SFOkrO3rQ0QKki6tl8u
PBTt9SAYUUvPiTkW4Xi1i34CRSoUDqQOCM/tXPeVX03ZM2O1+0MfdLYft8hL6abP
WHlleB0pel7nsltofFErKYYnZUXiZkCLyLhZ+0eY8ko4fxk02QblIW6+VC7ZFHE8
0B2yElWO9zgD3fB//eQQfFysOsrOhmQSrw4Ai1v3CgbdNGaHyJb9tUaM0rPpUXR2
TXjqo2auson95D1nypysO8LLflmoXFRBYat0Cd22boGdDj4iwzgZDXA77lTUTxcp
wzxv6QdYxPfXRpIVgZIGLYUlYyLUtXImWpzA1Df2Xzs0YpaccB3f1Lk33eP8Ftbn
P519xqBtVtZrWMQqX620uk5WEiECmf+MMxUGkLfvjDKKayY9KC999ucGtXjpkroV
TwtaVj93SUbxViTJvp058MGC18eum7lxAnEJ5/33Wv+TXfo+EMS30H5nEFg1sNni
P9XIsgAvxAB3EsZkhYiUpfnEdDFUpiSlnIyfLgTiLsPbXLzTC7yqDtayXr+fZJ+U
luKssmqzZ+AYPqmZVHUGNXi9FL3j/uh/2HZROwhB5TVkAO8RJogdtF9vpcm8wuYo
2FZCo16fsT/tqODUL18HZj5ADyUadad4MHIfI3dHrGCdRg/5pbWjKAWyl7TDqJ0r
xoJMiSu+n1qE9mctQGP9Kv6jOFFeI+dFrI07qAWVm8S4MCN2ipvo3n1AXjjtGeEE
23K/AVVlDiT2XYDsxCFXd1NEpyaigWtB+2nOU5h6XyFgwOLBPKxAhs6Yk9jL1KY1
v7oHhilf6NSQoHQd8sc4Mx2EAmrpRZAkcaUOYhA6WE3/l2jEL6nRzi37/rKMYTl8
I34dMm7+HzUk475oGh9XfyhbY0egygRFf3NUcsMe5129dMazBKdeEMxPdzxkOMAV
DlIKl6tIHRqYvJlnJoSDD5vkJhY1m9Ic8udBPk84b6pfYnH7TZZktWUtsNyOl6Mc
htFBUoONwRg2ElwX2RT+0R+L99+E7HcxftbvUATNZ/V/aSY51tr1daT7WmOyk1cH
Bb7WGIVJRgacpYMvd47H86Ek9ZJnrbQ4zRzlGUQb//mbb7f2Pwva2NDRhE9s855l
cLSceeGwYsZ0af5yxeezaIuWYRV/czQ3NqOZKpWLQuDZYWHKxQKzabHUuXDD7ofE
iNOs3kPqWazHn+J/K9Fmco/gEwPWXHdo16LuYEd1k8EsYkcki9bnUGLvnLvFn+YR
XS/UU2JzDYtQACvvUuNKVyQmZwODU1N8l6AvBg2Y8fV/gu6ouUlZ4qxUAuxKhrNO
mfzz52q2FLUFNUdIeeq/0n6We11d1ZRDkLBWAjUznNqprZbl9HhrMPZ2dpjbA1DM
NX4e7Kk8SyDOyw2feBGNQ+VLY+CAsPn7NbEPFBQ8qOcxw3DeT7TdxJNv2uc3cKlB
bCyr94qDVAsDuFPZAfunKGyN2WRoj0o6aEDfCQXGniLQk275HSccXQZPGrgD2q2O
DRr6XZaQwtNLxgBizCFw6YdCqfsoyurJCcqv+WYhpsHlplPbv+FbFZtkO5EBv4Ej
Et6FybN7lQruaoPX+gekBRsd81FpYjH/ATkTAHR4zpoDwMyJgEiTLSn05i2j+nAi
AAzlYIJKJA5DbEabEdGhzQB2FUHD8NzB8pIMM1HCioF1z3WwDqH0Z/aUGJZeVwE6
kcI+MrJ/aP6rRTOxPL193jmt+3CbgnEDnzuQS9CUhcEGvd4RhUFp4qRH/H9WCvl0
xSIR3lynhG9T1Zzby4KNI4hWbEHEraraVFu5EF+NFH/EYNqDAetC3Dn0O7MGv/IR
VvV4jezYdwkSqtF0M21D7fQrUJ/VJX2BfhIktSsh3h7xd18PBVkHTFYMRR0VgIM2
Og6kY/D8qk8Xt7xSadrvsNiCNLIhXhyaqdEAUWw63piSoM28KS32tQO54H26+CdK
rtkdUaJa13T+1inMPOw4PThObrN0Ws/mS6hkpjx0S+YMYx/IIarDc5ekUyzKRrLr
gAqRtNS1Dp4ZzN91hsc95mBap/uhZy78x1b4mcAtQV1G3k/F+xlnllMoOHvOt+4F
ojd1PIOjO3Q5MFsWkXbjITkIUdGftFS3xKyuh+WH4iN/lGzAnw2fRmghDX4KA3oG
jMyhjRV4HGN0XVkAGUqOB+1BNLMUA7ekz1umPMRQg6YtOkAsnfRyABonwcBVUN8F
8Ux8CKXyVbgnRFmm3gfMDPzUHYT4L/Hg8hQNWBVSwoKllobN4RhR6Gr85a1ZefiV
251o9oqeEFB48LKBl7TgVOA/9XCdurwJ/WxPOpfM8Z7X3b963nRdckd7qi/TbCim
AtzQc/NqSXBKpcK4sV1n76JWfosUjZvfbP/aWcOakTiPoQ6fJbYcYGHl6HdPaGHI
5XPNUBrdCM1BsRxmdLwagr+CibU0NfyvAOoHN7hbEAnxkMiNsVMs1lHZ5kjqve+C
0/90TnELGZhMNIHm5Q0h4lHOSnw0C6Lw/M6N7qpaWgtUUrY4CSOxCYAjg3D2Fwd+
/Lnx0YaNr3Hza1r1ONmTuIXRWI1dyoC5cmCqEypFDGXyunF4ZUvefo+CPJHpUz/4
uyJJ+pt5KLqQwLN8uy50uKkYF4Tw230rMBWa3M/vgFzFQeb9WpAytmEX5Xm4vDrN
cWMSMJsdIHwh6u0OCGROZ2UQLBQ5tuhl+HJz9bEm119HO6HGvVm2tH46/i3bpZXf
VOe/AZi6R6LNiS9VDu1oaPoOY2f9ScPdKD28cgBianGq6gERgg+oPix6S0IR2Slr
P4W7OGPG65F4MknaS2uKOwDOg2l38qgqyRSWqdC5DRgaHZlpRGbsxvlRr0HMATSt
kfji/et0h6mQFi1NhCMSJPG1rzyTtd49idaZ9nUNRJA0jskhA2MgXWjQT0RTDULj
uvaqvje9KjY4oz2W4sVbKdVLcgMHP3KdfvnY32uCnKny1iRTIQEmeUtMC0NDjbCx
bnmxsRpxnwrq98hpwf/W8Ly7C2Qk0qX/d0Jw1FKXsAMMQN9p+XjEMw5ktuwIlVK7
pTsiqeMumdqNgDIjkWCS/zEg36B0FDodjye7VWea+yzeH8giQbC3sE3tA6JwrUBV
z0Lxqkftgwi4uzoQXVBANcYRtWtzsyvWz6hmsdV00xTyxksFl8NvPpdHHAfu4MHn
/uPzF94kw4lMksPYvXsdYqijLI9rh2GARxTM0hUgNhNUBWP0myd43sUhFARkMOhW
Hodo8lia9HJOKpVwmnd0nP7+/HMRN19X8o9p66DL34zGI9TD0YPk7s5SwdTlb/TY
SzyFbCweAY6V1z/jpcSa85aPA5sNGOHhOwdMlYuaojp/zNYvdr2T1QDhIy/7ZgnC
y1f8Vc5cb3z5mNXmfMIqRUIDTHkTV/FZh89q4DVd+/DVLfWvG8EB5tc99JhX3oVF
unJB7Y4vthCggGnVUgOyuv/W+dgqGmU42it5A12wYgGN2zQ5wkEn8/PuanMMGSaH
K2Qqpl99PmgfCM6NTPRBrj6oTJZ1wKpga7JLVSIxZ9E1PUSeN60SmUz+xEFV03tL
x/EhmpE980meqqDgdyt/GtGnfjdsHqETLrCSVkHecm0P0Ko6qHKDLPtldYTxTpmP
jBzCs54Dh5/9WTxNxrTowy3VjAVi5ZRL8QqzX09tiyIbVAkJGbPtk/v6Xd6ZQOqy
k0ffQZXr3caqSrvU6R7A4KW6dTIfgsN1T3yznVOKSBSSPROTo8ZTVBhq0sp/uo3F
BsisvjUc8CN7zbk93ZAsh6mGrrD7b/mD3d46r/Q/u4b6mPAPutavo+hxAJmzNGIj
rozajVdFsu+fFQt+TeKEwfx0p83a28U3385cTFeWOXLXmaX188fd8EU3cGrC54BZ
yh3Z9tegN3jK9Grzdg+LzOlXFzdBlf6YrxE8OtsDNqO9jRmgPcUk/SxGE5Bi58/G
1hkBGE8YCr5063NsmQRN+bZ+6Ikpdg4M9RX5tPDv318crsCCdLtOv1f0MUHGpCSQ
/Af6qSNY8acusftq6Y1Hmq4nnQOddrjfora7y9LRNPJTKZSMcDUkUM5kgUgfGkLw
bkWa3zZvw4jhWeiRJiJPwfE5iMaxPqHAuP8u3YKo8T+xXelbzt+IND5LYSW942oi
bQG78qp9B0gysIa8jZZqiqQAoMSegeKctwaHdmfHRhOgwUVARo4AM9oIFoGZMwxT
LkOMto8o5v+eImuMxfBFBgXG7bFgQrkL6Aq6zFxFl/JRisow0sxYIP6ex3V1e82M
pctmbBOpNRaf598xa+S/90dqyqeqYC0jXREgsOnCH7nzeXN0L5hFYMYO5q/GdtZs
OxHP3ipZINdJqqkXfT/I/WoCyWGKHVWRukyR/zzvc5BS1BLH3Eht2d8vQhpDClaM
6zTIxISMJAGaLZiTHnxNOwgOSjtuAt9Pnnm/q1U+ahsIZXv0wlfIgrVLMCZAJzlP
mZHxZ+nIaGnIvLcfX8nI5qEboXcAUXCkVapMHTYiXFSH5hTmtUWakbNGHHGb8ss4
O18EwhqVrZx1ouRnAnorG6dVsHW4YhWPmwnC4eN5abdBKXgikXO5x/Gczpql0fnf
ETzb1Qhp3hRbFVyScnHRyrj6mLDvtTbssJA1MlmPo2Y+vIjCPwRcAGjIScliL8iN
f2fIrDQNgLoWA5O7mHthOqLQV9mAjPxWUn2pOjVq0oJ1NFteu3L2VvJtJu8ioDUL
TF2PoOsBjS1sDJD/XAiKh43GckqOgISDVTGmiTOb2zveraP94yLWirvNs/QUHXt6
VwunoSPoSlT42SZFfgwGqhCnEgPuf15irq51ff48dKBuVZ8yERlpgqwpGFf1bmvE
L4mZaFOyGvpv0yD2QAJ9ULeorbqq4Welkuqj0JjKAkM3LbZBiyvCqEfZhcLBXG6+
FSHr2wFa4OP+edR5fqTpZKPfbWIT3vnobPds88W/kRRAoteb3yyMFLuQrpE4i3Pp
pbRwL1hHOdCpLS2mZpx/Bzu+BEYuRqCDB66aZj+I/XVezTgnOuNJ6QKr+ETb51ko
hy+Pwf2F8tFBIW/fWBZDnnvvzvPpYOvsTESbwowUECV50SeGS+eeUbHg6uDEHpHu
wH12ROyEIb9sXjd/VyutQNAEc7uXkPrl6Z99LSwi1QAHQN7fKQ4Zn/5Pt6QzLhXR
aq2gTBXBdQSjEfr6g2PiiNjOBGLdls8jc71WexPlTS/ANvcu1Y0lgWWUQgI1UIzg
P5F8BtGC4IMLR03ZgXolPgBb75LxKYKy4+QufK+pyh1j7rjTp6UKjHx3ZeRqW4lj
FqQeWNfyjq3MftlnJeH/5NbfD1H4JiQDMuzowLrWsM6L2A6shjbRIGvBQhNKPswS
dgX0ifuIlgK2dZEOj5XwWIOt3EHwn3QBUwkaPZ1X6OUao05x2Kg8+05fdJZdnMaF
3K8uZ5c7iWUWSUHm4rPZoOxX8NQzaQFxCyFJ47XzVpXtqLhGDV6BK0fDi6VogMjL
S4BTEAb1r1iB0QScH3Rq/Vi+i+BkmpCgsB+8FVUZnKhlqrAWIn2+RX1Q65AbUGBp
3NZv9JVFH1W4vaRqIWFCdjfera5cRWcO+14QuZ0ksrjS+Ce53Ea3DxM1lBhmZ+5u
Qs/FFyMPF3nePXxG9i5k+HUVJCTUh7CsZHoTm9sbAVATDsF6nOlXc8UI6FbQ+dJu
H6i4i1Zl0ngVNcDgF0o8aDvy+RV9o6PgN6eEsHkRf6XrNWpvq2qaJUIXstyjlLQy
wpqL1B6nu3cIx/SL+aKIfjFH3/jAOQk1Tl/zl/T6GEP91ZGc97/FQ0bT3OdxQmjP
uQwGFQDffOTE8dhE19DEg8CTC+cPc0wkyhiT2ZkBaIlwjzImQaEU2dfLEx86wjOy
dqyKmewx2CooLFNu6DHXAgd2ZUBysUu0UgPiOdVKtOzCSrzKarFL0Fd/L6OFBZmW
/LlVJbkCDMPV0ctNU7SN0QgXJ3vFxltEb36gNOFO6uQTVwGV159AIVwjks62Lvyh
RLk7u3zsXXW3JEyHfumcDZhpQnjhZXVNxw3E2BQKuhI71WjFbKdbonDiPbSLYPe5
qVaZKiFnpxew8xo/U/+VRd2SXa3X4yjOGhOg2QexRSk6sCZgh5uj/xkVGmUFojjs
a2dU9R7S0XVckqeAcwIN5CrUSF28t8JxoMfnbk4UnlhNwNAFORN//hiXlITJH+UH
kpJ9CQlkWGvXEqnkBgbmVz6dfUTaWeBIS+imFF+b+7EIna/spw7OlvNbi4MulDkD
+y7fiBcvutRDdsyLnmhJ2RUuNED/eQNc0Qb2BAomrdYP2ac1u9mYTCUFXlYz+DDM
FpWho0DP5TiKMEgqYRMWC/gdZdRL7GjLcGZBWG3/WO5rMzxmK0Zu188+FGLn31sp
wYTR8W3WdO9SEqAR3R5d50mDijIRROHIX5m4PnzuQRxtbbPhfdrF1drGkq+UTVtW
U2FDGMXTHuS7Kbt/lfCEDKCv2DxYOUhbwH86UUg0XbtL1xJT9VztwelP1nL0wd/6
H10AhkGQwkHWefba2iCtBYX1OVZcN+uE7GkO+Ie1/zRYNEVpN0bMQV/FLHIezKdg
GMuQxpGKf/mTGhfallmwl/b3rDxGPBBk5XKTZQ8HkHECnmrHYf/9OvPQJIVIjePx
XHpDafcSY52oKihgWgUUS68RgSPRU4OoxmFN77a5H3JzMBCTwKafoBa7Il3gfwq3
p0jXefiXyPojRGfGYtvMQlzWrGOv6x6FRhtTpeIoNff88L45/pEL86H3uhHjDwqh
QSHR5ZR3D2aYdmrToIbmoi+IVrVq1dJ00jUSyIF30rRv+pwuACwp+5IAQeiKJN5v
M1uJwVp4tRANsrp60/SkYbDY9WJ6C7vxohdvVrACiNssbNiCWWbBWTVUBKzGvzid
koauoIurub8rIrQKaj7pdDVRevMHWmB9FIWjSLC7C0FOBYPO7R8WZV59ONuUrfcQ
IKqStJ3mjIdiibkhIGLwhsT/rQ8B6+yCWZiObxOIXAVT7QDlZGGGN0FpxeP843Ak
Y7t5JdcvS2luiM+B8jGnGqccEq9xC/hMqcjHdE/Cgk7+l0hexwcUxR92+E28FbBi
UnyEYROXwu/blNVZV0wx1pbe5FhsYawYj8UfrMMqJSf7evkt83eWonN50jIyqNQk
ZtmXnj8OA8MWsLbadYpzwQq7KT8fEufWn4ioRIRBs1jUZyj1IjBnlhgNuO0//WCE
WOHGg5gXufInCNb7q3p+S9hEJznjUJDnNW+ntrtqxoIrjiYZydP1aklWvLmAHhvI
UfkKmrl0mHNulIw9VvPZWYwZT9+hKFS0TLkaLrYtXujrSZWnPEP23kAS18VXwDtV
ZV2cxNvmyWAqdFqZWVqh4ZCExIHynJRF9+kcwH3KXow8SntBGhkQIbMm+sE+etN0
9pTrHBZbxql+kVvQ4aOc3GNa2O1upYQbmky8Xn5JSGQfnuclGrCEpl+xuH2+2li6
19cQzJZ0El7KE7p7P6eWsa53aW89fLk9hJwflHIHud+CMvgwo0kw0EvIc/N0tiIm
YzE2g2WcKCnf+k2zCdqeWRiFQlduujfDrW1koTQS3rEIBqbv/Gwj1rpb9WuLLAjY
QtjyE/aF/mVqPh2t2F2vxrA2U4w4XcgUe8vHGd7TnSqVCz2rKjWw9FZ8uu4Y532H
zdYVIVmIpKe+FO7Lsirjo7f+48uhjzS7HJYolpI9BXYaiOoaZF150GFE/7f3vNrv
rt3bRsnEzDrPFejZCnQIPjU8L0b2Io0RIpba/OhsorsVhA/ma+4AZbs/fHzOiUZS
yrzQY68bK6TV1rb4MEGEMBXSWR8Gm0nhKkfJIKtSA3MDyJWZyz9u1COsP1u222B1
UwakuTqB1+AYiHSOe8kDsjWmOskk8aij0ej+5O4j01tC/BSiJjHYd5Oupxn3kPf2
Dd7lMtbLO3UxOsTQpfyggkGuNZq8lmFPxwVFkp42Ty9uQ+hR9aDDp8p9QwAqjH1K
TCRD1IGV16/P1O56LRI62qRbxirPmAVdqM72/lnnrH7HtdjW7JwzK1V4TcTqFTBW
dx7/+T9h5t4thNX7IteXDXh7NcY2y93oKaS+Wfw5/Z4ZRWoU3QDDIym5yrglLArB
i058c5SrfXXbcLmx480esKuM3HYNGa/wzM10zKb4V/ApQKpUJDd5dVSFy5pr7NoW
hdWY2MTR2oY3HxpoKqPEy180NwN3xh5jXAJ9eYFsqVxwxzdO+klvfhSrBI2x1zAm
pasBON2A+VNmCdslpt37rZbz2CK83h7MjJGp2SmVMwiwg/mUHjDFQ19BoPjYZARa
q7GvqJpgErbKtmlqBlMeKbjT8lb+LZQ1SFMik7waER2xamLGdc/RbZctXUL7d1DN
0MUZfd0QCzjkN1GZ/mpYJPb6Qryiwyr9tPjRxLazPuj3O4P5McDerj9tOjVPwetG
w1FY+wPsTfdBVhNcwmUPgNg5ru4hAJEvTVuFc0g/2AzvrE7TugDpwluaYCV8Rc3E
aoi6T7R/gBaekBal4QB8bLYE9oKROeVu52mmRdXN0oDWAXeFV3daPjRuSeoDdsHH
ivI/WdYdgBaMuGQe4XO98cwtPYlm79nv8BCkFZbldYgX1fZD2jSCDyLD58Fr/OKn
SzMFj6GXng0vj86PkFLDXU1CXBrWO4o83iswqaUgDljJ4hLNmijr6WEuXnoM6JvB
OCzgQNBXRQu3His+6kCeQYOe51deTKB1w63e9FUtZQ1/za1czCdjA9Z6KgX9qLUg
VbN7C9Urjiq+16QBBYRnMym2szl/FSvu6m3UzMmjTUohzykHCCNo3qTFm/fRaRO5
wf7ulqgmhbT9ttlk+Gq99jOd9X1BAVk6UU+wNq1U8ITvAJgMZRyhbfClHVCa9eTS
CsGOS7doxDa2s7MvlKIZjjqMyV0iWfkZoTLhYzxcSo8mLwnphTEhr0k+RBB+KzOy
jDilfmN4tf2RPQJAzlTFSjr5N+MDbgEHw2jcJDCoyibzRLHcFDgDJevkrr8EhBfZ
geVtyXTnqXq/EedDXBX7bS/GbarF6xWC+lM3P2sAcYxNhuORvY3h/efe3rpnepLA
+2b5oaQtJjkJmSHAl5g70yXG54+3b1rqSZ8wUaH8MgoHZF9+Bly6sXorudYLTu21
QWYYw0/3CQb1C/TTs4QEIyDa6yQRlMGBYwRqVsIPHP3+tU27MVX0+5KwWY2aOl42
0Ik9xY87M8qvOp1L2WVv1TkiMu4ZrkhrLuT+QXlAt9bEx1haHhpVc8RNAgSNML9b
4qC+hOdHU4vJQBrxDf4VfH9I/kpfuxK71Cc50deUvttZl7xAayZZ5wahKShJcE5z
kF0jFmPxyXgf31s7idclkZGSAQD9Q55RDKsRhsdxDvLXEa7+pwQ+UmHNMwPbZca0
VYUOAvq3lbWcypIVkPPiWyO3MZwlrRX6t4Wj95lROlparrk5/Be6t8gONrPuhO4t
IV0Gmke8XSDgMhqb13bODczUUygq2e+TaGtnFiiKwJqKsmOlMX42CWqnBrRwNS78
kw3qfGPF8gne/VAksf2DCZXFGxGGTAZFmmmO9fc1lPcx245cxCUmdp+VoSwVWV9r
B5eEO0WL9NirEcbj6dwxO14evAx2gMMyUiLpaWv5O0DEvVrHJDwr8D+eDLJI/vgZ
4y998I8/ci635p+cnbdm15/MqrK/7rJQSY04mGN+zHagp7kSb2pc+YIQ3QlpYbAM
tGOSmVEf5AVsu5fL1CmMFwHwTbvWUAHuCLqbXQxUr8T0giaIrZJSXanF+Ek1bPdz
eQbkOIAt3EHRxUxu27S+rYt1NcDR0frHlv5x+CpdlaXxeFKok07yUxaY0z9SWdVk
emdnw5C+imQHv31JWhqmxt3bCZg7KgI853v49RzULuCqPOMGBqndVCDKy3++iipd
wHXxkBJ6hmN74z55FjwplxNJL5uIV4QiJTmtKN74U3PKSZodEzaNEIbvlt7kX/+V
Ed8vYLxrNM8GKgCynChNIxTz3k4IRk9kTNGFU7HoO6fqI4NoPCK2eq4bCYI4yGui
op0KoNyfVt+df4S6vmOBUqQzXUNppWUgjOw0+dJpczCzJX+WM06+8h2aoNr8f0ze
G7vt5yyaq/JG26YQ4bvFpKewv2Fs14JjiAfF1TVXsVwGTpRsCO/NjuU6ZOfhJ3TU
X5z2OvyX5DyA8MolorG7+4WPUoe+y+dfYfpbYRzaP/erF4SthPgF4U+YnmnMw0U+
/PoqUwPaRU95NH/oUFNDMIN9nJKK6P6yU4jCpDcH+Ea/IO9jpFuGbRlVt+7Un0wr
meIKjUHeYp/c+5PCLba0m2iELD1q8FUeSU9CNjyGLAf6DvwVBolV1pZjJkMhCBtC
nvDGCdPppJs5f11uYiQ469n25I8ZR5smD7bBQVd1CYvxpinlDxlhW/P+CdSMVc3W
MRUSbCnep4s9tyhzgKKVqEgUnn6U80ixOsOrfh9EKxbMlA1D1yPiPGBcaw9lyaxJ
SFGQ2y+y9FFqWhHTWS6uoNUpKflPCK0/yXGc2UcQ8PE7wzyCTcD5t4chaKqjQPN9
BuiMHyKNYPl1wixPSfUoXLgNFSIKv5VufOpxFEcaxIvC6vUwkkJ35kmgz0pVGQaI
RrkjbcWRJReMYKIQgiqlVIMjmBNZUffsjWeXXBNmdUm5W14EI261eMWJQfF8ph97
Ye/GPflEv8CKOCWfwSmOj/H45E5iPlK2g9z+OQlF8Zbwucm9StJDXz7AlXwUKofn
Jt8et8eMAsDgJ0bUE1oyP4+prJjVLloMvX0Fuh7UV8fqWfgiVXhCzm6tkmC3B7Uo
gh5aMmoefyvkN+Fglbgi4YeonMdb/z3icaUEcuWUddsJl/16QWOm2Z/IfT/Hr1BC
rQmOrgI5Vv2yN96JOZ4Fog7x/A6Ajl0Zbzoc4ElHDuKtfmC+RjsbnsJnUZYKxIwO
bZI5eXR5Ts0EXaUYpe/dmEUfz4z3XDCHT87eQk/Stk0sxhI8IAJkPvOw8/1sFdQk
id3FFnyyF6aiuxFORisAU6Qp4DnLgH46XfRqDqpmpdkr9NSQ10ZEJseAh+p7lrCS
Ybvo39YAuAf/XjeFVkTttMi0LrQVhbujz6ICT/sBxGEfUlZKmPdhVXKmikmFkFAa
+JYkPizlL8JE+B7F+s7M5DB1veXc3cdwFDPNaqmuxTe81Py8N1f69gj3fTVeHXJ4
N/wlnHCj08L7WBZXyXyIto6gq/lhelI8YZ46/qnsWGYYcDmS2FB3yAY4ye8xvNkM
kxgl/SLAcuJIpMOYmZmwMjmDofKKfY3QcuH9ViO77Zu89RzsuA/oXAhzvbnp8YWS
lIqu9ZN5E1Xlkk7AUWi0F5e1Ao67YGIucDeflrMJ8uXd/CQglY5EqVCbGn/A2Eua
8qQsF82mtnchjZ6ULg/MVt57TtiAkGriOFuowk+j5sRBTMMu74AXkNzpiemMnzc3
bqxADXEjYxAs1g/XzTb9dZae5nbBBLNKgrKfED5pBIqOB7AZQv3wmLAZlqYceZjy
G7b4ofzxVxDFlI77u4CWZ1AnLqfU/520qFCuKsfRGvbMZMJ5ZbPKB99Cqan3u7Ut
WyGn7q+u4Y+QpuKBAvjzRuFaCZ1GuhNInf+AHrD9kTIim5mZDDMUGF1JHH5pcNHF
J25DB2yyYPVQKHSQ0LTf1nqEQW/r4PZqtiupqoBNhFDDyzSEm+JTgEJl5daOr2Ua
ytk63UJ7Tc3RM5r+n6hR1w==
`pragma protect end_protected
