// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:13 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U6Z4SJboNZjz6xWowDpn4yHsQNqMRwdsHvBXXaPf4NqRTlRPcsVXy+rrS+kwoKGB
+WLInxRj+Cb1S1Q1ERVqg/6Obp0HDTxoCwXLRfDMSV7UQ/7A/2NHoHfx+VvuUmw8
wDTYQutQyy1rorgEdxj1WTfMK7u2BvsPjKsq3govUHA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13536)
Ki8A2ZuJlgt0PErkXOf4y6TomJCg32oZPUijSp0VNXyPGUzYG9kI5YhdnzOXIuBQ
ta8R150ZSxQiMv0f94wyCjma1eXtpX7gPv169k3jVRJWOjnnhkbDFErdtI1PTVUK
FTsTvjlZPqWs7khi8DZbFT0IG8wOjOf21hKeXgK0VYs8Yl/G1UjGHVEzfjakb72j
4ujFlx1pYxqzRnXWRtXC21Gz5YvYDB6fZK4ltJPqCB2qTlzu8CHBWSuXVCMf9MRN
fyrz+wmGsBTADG4izHY07KjQFPALhWLEMVIy79duFB1tcUOyM398d/ppOTIWmFZP
G9VNndiwQklKwoMCWukdyZvZd4WNF47hVdJ7GVQvhmpn9bhgXcxnmUMxNFTtz2T4
y4l+qMQmYTH1ufNQHI3EaIjmAQ2c0bhMT1417wgf5nYZFkilU5+cNrKo23u+BcIT
LYgsk6v4gwWmWTujK8a4UL/zF5bKsj2COfrxlQBkNPrjxYRJwRhLmgOhixc/xhCm
DwKhdio9W5doIs4pdPtDPQD4lWj9/55zs3CRWNosS4QKfEmsoJDVrXFWuhikFURI
To1tZeikgat8EPlt3HdfoWURPrHCQZm7VzCW6BktpOhJ0BwZRs4TsarD4vIUk/E3
fWRlTUNb94LQb0YMyvxfJrHoGkfKhuCvKYuoBLmEtTMdz3z2tG0aWN0NTeqfn8zo
FzNDUAfiaoKIC6ftHjn8TPGg0RRU5vEQgm4pI8SeF0k4ScPxzkQiWVUQ2er0sv5z
GT3UV1YF/tE3KZbX37eS1G6GgxiPEi4MlEX/3e355wLSuVd2OzwegJbZKHHyVZsL
dzULmaMEJ/sNeFsgL5GxtU4PMxjLDFJBncMsLAfO6uaQa8oMvmPaF3nKIuiDi13M
ptnQRLhaTNWJhbO5lTaD1VKcweBnlacRA+/bi/QVxxoQwT4P/y8vsTn0zQJPaUYK
CsXm7GXwowvzFhL0mEqDOqZaWrte7kR7p0dDwY1Sjh4FagkwhgSZR/+FVMYLyVnh
5vbDq63eXLx4bQ4nnlh1/yCXatlx/dN4p5fms03Vkvq5taolLp2QULlKD8vIjl8E
uPQO7kqlEJXalAEvZh2WQdH85k00Bry3SH2ni9+7j8w7/zBpE+/WAM851USkhkiJ
zunkn2IYRi9ubasYwWua2OkgPYZiP+q6OaAFKVxM4Nmam0f3aQW+1c5t5vDZrmFd
I9G5m89Lsgr22VC7EZ0DSMnu532M3nIquG6tYeE3MBq6l7fHe1nt4croLHK3bgPw
loIKynmWLvAbrOhOiVQiTpOX9MiHR44nLs5fqEdDhxPVCyc/fxBymAR+a+N8rpEs
3FeVFbyXV5TM2yt2w+EJo6QDzoAnGR6AxM6trOx4A/RbtculVJhXJy8T5ay1dBNn
B0ZDbWXjsbhmRNGCXI5H1Coj/vtZNndDx+a8+Dhy1x+i9z6xUJ9K3uM5JhP6ub6L
DkVpHeW5UbRK959ez7bEAV1Q6rbCEJXTSaktRT7R3/JdVunaqGtpe4W/Iqx8C69I
kcQuN7zFZzR1t3DUmH09qMm/YPh0B0mzQRhkYMz+v7NO6DvLkCH1tq9B/2/9MCGy
ngyQQdZV17SS3pkZL0Nm/dh5eZkbqY3Y9zjZ9N/UKNhcsX1hgrdg85SO6rhXcFWF
UimLlHyIm+fTK5Ha7raMlMJeT7aNfbfT1i6L2R3vwTNhsz06IRfiv3FKuuskebN0
oqfOyzuoHaa/1OIEQiDAylm7wxbHjRBCh4bz6kZnkjJaUUnVGgr2MivXSonNKu6+
BtEJaLLCgqbxU1bZLfizr1IkhptZbShpQK2SasjvKNXUNxza/sBLAv1+j0GwHVdu
qYJoj56zzJJafCzp3opXk4aIhPYA+wWYO2NyWnX+mb2OBLSFZccyZ4IZppZXCvhW
GxZea639KflHeGc/S4ikymwUiJO8taU/+vwsTY0+jFz/lS9Xns7wjTKNDd6RwbDc
g42QQOxfwuMFxD55KB+CnixAfMaG3mKXvt76EIQyHy2XDnfbpAdDeHfXw7EkDagl
PBmo7i6F38DBDx4y6Dqh1EVhKJTSJCNK7WopKHLQGKzn/P4CqCFlAKunEpIXTIpG
y/SvOHTFdlbZw834qlr23O+R6gxuRm6ctFpQO+Tmrfx4Wvsq3SLUFglJmA/Za8G4
kBaxixnIMlsmk21RR7JiWax8s2goPCiSHfxGTRJvw8bWW5Trg5gkKLu0SfCRBawV
o+rIfZmYHFVKDW77Yct6bNy3n8wC+gJGI7Tnkg0uubPMnPgx/BBFo/6j0RmptBS8
A8qW5Lp/OeBv393vnnlzo6QCYsrdA2/zVVjbnf/QHkSyZ0uxZR4uollPJj2CPWYp
70rXIkkWMFlwzN3vQw1WCLu6+meZepWhWRSskibqeGLn0E3YylkbqFzhi9CsB90Z
xGmHDLcGR4n53pPCkLnN3odYKggDSEaO2cXIE5S8wHA/adQRxe7uoAltY0RTQ9d+
LbVpE9nsGSBiQ3FSY7mO1oGvZ7M2IKExMb+/Epej3FZbEJkASZhG8IMHmgUNabvM
BjYy+UW6ToJMzZd9UxbwO6Ba2izRPq+zWuq4Vx0gy9a5/B3wOxKS6SMikSxExggg
2b3L50ou3dEVtRA1vvcUVAFb2bbNpRvZvSXjMJPSVlZyDnWnh9BrfFz85iUR1ZHU
8bx3Xyg566CY5ZZ1WT9O7oHXOGLa+AaR/mpDGQ3wFHBC8by6mbBW8WjPM2bmMHjO
ufPCrIoskz4TgWBmu3a7TvPi2ngQyvDrkQLOjKPNBDYyR7AZHZgp3pU8ApjoKNmb
CsNTnNJZrpsG4zPkElRZ6OQaOL5HICfR3maSB5UGSiMDcnuUbGYHNwWI+nZKu4RV
UCZeEP+p8M06Wc27sZoOr6vmMW0vj3G4y36vXTnf62h/IuW0KTWvc0t7GSCrTtYZ
bpidi6J3CppmhOYWJnv1LEOvR1RpRPeySqwR82m4LrFybI4vDJ35QZigPVIJTazO
NzpoKipudvHX83vh6WQpu97kAYm1UMhF9rCFkW84Tj9Cc19XOnw4rlclXUNDif3k
VEfGS/buDwJHcZR5xM8YWz29gGopBlDK7yDT33b79uRlbGy3njbpICq8SMAZiwYl
y0BeaR+QJjV2L1Tc7yhbaY3H4URUiFAJSed8bA0MEZ3IauMlpI6x+Iy63HAxOudU
DVREniwzbZIPn92rwDIrLkcJgDWR3IXhPUNSRK8FdaZ8zy4qCbpANG8Mh6qMyart
09ESKEzk4ctsCRstRG2nTqbU4dtBM1UzpVgv00diikLp5+WsnyJiaOwYgy0IDVRj
GYi5vsseoNXPY7UKVfiV8glQCxWrm9yR82q7srmp4O66ALLTmkaD/WQfZIWj1eo3
a7T1IkNrl/7bPtdyNcUt2gLKWIbwXA7a+LQ/hkSPWDRhdyFDVa3GnGIHW0yybjj1
nEXP4aU9SLHtOagT9HrrXX6jRfY4d1ocSUhMfXh1bUS3wcYTUbcr9uiKmUHX6/tV
d0M9MaPLbP1UjlgO4lLAVvbTlB66pddZKc+TPjMmKbdGxrnRSpggNEwku8awkUgK
0ohGxKJkchLeAFuECE9S12OmhypbDu4OITAU9tdOJUEePRz3Uhkd/w7+cV94oPPa
35rFT67AYnLLIQcnMG5dUis7BRdIQbeQzv17ALG8YbbUSingIlKl87ZGtaQ3uF/W
qWJuH8bT0fqvIdlyToVZQhJSF6cY55rkqd4iclkchMNBl6zB1UxHFjnEGAdm273g
vTJl89T+v68DoqQpbZ/xcPbvZuvmA5I/WlmBME8/hee+xqZN6+Fxin0ZfPs6gRm7
4SY5hJ1W13ROOC/kEkMB3ERIL5DZfXY8CrPzPm0ev7RuuaiULuFNp0WoYvL9+CWK
IbCRIsXJwwVrXl3+/rrzeoXgzXE8RTQO5BzfIrsCfCC8HGrw3QmtJGz+S4hIpoR4
7aiFc0ZFhWSrc8bnKTH5t2XnvkBK76B1c4yiZ8afJVhAHRZcHvn8GFdhvwEuz7kF
TXoo49emNPMVPQ4/Rs1WIj0wuTsrpTc7xeqlITJTqnWATjzFfR5FnDdQvanwxqrN
dNd7Wf0AGuA/0gccyhOuitgC46wGxQvSeo+ZvsAW9vUbi2YtzK5FKACV35LcTT9E
q0DgAOxBpu43DiLrmW1DEtQ4xGa4/IFwVZYNeWsV00vYy+lMaxBMXgGPU+zMgg34
yndEpEMaJ3HnPDl3Xz1Cpgq4+c8GMvuWh4491eaH8q1a7ITF3j+lwMJo8JW3ksN9
4E9DezfzYOiaXOx/gYrWSBYfJlnbszrHOWjoO8HC/Gje+caqSrxq3BlKyX5Itmhv
zG1b4eU0yhi1+nyYZsdOTL6E2eh4B0xBwtXuByMTZ1+4EXSTxRhDhzlB3apI46gf
N/x8IE2zCzXmxZNesAx2EDmhkAgt3bIBIeRBW7G9fAHdcmALMDedrPdddRA2Ruwg
+eePziic40dSvw1c2muV0U8FpaL7CO5HJQO2LKfG7Tix/+u5kAOmRaAko582l12t
c9ATVYWhaPoqE3WIdzGPI+n7Ux4RClaVeNKZeuIkJQwq6xB1pqprqqeETnU2lnyH
taeasmBEfkWcaKqSTPOFIOZK6s2InuFDWTJARoGFG900zq3HxEytCDI7ypAqq/1z
bDRvJ6KdsjxXvDjDYloblA+SO172BnrifXVPkfAtKykIfCUdwi9uCm6On19ly1zr
B65V/vHWSR7E+VPSDHUDsotbvRau73NYWNPffnuAjU+FtY78Bo0HVgO6i6wT4zzM
vqSb8Z7F+vT8YoDCAVS/ZCCaqlXz5vub7iXsCGttFmsqF/2PGrBo7keJmpUkB7+k
B9xnQKLEBNQquZjvNRE+xG9vk/C3o7Z6lzblYnobZJzB7hYrODxuI+E/U71jEyQm
IZZyL7Q8Z36OPVW8HAR9CqwxOgnV7KCwWBBpflxNIPst8Rg9h5onzsFQwuCIzpVK
lHZYPvvgTzYELMgmlxoc/O9be0jwHNy3ValJaZnBeeH5aDBC2w4bxhoEsTZszk2S
uF86/WKkxMuwOhkhXmuU9lGiXABV8t1NmE5VsgWG2KyjQ1AVj3IuiFa91VMKnxuq
e2zcwYMmWyCXRz450wnyYkUwkswASnXOG6RiFNg+cpzNaQhNSalOzPf4zAH+JG4s
AVKQ3RaL5Gdd0+N4Idix4YpZ/892ZNQBuXV/GuuaO63bXuxIYFAYW/ckagteOzIX
ANvW/Yv6DkwMHh1R0J25ErNuzHAVS6s8O5ugNRjYlGWeAuJfKrfp/a6q+poj3yLw
yu4vYrQFcPBXbvHTuzMRm54HK3Fp0VoTnaUMxTOyQQlZmJaA1aUD+axKmfFLC4j1
4rpc93SrPADUhbP8+P4LmLGBebtb7k5+UYEtm36n+lceyn0LBZT2KhfRTh5zFWV5
aN0CsCedto9G3ynYTDaon/8BXu2CpFjpMRU6ydNA96sU9lOlxTBXnauU11jQ6PYv
tWiLqIf+Lqv/q00vJ9bBgAcwBNrhUm9fveTB75ueUWLzfMkKW7toEo4MpcylL9fC
EaGtzodDgjsZwMm6OR48caLvNrQCe2BnDtwB2fB+PhdZBom1Sy+s73RnhoLZvgwg
BNp3yxKuhTdqmxhm80WKNLVnrZ02b4M6A0MRD5i3qV0DSks4wnTsRWyOP2V08/D/
I3LrDkgb0r+GiMghJCqJy9Fwo1pPjZiWkRxOWVF0iQOYTjOqbfv1HyrhuDcbne02
9nCwbRFTxsvrev8QhL5NJsn/gbPfbFoop/zfSj1B9tDK80zx1jZuEmwcvuTh/dfq
QdkX/tKNujnU3iSw+9WRCUht4gW1eYlBNmKebhr8I+KxwVQy61xTR+DaTRPg0TaZ
E6PJ3YhH9AHxVBeC0rX1HFUrYqbI6f4HazvcQ+LCRaF+ZKpRV62LqokJIr1hG2Eg
uGBf7Ashwx9wP840etIuNQwLa0BISPR3I147nlsL1bqQl3bZ7L1M3IhpN73y0jQh
SNJza2KoTV44+8F/L3Kxge+iJw+RHdmlDm6bPOqU03IWDvMPyUYocUQfgJfnkM6G
lnCtuAXJcZ8Tuh2/jXQdz6LPPLmsAb1EimPJEurviPfwTxJi8L1s6wxVexpVMrDR
UyLU5e3wv957HN7Exj+xK+tJLa6JWz1/7sVREzMpim4VWwmhha7otNHmpyR1NFSg
IWBxYoiosL8/C8KhFG8hNgq4ZUWtVDFLhz9Lqgrid0HkUhmB5VM6wHXGxlctnLMo
FJDKMGUzYr3ss5ItVyff4kOwSMXc/uo12vS5vUcQY1vRihTr7GbqEVdx+fbqQrMI
pv2qkkDE50nhu76l7e2lM7p/Jx0qWBEuJaTB41maQ+zD0jD1MZV0ecjYA8mYTH73
OpdDDjD8COtMmRuo+Fn3UajgSTH1XHHuJh68nIWdFqrC3vmFXGzqIoYG7KCR2i3p
pkpuDmkAvL6pEqP3VdB8b73C5QR3EHnXUWtOlV61uj0I3zYq4wtzBwSn4rO+ojWe
N/Cexud0kXBda7ew1qQALJEZVP+BEFO+4LEsYRuHcC/LVBgdhByLALTfAaZcscvi
Q13A4f4Ft8285iXbyX6UwSDJMchN0E/4DtwcFVGl5Nil6pn5HqbzYs9sDDsQwc+M
skJ2/bgaefsrOAsFRLdAYPSO8tfWHKfcVKIWBnsthuWm3CNG/cLUCAMOtJ+S4GUh
jVnEVOBNraXuj8q36bS+zQGOAdxebNzZSDyg5I5WbGVKCg7SaTCZ2hof1YXzm2mL
TpFP86DJ3tbVy0AH87DogOzsuVcHyEk7yOtLMNz2sxpHl0iUPmXhMtokZOrFl/9/
b9tT3EBa2QGX5mxz6WwCcSz1zl9v2x1qqec5vdio5P3vXjabvMtQqv1cVn47s4a7
+JBArQQXHlJNBBSxbTLPh3EdQrVG3LblY6oVSBlQhv13LDqSwkN54IlkyeaLwoWM
qc+LI4lq6XK0bPstMemuUkJNExPtoN44dFliBNmUgCXPQITDv4/gdT+7bzktQOlY
CTaccXDqiPmaUgHNhgJRg1H7N8+H1eeLFBGY0+/BSZGkD4W1vxQypG15PH9f28E9
EnWcy799FbmBFNrBaPtDXzzPwd3psRKNBcxWUYF3hiPGs+qOYmgzoUJq0w8w7+jY
YYw0voC3k8vRsUL1rqSvkxK8l11ICU3gebkVFpAxy/4R6AWu967wdcdS1OvGadbP
lywPf3e4ziedZCKOcAJCMrBgQ9so/CeLpRXLsWUS1eSP9PalnxztoQAIzn+QsqSX
gSwT9rv/00T/LWEOLDNVbq+v1GukpYtSR4yBresSEzfyG/RJMpll5Jd+kTciRwJr
mWMdkqCbN+11eUBC3EbjgzgOfgESCO83qgYa/TNg+brY0vhu9OtmwFjO1MCLaj+z
j7uWpDtuQUrGj76lXmSWziwdNHBFqdt+qomeJ2EexB1EhViF6KR4X9ptOI9q0mRa
OfrhlGnRQz7StogfZD16QKhk2318z9QWAnprc7vsQJZdnfCid/BIzdbSZLn2tKpb
fr5Bh+VB7ONg3C6jjn8RStHTvpbTWcZMRPXoM6qAStiK7YZpolMHSwAN7horhThe
gZCoIqkFGLFGdTVatbw/HirXh7zXsZCnOR2V7AS2J6rzPuS7Wx5Iwly3jJsNmj+i
mZPjucd96oAepbLt9IelFe6SBSBMLQ+EjIyaGYYtAaVNLqYOSwa9355nFzEj7oUB
eVUgCpADgiQ7OwSxh9vbOVJBDfztNsf5ccPG6sD5/jRGCmjEsvHNfOmgRb1dtqkE
5JuUqCCbaGUd11ucbncpgp1O16IiJy4qEzbwWM5EEwXK6y1llE/ggRAXJILnsLHK
/dEmCiWZSzRl4clOVTCMPgENspfP7AOkFd6j7RqifKujHgSrNTd/iaCRFKopOfFQ
J9flmkPVD/9VxmyN8hJdkR9ofwDHsdARoFkUIygIL6tbzZONJaFC0IViSf1xmX4R
6H9HI8IPh+IUTU6ooXsOjPvb2FMmlDJ45iqkceDhn73w9Nq2kagCNNa1uqjGLXY6
MIpgh6Z8csMPCe44bjDCmNn6ahCTsD1mjomrvvXqJSDGlL1ToB0yW3NddGuXo8Gz
d28/Do3oLpFGmP7d9Gfa2jpM34rBZfXQjKqAcCKAOeldHNB3g2amn5y2hiKU9LXb
GxzVwdQdWf0koPb5UGVGLJY/z96uVNl+z5i9AlZ1xOoxHmnpnNGu3sqrNdwU2NUr
Af9EJxv4ZW/O/TvIcKcMuexotq2Z9qzdQPDv47F+uGppCDoh992YnwRAu6P1Z6Hh
lEsddAPt4Eg2w/166GeVypJ2dXcex1/DDn5KhcIVWxqCAQ5DWud4Zb1hmKy+eS8O
ept3Z5kPCUB/OjcFk6jzSPgWtVLmk3/uPAuknqHqg2UbBmZQT/M38LhE+9gF9km5
q1ZNoBNV3QYh/b/FlzHNvrSq/iaS0mFI63i7frSlTg36FwfkJE6mUBF2Fz+N2lJQ
Cn6+kiO6t9u6FrcqjjVfqQy+hoPtmRThKTV4BEFxFG4vc74ODDB4mhOm6DM9i2np
Qsgr6wf75VjFpRYdlhiGNaSt4nc+HKKWUs4j2sRg+GgJIGNdt4MG9MoGj8fgT3sO
c9a+HtAP5XwoFxUYxBcRNKsFpR3M3EBR3Xrte/lRHTo3a3KwgLVIQ7f5CA6u2thM
ZllF5ZxhHhU4x+vBsOh5lCYiOEtCXNwPscEJVDYkemv8IaF0myaZ50l8g1qwah6U
+j3tVMNc/cuARpk3rVvxgMbwlIsRtVOzFQpy01rvOv0ZSn9j0WUpCvurrjkDnIIK
3QMCittqgzbl5TT/95Axh/JNoQoW8OzsKnyAZGtJ9HlGHE+Jsyyjk5nzyWHW+g+D
QmEAE+s5TsW3CfyB1hbotktxvNDBrKGk3dYcXyTVhj+BwqjFLWEF1cOzPw1NlYyt
cTUHf0WIZoxBq+x4CU/ifzYZFg8fWtTuvnE5brkUVkdtAjzShJB76dJXhR65P2c9
kvtKTq/2hpKowYzCJvDmt+WblFfMeTxUyo1PaBOSnWWE2AsKUCCT1oNCUeQGwdwB
G8RZGYP/Y34Md1OUc211bEl3BjF9TFuaPCf6seFQTqAJ27zpfCjfCLkN0aaiTBww
F38+HblGcApdwGLlH4krhPihUxldFk/cRpHYLnEvPbT0J+R9QIBYynJVH2PiOznS
DsZzVQfBYexHoyHI9HbjEbQtDf8nm+YgS/70kIuBfAJiNEd+AO+XAVBeT8QLvD+4
GhEiN0dKhSngCK7xrUnvH7frm4WKn4zjgiOIQs6UKv8wtuJH2rKux2T0KM8TAeWk
hd3VzcRYiGOlQBoBPCq//8WyqM6Hb7m74sn8q6DSQ06/oiZTfO5w4EZWkaXiauVU
nPMxoIhF2AsKSFe/Rs5O6eoXwn0v92Q2eEi90gVhY0aLzJ+ABYvq4OmbHpNaE+ln
jv3tp5sqpb+mOlqxZx9pIF6pQJaF+Xs9+uryC6bW0YdrRPpiZvhNR3hoozofpm6V
+vr/2x0ywfW+OfQlGmFhQby4rQoKhj3l10M4eBkWsq/PQoOIYGzkfQEFBYUXcU+R
K3IsCNR3AnOWuqKw7wkf5KPCXczKiIXPK4mibi0827uzf8jkKsXNPElK7XUcOpF9
C7SEFQars/EPuxN/PcBDRV8Qau1zMd4hTEYhn4ktBomRiM39ahOrF4gz8E5X7ceg
eeEAZsFgWo5ZaI23Zjka76XU8qCngjdUTnE4UdEsJC86qm4S2BiJ8qDRPI+mimbJ
DPkalr604p4Tq1sZyNkh1hNjjrCdSRPj/RDKaiODLmFNk6zK53ugzdB3dX4cnc2z
RLzvOWgU7/mzpKLNMIxhRVduwOmup+UR0XtcJGzTgEFSlamO0HpKrPprr+AsUNeT
utOUDT6nOGq9IG8YCHaKcvuYdAV8cyvtiDd7UFPnCtqawlBUofur4A0u4ClteJ95
EZOqeHIDzGgJJQsBS3P7oxe+pxMOJk3L0T8EdbfQm+d/2GCQCajqwb87L0KGjjBY
gcXUDiCmviCOzXLrFwJfL1eXXESz1YsMJIhzwealWOyd3SUb3iMkyoWXWbjRKF7S
DXytd7e3lLhHlGgbx3I33hAI3+JnoaKhzX6Km8JHWd38NBlrv3hKr7HlMql79Uak
nFLU/nO7WAJFTsq59BIbbY7FWQBGvallsl8V9pjQ6wWuYGBDA6tsZ4MqRy5CtU9b
PmupQLbKDSseU+6KaheYV8fs6KCM7ZF1vcakOxW/rYxxZF9acX+TPg4iRQM1digc
9hEgU86aKKplzpDYXra5SwLh8gvGsSWqKSie8w+gM/tkurIYWS05DE8ts1hTmtcY
YGyZYdzfVU1S5+20cFdaG2yDIap7i+I7z4kQeljIk0Qgm+lWjqzcnZANH+NRUoNf
ou09dPYMO+Ecd4lOdSSXNrwI3bVrH71ZkRyXAOCzt4qiMbRYoGsUjwVIUOK34jbV
FSvE1BdmoXbROvDhBwXzeA/X6limTDGXCBcu3NrZy4eaeRTmU5OGw0tqkS6hE9rl
dEVE4j1Ad3N+7yj1DorDwynmLsXyNQtpI9NZb2bV100Lvh52Tcc8MxwpPD4c1qSW
VBo2kJKgwWEeuAGKiKjVvJFi018jjl80Gf/l68cxzQ90oqNNkqnu6SyEucc30UzD
Rpc9+46YXzK7RRtdbybbg9eLoYe3jLIyfz+aJLxxZFPCqqhAGA2XKMCX+GUku3eM
ET5vdKDsrI352k2ElJBx+lr78lpVQOzGowTasFJ0QuU/foIgyXFvHrmEE+QLyt/Q
SDuI0TdtRxSBfNlp/iZ4kH9x91m4YK+MiTcIaeWsPivpNTFZh3+uO3tEqTDX+39S
+KLdoz5Doda0FztiK4wdTpxJgtpLevoKkz4nysGfOGwJ9vYOo8gN+tUJJ+BAmX/W
44egN1EfZ2YxTrGdbWfbzJX6Lv3Sf7YOk4KBEZul8qqTW1K5+EdF8GKlGSOOCg/8
JILBz8AHZ93Vp5c1sL3wVhzUpf/EVsI3o9t5yeUDzLeE769UHouJWbMbKY/g/XQW
BYaU0QRQ2Q3yskorzPc0Vb+NoQ0T7JAD1eRZDBM1sqM7QPYDAMjNV3Ou57dEpx8r
gaMkcCp7UZsSDu/GVKDAp1X7tpyx5qhEPXywgWQHtbaCwUv2Jb0TRTzVjnw4qADC
PRIptTc5WnhP0YzFwNwJ2Uc6gaTXzwkuR56h6Qjolc38jS0kIUilIstdbqhd1kby
YtRekCicEPrwo5ixSe4dUfYsDCIA48UWkRDYXYk2uDo4qLp+DUsr1V2Wcd842W0L
t1kkuEMaWxHTgu9qEZDP6krQLID1h3tltcilOLgHtiF08eO8hwqkbE0tQFvyb92c
i/Y6y/lh2ks9W7YyrmWdDgtgCMYJAcgMCL5oVllMqOxkRypHQI8LhRehk0pvgbXa
P3YbWSOg7SJ3R8QCsQyNySSUCWRcw1wL4eVIlticy1iQFy+DWaiQ1VSCiEAcrhu8
6paXWX88r4OPowc1WcAS7aZc6kF+BLQBc2qg7ObIw80PQT5V6n6kqRxCBBLvgugC
//5hxuM0BFWZEXjbDyZ3VRjreRvgOPYWXIYcDymvjrYA1LMGXJr07kzxy5MRG1Wn
Eqw8lJQCPXIzDIl/oVOlUKhWd7HMF0HY0tQbz4DBR3dE8Kvtq7vfysdoNK8yJdpz
WbaRIsei9JN+m0uf+lQYsNOKGLwNQLUVqgHvvSM4rzLtPDjQddtLsasjR7z57A83
aQJngb53ZYArT9nP35a1mLQFRYlVx30mstR22JZXlfjyef5W6WSqk2ppusibhBFt
BNSuQ8UwW/I3D02UX2K90iCl/3jvXpYlOKETfBrJ0lsZqginOFe9CGiU4jS32yt+
bJBKtpWKwAG9bFidCdPd7tIzewR2Hzeo7Nm4M0n7F617OJdwaSEstcQQ8U1muECi
dzP+HY0EUomVj09DcLYIDdBbPV3IzaROGUAnPDyopueGVOtPJ2y0T7yYfgO+bDJa
gjtK07AFvj4rjbQntuF/5UKWKBhsoTUqlhfoYSb/sbMa3AKL6c3npcAWlFE6b1Fp
Zen6uDsOl+iLUlfh6Rk5MtuDqsdhdWpdh5wunyGMLBWmNTzty2R9KDqf+uGhZp7D
4Pmx4dkULbvjAHVD+0E+J47UJlIJA3aAVmCUTcZ8l81DUOm/kvGEqj1ItsTa8ijn
rqrdD9cg4mUZaY4Yav3etRPVFlj3vruLjoTlgw2PV9+ijOaXxr5pxX2dDPhOBu7P
sXuQiCLORFhjOAdAOeAe+7FxtASvBXIVn0LWepXBz5oGuFUKd2tpglC120EhnSRF
7b8nXN+QbWFCYibFXBxwJVKCQodzjzlIQu00JPu0IvWCbW29KhrvOvlN6bD5MGm4
1m3GTQ7qUuSc71JCg1IY2gW9IG2FJfNAlvIjv4x5PBXo5Fwimv41vpds17J6ezr8
k543iHu4a1FNcqB2gaGnvFdwVvG+Mg8+5PROtycloGD8H99xf17B+PbwkoEMwL8p
+U2GYiC48ZJcWlgm8bQPVwfytXe+oxNzKjRINApLKTVFw5PdqKq06LMZjfQqckpm
fh2+DYTONK5Rd69DvC0d3UXKIjMVvfl7JLozp2twigonJ6QGHEk5LAWag8Bg51Q7
7yrPw/FyRg5NnSiNjakIaztrQtHq/gIVP+k3cj4c5M8k4TsDVtpkdZOTpJ9vNQxf
6dSp5BhUbTwYpAYsS7TsWBZj6GbGw0eB+fYpgEzHMZkBcSsu1Uu63Fo72ufACQlv
NvB7iSLm596f96YdWmyW8KF9Hc8iEMd3KPwWk2g8KdpEzKPbbjshQ7qWr0Obhb4o
7PwC0CnGd170biisbn0LsRAXOJCrRH1P7xerh6ndo7w8pFOkmqthgPxyY6J5ZIWE
6RHeMsEHybXWBhFrI31jjhhqHVaFN8sVXYP/vfl40otWpl2PskyswqDpnesW1J6u
Aw3AvqaTzqJ1owIM4Q3JPxE+seQbvqzVN2CHcysQ0BCpsTZs6joif1iGphoP0jaf
knos1SNGpZXPE4BNonYRDsMiVni90ezIgrvuAXgwJPxhz4CXNhNdC+6Q6irWs913
/W1oFyCUXvxe59CjTFWsnEwidjrJudkqpj6hTLx2j4aH6fLTYdlkHdwd8rBGVMRx
ZkuU2Ja6/ceov4hv/t7YLPJHU46kUZQvRnzSS4/ApxmOT3lGCSavbTKw2KqkvEW4
iZH1fIjrOMNRRK7ATci10TqDZdF5zPRE2/+bzdcV2h1Exty84ryeyU1Q2M/PPsnY
xO4QbF6L9dXxUQkyVS0lKIc8SmKJKj1aS2h6PbRkYna8LaB5D16PYr4QDgZfMDgz
luRmRmfnOH+zgAduzi2ocnb1ZE7+968JrsQugq42Bhgcz/OdgtftOOM/T37o3b+p
scbLz/tqy2WV2xorWBmU9IhG6OpjxtlvUBRJDVYk6FDAHhLZtuLGkgYtlVeEpK9W
U7e9uzb6yo1KPfHO1TgfJTOTdKrWwRZoKWul1mXAFBMcL+7S88dYfzcjcMrTwxXU
xl95OA3zBbDvub7JweLAS028aBrv+42ONCAmF6imvx3WPBS98oUoNPkRaMtw5Q7f
ZvL1WJd8xvmic/GWgZgalNdnpCs6jA8YvFsw5mouYFGnOgcS2L8FqlTmFL68GP7C
02UBPG8aWRocj0UPeVLE4dMpX9RjsGwI49uLArzTFRJ3+Ni7+6ynFmbdHxp36Ukq
E3n3KlYzY7mRpxxLX2zmNzDoDMzGZCButWbWSvbmGpFJqe9zq3GRKCf+hbKItZUQ
TtiTmY0m02B355hb8XoLVPAqnPGSmWmhkYPNHf/3AcEmM1l7J/61iuaPONevYSEn
GPY6W3V+qP3Up0MI5ipFa7GGEQ0SyYSqAXg16hGntNtaofj130O+VsIxhSMl/38A
XdzPkdu4cg340CwLX3+PW/pEOZ72M3TZ26oLIQgEz2tJYaDLUi+Bdc9nH06UZke9
ODJjbYo+gADXjW+vDjzhspNbKENA1WhQg4h/6V9eZcF13CtT1xV579puxQL6n1L9
qNwhL2exFUazybaeH5C42+ZsExn/bXWrPu7YV+O1JPeg6OZfHV7hM8gabfgHQK3M
1X8OH9Gkslosj3ISLwmaK/EZpfII67pva1iwfws2KU8+aCx9URAtCgxyiABkAkVR
dMmM72oqKVYHBGcDPPzl08jrPr9jBkUo6UZp+AICfv2UzqYbO7deCF3NyWMXY6F1
Ksyg2BqR1YicevIPuoHfF82OaCXtfYAsGgAsYS52RiRNQlpgMVN79iuuDsmbZ1pe
RQYXEpfk0znUsWpbPr4muN/lw8khFAUFR/i9Xj5Gk2GivZl4E0D8vA3IymD9Lk9C
FM5dtTa9CF2x+VEiW8JBf87QryHf8S1M6GhmJWcX5pW9RLzVRHIVbAy+NTtcdUJj
EdxIlx9lVIvWs1BmFAtyEZqSSvNEROfZL1QDZxTtoyQ1SfKuuMSQNUvP9rm0NFuI
BAWlgIZ1dQqeQ4+w+seBJ6u+0QSIygKNfZaO+2W3rYeNmHaDg+wPN9CDiTol7hb/
4AXq+NGv3GMwAHskIwPbVvn4Z0dirNEs6GMoS7xEs0CSZn3QXKCYth2GrFzksfn7
04uBGdJoV88Go1nusVNJn1fX3OZJsmxeVtK23IDdOrkLC7qeDHDn9I1bvGbBKrIL
st17IjVc9Iy+kcNvR/7mC5z4NhmXyyOcbcE+5SwZKo9HCfaSwnkWsJpYdMRTmTwy
HOTn5BiXqOBBwJmYAG5eO4Bi/m2sogHN2fEprioXn2BgAHM5kTmcyK8OMUZhhuEJ
TxJVnNDq4YLir4UQslRMtwYN1I389Ic6S13UJ6Gdc30JlhoNwqfyaYIUxSpgO2Ha
2MgPtZ68WTCcDqmsc0bcmhBIjeQFmD9llBN1hI8z3lnijmUNYlvoaKHKaPKXF6KN
8GocoKbsXbgl3XhFUaHTdAjIUTmODaao8zS+nx4Ni1oRX505ohzgUmLSNnJwoGBN
4aWvKpkjSXWwWFX/bW/GTpX9NXszQ9dlwC4A2hxZ2LDSaVmYBqtyIGhtPX401VYp
JiOFOaiWar4i/CywIRDr/0w/y3nvd93aRAOe5PHWA23npx+5RTzfppJcmzpKBZh8
P/Z2D8aC20suOmpO8oCBMUMlAy6UXETKqKwQBVHMX4abG2GHjcRUbjHlnvx5c5yO
tO1X3x1iTkZBZwnuYiEyCFPlHLCOquYqziOaQR/8y3DA5qJM6tAzU11LAuZq53oe
H0r7xKAzhMa0ORQIlyn3KTTZfD7prO0a++HNt9XoXyOTf0wjq8dKEw3lMsrquQ7X
N8tBFdiFk/0MU1rTXRJ7vEm117qLKmHz9QuswNVjhVJkSvpEcBFf5M5gPKaxaytc
ssHGNJQXthDEXc3a1k3ogRlBxuSjsXHssIeDMT57FX59JvWZXbPFx5Sn7vY4qSTj
XJ3yzSFAQLWYQl1E3pJMEv9DVfP9sxGPE2leJx4MhVBCHmFMPf+HurDGDaLTzNRI
KJs60/tVk0euT5uccYU5a1Lh1f+NnGPOigP1u+j9j2cgMEffvka6C0Jl+nbgPGZv
Jb1hznmMzNXecTbJ9WSjLwZ2ZKtvu7K4wMru2LdPgb2pKJEsgk+hIu4+Kz3yLV1j
RWyPrRDGA2HHVb+YjTPjg4N2p3Jx/NqFFKAlSVS2ksaWBNzMq84QjFuQ4iGmN8kY
FGgutQRyx7zbPgfBoWqNclOHOdqa6q0xoW3OA9s+EmCWIckie0aZFB+ntiSSAmVL
hQbBjFcziulmz3q//I3mRaCxiF1e+UBcQk/wRpPGLhJo8HqwyaonMVNM09J9yFbi
F1VuIBa5cKSon+GcoLFO3znODegZUFVuzUgIiMmoft/ol4fBwCuCJ8/8Is42TQ4a
adSV5QBkEcAiIhJaFdq20F24hQwUGoaRftIyRxY/ijTk4nDe12avqu8xwUJgF0Wa
xlb81FvECyqlOajwl5ltSrhazmu5D+9YeP4VeZUagnrM/0h6Pf8QZ/Sp1zsKdEZk
YfSw1aKQNmSLt1QktU/w+ol2zbpLjbcx/WFtIo8tuDXg6F4cQhsNDEQyQnGuzr/B
K7y6EawGCogAQ8h59TiTrRkPy0B9XxdxkRGz4XtQgprehQPZwa4p0A0mzQESOKeT
+xSSKLWgTKfFUJakxSz9w85AUdFICxEafo8R3TCrk830tNQW/g6rNC50afGZ825K
S6VgF7QgcaZ4gbHeK+RBjOH0B5DNAXjvGRbi+CducTo6qWOdkGkSw0UdL3MAL+kw
FYHOwIH/sAswursgsKlLmaAkk32SnU3QF8fvOezq3MUTWhBc4B+vrH7E0gSWgUk8
7qQQPUy6YoNQMTRSoCDfTG5OHuRfnBsLjLoen7KeJRLck2lKFbrwtZS22Lb2RBpm
QxM9LEJpKC+XMS4Cpvb7ANQB23ryCn6xn2SeFOYXnZA2x7qbfltHhAOleptz+0c4
Q/6Q1ucrqMMmSdG2ysmiOdVMcNoE4GV+gw2aSuxj8BTzETniBR0xcaH7r55nvKb9
xenL6bn9/Ud8GrHiTHLy/QQ6AzeXJkulpBA1ru7EzV2tCGFISGPoEsoficW/yLf9
jaU7MUGHgsT2Sth0urbed03WOxYPJAd7mQqxBhR/ISDetRc/+lBXgAHyebbkEElC
px4AR5ZYXLIndEJwkMJW3PiLPzqxWxuxavVtDCpjXUk9TR4aDSR5LaEXxbcx/vkR
9ZJI/yQe3rPD5txEwz3OMVteXYvhhupaAci3zNIeXdVpoZhOVNMDacEfH1PIk62v
MxsMcF/x1mA+OicbLtWa0si++XNgWAJ0ITKRJqqsfmOOaxIdZ7On6BP4r0SPfW5K
EmV0wEaFUsZRgUC9kBRCvzQz+k/8UFrx6DDH/88quWrTjVwPHx6risJATd0MP2sw
96XWk2VHsT8IOAi0IcYlj1yZyPmikLPH8nZ6tfQoNzaTpX/r+y2TbGTXqrmpr0tr
rkiZ4aTkAQDZuTE+7Xius5/0S6n6EWTT0Kdd+W1KgjJtITnPUClKeGci4Yico/xy
ZGSHbqmIcjhTBqcBaMFiuVTYmw1nwFz5sv7Rv6c/dM3WfZ0wayq5L4pcBY6KcW1Z
3OOqDLTNx2jOnMtP1QTHEYyD2esBUZ7kk1MY4g33gXK/9iGp+D91zOmenXMOQkkT
841nA4tT7RtNMayc3rOlw10BNJrOrJ1NIyd6r74wTIl3Lvq6fJPsrdNf780ftNh3
nUhLmvWdSCuwrgAgGdVgKG9YrSeBePPOMihA/azudA5EQ31abE/4c6Or2oh5UMfT
CQy2QI6N5ATfoufVCVDHCAu3mo5C0GYlxWDpiqWXHTeWsezeIWkuSYmP8BM4j6LM
GCE902kDI2Ysc8ixDAy/lkkwne86LPPBXVLu+E0jVmhgKN34F6lf3/y0DCdVaQI+
nFyebCmeQ/+p0w9NRx0GY5IspxfPZgeYwgBRFqp+scP+VIDvh6Ki/xXneFGFL5AW
HcVTZb5xQ1r3AODYU1jaGKQGFSOGb761iQDbe7znkYNr+3OM7taP0mphmpoBw28a
6SQzI3rvD6IKjP5g6/ZQ+cCEI0F49YirbM8qMtAcCyKp15DKzBWPU0OwBC4d/qvt
jGq8iy763F0+LfZEj/KHPbt7mZADn7rSw5YKZkyX/YynH9efRcltWPOId3Pvb90w
Xk9PTQEDlsCxTgcWQvsP+DeDnlvm37gcSDhg/zukkqxdeY2hmNlCEo+OoH4fl0O+
TMwV6B6UbS3hyZ/D/gtIfToifVqmGSG3PypkPelo9osnB9KtBYgqO9sj/yOX5wnn
KWhD4Qyi8sgrwtVCyxDuuSl6WL8UZv8PjSsAnx4vG3nh/2IgNAs5ryGCVSjs3rlu
APMBcKhh7ulsfYUAL4+XCqS7w6EhCGLnMLQs7w1YDwiKQtK+ge9II6UZiDwutXFU
APGaCwIfcrpX1XRdsvw6NjvGs1/AMqdgfHswbsx/KkbMYv4vRChgRtM4sSvteAoJ
`pragma protect end_protected
