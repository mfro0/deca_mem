// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Swo7qF3bd2n15kJv+pKi3ms+QuxcZXcq6OTuHZZ/Qh40BeZ7UO/g54XkwGYHtR0C
v8534FTutjNaWO7fsv4wFAfMLJakDdpusG+vOiaHnVG0jRCXrXtDBGtLe1vEg7Gl
mIovNAwwxb/UHke5wSi2w/KqoriZOr92EiX3ItsNjvH9RqImnFUAUA==
//pragma protect end_key_block
//pragma protect digest_block
DkcG2l5WLSo5tCeTLl/yfXtRr2s=
//pragma protect end_digest_block
//pragma protect data_block
RgFFIcEzlYOx8d0QOVvRB0ToVRyt1H1qcEdhX2/mwBRQlqZvsH4ZIN2EPinKWjFt
3iMfSeHK+Ai+VFDraIVYH90FsPG/orcO8DYVcKVgHUi1gdFFrmoPW1d0WGD1NfPT
6PW1i6iejFRM7iYTfNj4g1V59heDXx5udJ+LJQ/7qngdJvnVEFYk/UHcI0P7hYEg
5gFAQBXaErrhYmagtKiMly+7VVMdt26AS7u+6+rHEs5/K27ObXIJvCu2ZjQYkiib
qSiYBrjWnrncrWW9B1KGGsaYcIkuY1tnMW3PIrp1PYGlih7sVLGnVdxqrRT+XMoQ
KpKCsm0PbzRhb13i9cMAhm8QUK3XP2CTLWbledw0Jfx8BZHpDxqrfqWKS5i5B0lt
ImX9ApoMUtjKf2nnwp+I5EAhdcU2P0FYYRHsAmpMvI4q6RA5AAOt2tdsuuy1j5hz
PUA1croN6rI0epVyLzW93sv8ZqhxWBT3zdQ9/jUJzYNhMClg730qqwOlkIT7fepG
QHc/msmTz/AQOk1ZXtFvL2j0oz4GLapgdEHNnFewxEdIFdyzyi4ZtaOhNR6PsshX
ER5zatc7Om+1sXxtXiHUKTLEGuMuf1isK+xZ8kn9EOKiSaBeZez8bfP33yqmWwvh
yulL26cYpnMTQfRIR82svqIBgvU+LyyxYs3iVSbWoDnRpDEXitU21jdX8XeyWPVY
0hqglcQD8032U0HQVgRJOvKBFmyek1+oaxAXMXt9UN8tXMIfJKlYBRxQcUKIwsTn
uYlpX1yDw2izAt78/o4Wtpvj5UQ8YRo1TRdbVTR/Mp8K4YhdFZqM+/fKLgAE/JSm
eljxpK9iBh4hTwy7kH0b8sQ2QpqZuarcaWDpgk9WNJwg9QjDCx/SUwhAS6JyxHmL
1v6c/YDAi4hOzZVhDpSQr8wlSvUAb4/BU77ccb5FqYoHol3YoDFsEqPaAX/TNt38
m4KjMTVQEKlbm21Ac8O+jgSjtpVvkx/a9Lv3mKXdpT7LXAbQxLdsJj0tzXsPSaYI
ygk+ZFA3BKNacLp09HhwB/XLf6DUI3n5g5fAgP09dNq8Tsfh0chTO4r3BhSwtaYx
biZtsPZoQrkcmY8ERmi9JkmlkzkabD3FGze/NFWsYCcF+nocSuJChYCjPblMjUmR
uTlKuhlcPC+Z9TgNug98VHDs2Niune09362suhP+dSSKg18bsW2Vl08XJTQSrZEm
brwDraVHC8shSzETsYeQry81RnjV++uE7wyUCuMFQG3e+WdIY2swjY+XPRCYiuNO
Ev5ATRdv7AYoNV8yNl59PCZCtjP3j05N0jmisWXW+zZtPZEcAqik3xiAX/WDUTQi
YIRmufI3Z/sr57lvT2SusvQppaYzU04oBuLPcd0njvsErQIXEVLXR/N+gK6bim0E
qvpnZwlRVCs+V+c239rawe7u/DAZ21L6nJnDMgtx5nPKr3gasDGvj83RllJCdwRE
q0818CZmH/J1XJfDvba84FrxHh470nPm2JPvWynH1r94rusYAXzSXYjzi3h9p2Uz
0UXICYjQkrk1SzPsY6jY+tVGbdnNOiYOYEPxeXZ4E10bBXn9b71UXirXcEIx0VEG
prQEreM42cP0pdt2R8mD/e3iBd4TraAiFi2HPW1pTopbCwKBzzKTH9Les6lxGKyj
qBnEEfvxl5ZFSiO1+nTHmWDGq8KJAVwjzteiBPYYMqRS4NmAQpqHAvKTQ9MGaNQn
MvVLQfihwcNnIzvNEk+PEN7Ukz6JM5W26qecZJtkeXgLxk/Zv4HpvAzQBBuLYc7B
v7JlByo1023Yy8Tbjzj7LniBmAfDqQJbY1GU4btf3LD2Vt39ftLEA76AuzLhDQGa
LtBW8O171yO1PZ2Vbd5MLHAQ6abkrN5l9Faaw6AXBf+cBPGzMiRbcC/LEsftWrmS
ASO9B8NiN96HFReoF5Ah+3i0HbkWKMuryJ2EHho58iKsouGXJNTqZKoYu0HA6DFd
6glhaDF0wOhgCPNxm1oQrma4zGdlLUUEBV5wBjka4SEBxU3Eq1YtcdynN5CObSmT
loBgjqpXprL2DjTOfu4RDVLvRZ4PiRlqh3WSa9Q75eO0rFz0dRPJhtbLnxzEGfpV
/hsF4nDuRnEnxpfVxpaWW2Hb36SPySOxJ6GNwgA0D6YDWyBy4EtdNFiQbtMMa8/r
2fITTzQqMG+Nm7ToPdUCXuV48IWQoIihxXQfqEYmGobJVjfqg7loZfb1ZbsNuhUc
g5z8kscU4vT0YU3vfv39N29qkFL2ncoMAr7I+CpxoAc4qxIIAVfIXr2G/+ePeyds
0ySGHC1f1inz88xpBMVNYGYj+J230xBSudKppHGFqP6+yLkZc/dizMd2rpStIBW1
vuAxGLMI5jsXCf8UGhXOq3OKiaYYu15tKaDqc02AOfAThw5VmRF8V+Ay+0k8NHKx
9apPEHXP1VUzmULufltKNlJgVdasOC/MBMoGgBFGZ6X1Gqcqb1Hetlw7YLjCFjh1
66Ox54LZynk0c0blku03nOEMpBTPhLoTeahgu9HtncscUYaKrnltl6TffQwI9tjp
LawwSmG7UaDbRoCyGuuxc4wTDgNoXz+7Au1qCG2Yb9UlAOBqq7b4Afl8VygMszrs
XAHKiXeH1SQXhL87z/NqYeSVQJse0EFGUGr4V6WCn/b/Vj4EyXedpulT12tYJI4g
tvIfZQjmjqTY6ZdLZSlGReb5QNR4zgWgsJjdVKOkuzkcSbzolccAbSOHUr03MxB/
1D5O0DOWqCh+kQ0HRQT71zH0hm4PI56e2+JWUcws6cTLJ2jSiDSV5FTcXQOP+xkd
parV+5js5d7UYM+STirEUnjLzvE4rIUjdT9GqwflhvJBzO9FRk72MF6lWU678YgY
9F7zwVwbyOI2PmkidXAqaw+9p9hevqIS83ZBKlb1tTOygkl9AqKskvSMRTMTaMdP
R5ZDJvWWf/Xx/1f3ur3cfHR3z4ivb2176hTU5uEwpzPPZ/rpG8WAKNjVWUg8aE2W
rT4ulYUz0e5vCz6Uzm6k2AEQ7LYo70Xh0s+S2jwBE5/rpu82/Hzi2G5pbyT2q+nT
hS6Y+7IAt9Ouw8RH9r7D5Sa0WlUbfq8b//8ajNKE22HdgZFzECzpvuelglM7ewq6
hV4CKQ3mE1Q/6MYQ36D+cp+W8rTm/TxxLY46NAp8Q3kkjFj3tZV/61/M9Tl3lMmm
tBX0hG5ZJSbrLfh3zDmRnGZAFBO1eKPzB7cg8M5e1IHqzTT0xJ5osq0iZK6lWrLj
R+vCftbzgMwRnMeDj6Kzf31m/mYkr0uDKjmbTqwgrdtN81Ct6OMe39qRAqyQ+8ka
xpzYut7B0r/cjiRnsWJp1Y5z++O1Q02lT6DarifPKJlZIZBbaXcyIMThXKzPt+k1
DfMVHdeXTr8OHAFOQJ00l8W+jDzj2CiEM83CkngSSKbkthL0BOutClZfSrZpXUSg
aRo2ucMd6gEm8T1C0R9eH6gyl1nd32tS6ImLMKZNqYWzOBZhsnOoEroMzxI7qkRU
4va9hPEGeWIxyG16nM7ra5gg+WEr4Z4jtBhQwLvQ7srIAO9X3mjA5uoke1JzcjOD
gK0yJhDJcQXt1qJ6TqPKLh1MeopoVcSt5hZCG3WenazdikrCsZtqdRHew0OKWDLL
GZ7A93ALynS1ViMcAa+OE4hVGG5WL00E6vEbsao84f3qlfwdwzM9CzRN9sIOA/0n
uPMHlHleTFXCyBgu2vNcSn2e+FoLHnHywM1Ys07QUzVoYS6WsdZiyyQkstoYIHuX
+7oVtyQSB1oaYbeE9HTQntmiV3OHvsCOIQgd9fcoVecnkcnsWLzcEAHboYma/V3s
X6TKeqvzlx3z1vKlMjI8oUOBFYnqoF5rauLruIRiH7uc/IpP4+4d68pYtOeSB3lm
ReFr4RT6O761331uI6buORjp/L1nUwKQNBX1hA3fD1fm97DkbpF2MhOfc4BxW67Q
GPmahirenebpXM9NLND205RTefAMhWwYVmofy6ikK+LtFlSYNtx1tmQSgONGXl1x
qk6aqszo/EUeBwkiLNJ6VngAXHGIRv20sRNMbf7mmUDZbR2agmLXdHad0mLAoJcI
EqKTx739uIxH2Qjcnu/XoVt3Vt/ecgFaEyWynQnIHm84x/lPqP6UP9vVWMdTShEi
ud1LA572wZmR29igNOQfyRkHtuj95jUXJeJWbBUGhsyFUcuXuL04h83rP8PDEA0F
VBJvaEKT0HDpJw6R43TdRQ1pLOrlC9C9oB9fL6p2Jx3zmRfivB6hsFafi2nPGz9l
xm+CKqDjJYQhanP8p7mleZx3jUYfrvmCjER9pGRytZIP/2jUnFP7H51U/mMk7vJT
24SAwSg4FnXnQoIsThicqHevI91nHO0UD6a1qngL+h6M++xNS4d1feik8bYO6LzY
b6Iki9WfhAoX67HXTfL4SAlfcolPXpVsNA6SL/oA8IRc8JKe0dc7puaAvlk3a5hU
Q8LxyC9FiWvJbL8I++rqYMu9zUxOOwqfTENbyw9PVgdRNHBlGyfzt9D4KLD7+aRC
oDiZsf9XhqK1PLZkaj64bbISTpflqgd5xbj7KmABmZ47pP+Pb6sgujWyxlsUDGnv
kM92fYJqBCyZ0XQP5SORBHpGS7N0HPwrkhZmWqaRv6jL9235IBWG4GSntVONxSMx
Qxdfdl65Kd3AUoryrVWvA7o/8uxMnWqkBNzV5JXJd+rI0JlSkMa17/GFNZscREfJ
4r7tPiRVoMgzuDEaAKNLm9f902Vym5+FT/iCTzm19/T8aGbBhd2Ob37LBt1OKCzy
VDoqJ6z6K/6TL73Jn6BgGqMhNjsujMvDv+E/VH37AHbgcifnLCR7e/mb6Vxu/r6q
QYhPOqxeX92Ml5HX13t2j7wvYkD3kAX0oVvCxaxoxcD6t4s1wwelNNstQlsW/zDH
Es8yHeNiJDVsQiay6SYbWcZshZkbirlgQmZ2Pkgt1vUH7th5RzSCOLXymi+zaeJb
ayp9e9O/bQSMOhxSmIzApB9B9Op5s+j1+RJpMO13DgjrkfZz54HJVwy32Z6eRlnT
tDpmwn6ygTQ/J1Upp9cfJ5yf1jxYiWh+ifuewUNC2ilT2QzxsRNvmioQc7BxAqfZ
r2qvISD1dDVr4Gw+yF8jTbYBy16MCRFwTArsZcXvfvMer5gLciZv7NJ88SJIZQH6
PgfNDiDQP4vEHwBgMYDedQYvQzgMeUFppEB+a5wXyJgHagfDWfuP9vRmjV3Y4oaN
pDeMxh1Jba6IOdeNrPuwtfyQAMlsrK1pswNDo39Kuv0FpZm3T42kSxNQc2YFyi3z
D7ZJbnwx4BTyhmwsPj2xxCdozZ6pYeLTYijVwoLE2w0Zc0nPYLxWuJ4fIsq6dMUP
y+PIvMK3RGYD/F7MxcghEkjyP/4NSat+w4/F2NsHxn7FvRy/Pf58L1K1TYsUnarV
9gxNMZkzblRiyl/BtiicYCjttySXXQJ1LFxmEkehdEUwtvDCE6fQNgBb7CP/G7HH
x5sSQJ6kWVoNCRW/ZGPOt8cSwNVhfS5kpx2tLGrU2ZhWuz3pkefZqIO/mIy6uE3s
ht8dI+BxP41nlQD1Y3uRTFNXYBOjmF9qMK89REx4imwkUFIvt5gWI9lIGSuKaxV5
ZdCZjO/QHfU8JGq4M5yALFzCOmpuw9aGN4sK9GONYwy0aHBVRlG0TKSkBPYqvjW/
bWzlnTaoOu8cPmHdq/Omaqfvey44GK65A1hlV5mNOa5bYXFNAa2ddN1DcEw7wda8
zGyrH2+qdW2JkDDpNgXMQ87I9FaRolToa4ECEzkK44RRyUGsQgt5ReT4/aY1A3IB
yWT7yxF/iw90G+zvC4NLPWIxb3rvM7dwovuMw897P0vcF38tVdhyrukUb7KNUe3b
ERVGM9T8KyHP37C+qK0S+XQmg+qNk++VNjp8jUAFZ3RNHBeRf0nPajC8BOVZNYFv
fLNuYLBHcKIlZQllE4i3gwUOvV2OOHX0IN/MQVmXZ9cS/aSdzJAu0+koIKC6KdE+
UPx/tKVeKCqc6LplHmA2OWWCLSgDyIl6W7qBsFD4UMnsifMAjH92InIVnmXx3djL
/GuRfhRYfUNLyOruSp5Ua6+3Iw+0h6sMj1fY+vx1+GtXMWgfmyi/F/Z4y0l7ijcM
0viey+9NDytAkwcOnujTl/YEKujCR8IBtPG6QoVaHDuuZ28C4ntutDqvzxXgY+dR
gC3lwd+xiZNwTnYIku7HAE6tCTJvQYcjsYhyn0Qzm9Ah7822pOa/CrPvWixsElwg
REv3dRBy/xEd9LN8rm+4r7/p68L2HMTLuLZz8CAzaOb7JXQlTEV/PzXJ2lEWHvMy
Wozr7JgIbqYx9Wcl7PkDy14a/Ws60k/+SUblQ8JmdIFO+GzPv1FgDXZ8+Njeylxp
1oaMmd18+nlLsjotqKLtCuKPzmJdfJpz2yL+ATFMO4hB0dTlsUqVqQ9zOiV1xX0y
bQXWEBdaEs+8Da30c5wTkNRrT5etXj6AbIPqKL5xst05+ZBrqQWfm9xMVZGRmqIX
PTmgbxU6EkM41MNOnKtIrRxJJybMIJ9NB0IIorJU9eL4adTR91z1Aqt0I3txLrlQ
EyqP0EPor9QRabdtnVpwh3xLXwLTpSopOBvRP7Tm95HmyuDPDD3SIQi31gxFpIsU
LgNslrinUOHW4ScD+AVkOJpiXsvDrftOcS4Yl1oDfqwAuEPMSxoSiPx17N0H0O2h
kDHRre6LhQKypI7O4huTDITgLuPfZAyOfZlqdJFMdSH/Ub91dkwlceYcRfjTYHMs
PmhYeqX0dYsq7NVJTxb9EkquZoQ0OXsXee1Wz1YkTdJGzS1MWbvowpZeluK9/3IZ
yA3/sTX6egiNU1o0txoyi9Ir8bnb+/v3abHSxoqLZiUm4FGsG6wUgEHysAWRo2Pl
ow+4Rwx8ujJZ90GY39yqwieS5EqFzdRD7D+XTb34UV1V55gdRdbYSK1Me2ktJtmQ
8cIhWjqb5nE6ZaGZeS+UP5144i/hAG4O7JMGGxMjoToKcVzkppDSPFgNOAhVC+ka
7ZuDTg2kD06TrhuJZVKL28ux7bL9JkzzdJLWzOXsGVEqYaYOhqb9bnOpDbm3wKq0
eT3YQoNJvdJv80ZjXbqHFTOZRttcEUmZfun0ydeCXvSz264Wa2UFgvlwLesstufm
kNJmj1ZQLCuECE21ijD9HbTa+HLvgWyVYEusNYcelajkcH8aA/7YM2CvhHue+O4G
RkYtokK9vMB8cXHraTEaBuB+YY5bW/bH0abRX2Y8aU33/55Hy/MRPiz1Ie9eqNI/
Y+3qN/rTWob2sxkZDGbPiD9ZivLbyYpSRW+Jcmv3xYzE27g4L25qR7XfYAdENKPC
YyclUaJtz4GYjgRfP6a5Ru7Vfzu69Py5ppxBU9e9HEcSxQXBsgj0MpzEltGI1RTa
2u2Uoyu9QU/DoMkDjOO/0LkQyaQn0JdtVj6ystOhXpxMWRkT2cpaUNs2n4NryEAF
cWEg8VUrzbNX6cdXdJi1HCG5+iJeV1McJxnZWulqtU6hI3BfCx2N84XQmaqAlsE5
lhJw4Ue12Y4GZ9ZknzShAiUaeVKDrbiCNkkbnjzSWYtmoO6KMdRVFQrvUDpEO+9m
otD2+9lSXVZiLwec9bPYCPZZcPt3Wyw5aH+0ApS+MPtZ7eqSE2BM0OgSidbsTFMl
igiOXeR8g/m1V73QyqbM2DLP3rLL2sef9ViPzJnD24lmtJ9YuvTUeCHTwWQIQR8N
jmAOoJlO1PQ9YMtXGDMaL6BBkjTjYN4zn6t3mvSmhflDGfa00k/HCUUqauf71Hi7
68RoAVpv5jEfNtl25HeEUi10PtSGXCNB2yNqDdUt4gV+H3UO6FyYGsKH3sxG7AnQ
yQjEJ2npYH5dRXy1k1kiVHsHvNi+Vnf8FOw+ftl2oHA7eWmE7rGJwR5CS1t/s0gj
tUByDbeuthniFeCg3NYL934K1R+Vc1I1FDlYzhAmgg+JrVdxNUbnkuoF+abOZOu/
UyGpLYBm1+V6UoL5HAskEjjLxxcZkd9R9Vytc46wgwHAupmy+42kun1g7c9YW8Sz
h+obDHiwLyE502UeiLyOLl43FfYIuAiRy45NTF6abUJdGhal2pY04JGixS1PEKjL
NRI4lbCT24Md+cgB4nIGjA3JagC+mnBLufB6fvouM9DzdBA+oCzyr3pVeVroUMKz
59G0NdOOe3D83js1EyRXrWqP+nN8f877F3yOQQGUQO1YfoA2zgXr5096Dp1ov9g6
zcvZaYkPZ7z5PaDYM5VVFL1XGob12VIoCIUouTt9p68AsWZIfMdrUl8hbFVJxgYc
aUBpKQFQJuzO0jiZjYYAY03HUd6d+bIIrkzy27KrBbsnxWJ8dOhjEe8aYeC7Zvwo
NvbHM0aB3V09Fw8sk6zNwuMK9vzB/F104vJpWVFoYeD8O6xKrgcd+CYU6PRlEALN
JKd2S1AayuJMJqe/FVpvcLDSbo0c7elqr3rs3dEggWtiVBaiRW+/DEPuRDVzWq6b
JXR61mODlpcmFgfRUwFzvs+fhu5ePufk/Q9xd5dOXvrZ7R34fuXZKdF70MrtJqtR
nSoKdUq0EOXP2HeTvsl4c1Onl8cwIXRZAegV9fAfyWjq3ab635COAjJMbbqGwSfF
lOb2vRI8K76aPn4XTDifDwbGLwjy8Uxs3sJ9pzvfJ3Xyq4LDSEcbOQ0NFg5glhdh
cezn9OB2eLLHlAWFdmoqNlFILr9Dn8I7dbMhpqeVvdpH13tFKrom1YWnMVyc0bhJ
0gg+DTgJ60P5vF8S88R+FHZT+nvpUK14FyTwCeT+cuacEv/y76vTBrFkK1UzqCBA
IZ4zhZyjEzuaUs5hI8yX79F37WVXRVcSuGFKapglBSFtZkH3uZYo/kMo+IdTnJ0S
ck7mK17Hq5UsyxFW18i1/dzur1c+CN0yPrELdHwaGOBuNkX1mQyhsgASLYyUQzmV
LQb8l8V0XYUq3m+t++l8cK6+3u6S35idWhGsKgIp2dP+tWt7ybuvWWETav17XjHK
U8mtRv+gOWAiETC3lJ9zBdUK7NlTZbjteSGj39nBJ06XAU6BXY8gR7J8AKAVXkcB
sQyFRFdy8fSALQKNTGrvx2xyhvwJFzWpo1sMpvzDGkW74R5zEgMaSeXLT4Gc4FM0
wGCY3SzYYuf54TZQ+ZVnQJiAxwR4tidkrxBclCQGq7a2p6gbPTkn6pnmGRZklW96
micdGiUYVj2a7Jd6dDIC1vVvsNGi5iQOlJ1DvfadQQrJkAs55roBvXoEiIWlPHjI
IIUGZsX2+AhhXxshrwFiuEL5pRVzdpI+aIkO5OZOd2cGgKJIgvUJ99Hl69gF+2Ol
vcyrRhNxNRVqqdNVdCgLNOzinsHNp9VZ19Fk4DdgveR3JH47c7+PHAuwwjH6M7Bw
70+BOSzaJXu7Zib19r+Hb2RybBXmFBxBrPSxo7UunGr/r44zo4/91G/kk/OmfcLI
2CprePL4u6tfz67ynjVvGFLtHKQZPP0P8eyY0S3CH5f78ZhVHfT+tc6iggMMjx14
m/y9UHuwo7jCR0dCbutD4jZVNopd/u141nAzSDZ9pjKM6YequoRmE/Vm2aStGzRP
woKjUVVDw0cIcOIt++qNkeG3wlHc6p338wr8vzoXRVxPBBtmbigxABd6Osga4ll/
0dK12aYMH4DuTG1CCL5+D5EVx8bTJH8WtpAJGw9EhCbuKeQspeTySN52pp7C+6nr
b+zWh+nORHR9pmPfva89R7RNYadJTU0n/Vem7HcZPqxUecQ/wMeDpyEa42lKPruo
UyBXwEtkiTLHbmZp1UqXz7D59peOAJXGPIULm+JGhS4h1dTTNHoXbruup3wRYHNE
tpzJFSpbzr5NJdLh+//qDdJPbb3IaMY6J7mE672iJlOCOQ0+x4ASDmb5H49KMEty
qtpf6OhiRjtpPUWbt9hkMVzpj6x4m62oaoQHHRcr4/YmJI1U66vOBmjxVHf7+i60
zGqj1Gw9y3b6F0sp8blL/fBzdr6je6gncHFEC3ZpLFirVwdOY+EoGaxuZ6s/YHdI
aN9HzwRGbCSzIc2cgFQ6P0DxLPxUB1LRzKB+jR58XKnp9u8p/d8drko10EK760qP
RIDhJtW4nI2GpnX26MnNx9oMVCdWQJxysAGgs8oIOu0c2ZdFzk2ZsLGguVHc6Qqs
4ViqYgAL9uy2m5RoT/7W8zCwWrCU+WuR2+2JRqmqRe6NBHGixCDJw6POCZJu1k3V
LQNKmLeUQctxfF3MkeZ66ayiLoe7BJ1HBuBPA7tUpSKrTbzFobH03Ek6tig/ir9+
h740aA3cf38wzh1+V2Q3na1Ry/EnXL0y9VXKtFYYT/wGDnvXWiXzpVO0dDq64mTS
sCUHNjHA5OrvGjK9lDbB3Kh2wTlG2Wgr3BWRBvkNbeqEjsIFHSniUxPuPIVB3w3I
913kmlNoT0V9loprMUvymADS2Iv8iykpnrA8QleGPuSQDpElRsGtDdFbFvoJSTho
l+S6jS6gtihYRUoScqR4vRlWblMNtfs6RBIKGx2HO4m8W6rT6/U7N7BOVGZiuU2L
mgAEv3OiiyROkfW7otXfajYWA4mYNqiNI93jcUapANu69ZomGr91U6Bjmk/0MLRl
SA0x9iylZ828qJuh66YddZXWYHG2i2E55oznn552dvblLY/Izm4jcwCJSD9/kwJj
jljXklLdJSJxWDHC2gEPMhtc+PncwrxAMblldyQBLkKZvC2PrKYtnc1b7XSnIEvj
joMxcTXYw/Woz+aV3jUB6whYOn7T3/Q36imzQRpdX2CLExWUqIntlrw5drMg4CrY
Ao6A70W+L9sYvFlxmWoLJrM8aSgJ+EJnxgfaabTqNgH1nP5CkvQz5Uhf93TttDQg
vO3MEpXXHBFC2TfoWpT1TfD54cD0z/+8PG5oMkiu5kFnMpMOJw369xV89x32cKjB
v9py6f6BHqu1Zph5YSIV+hGbeC7IsG1RhxIzcJXgfjI1se2ROxzXgfSN9fHvcINf
CG2Mv5vW5F5ILD/ufxGRZmgSHFUaI/JMQRBEdDXuoxEm9NiSXjnUALsAQnxaXKbT
ODGq0osE4zfsYH+wTXe7YqystiR3kHNiLLehQiFF7bO6SKYfaY0aFtfOV20H8heL
xD2dwsZaO8lzihkxTfcnZ1mgZnoANt+oczMmktgIK17/uwmoXVts6u59YbzoNv7m
5lcoy4bbBDExdI2YoxJH7i8q5pSgs9PWvim0DmUrvHQ6G/GgFkeDFy7VkbWQKSXl
HOZ/fAek7ReA4XUSWhxbxN5YazDMhHSwRyEFRvgE9sXHxog7d5y77GqkYC2SfLK7
uWizyLajSN3NfGeH7lSmz0vW8EG0Uz8pbuwkcJKHjpEvrKqnxhTMFI/+CIKZcw19
lD46pD+DJ+ncNPY0mJJn9VPgSzKGf3yL/+qCwIQ2P6H+g4MwqSiwrtidlDNeQxAx
OVnkJC0mzEioGjzq8J434HxYMykCm/naqaMyBVfKXpcG8G4wZmTvFpDlYoQJjRB0
OoxP1y+pw8YI3EN033PH/irSrhpvCnc7FDDhNRm0T88tT7twhBIsRa6OIOINY0wH
CiiAmrr13shB4Rsq/kPweYeuHiU8vTphCVtTlVLLn4ta/n0V+kHmhwqlWBgEY/f8
Bs0tBy92TTKK2t/iMX6CYf4bJzo2027JkytCOVv/OjFTFnjPCgI+4lFYmPTjjfmI
UWqeX1nPHUZDaFd5UjO62TP6OjlmUPGnpnXuw/Xijd+pOUh2EB+HS4VP5noE09aK
ovjkpD/+IfQNmQHNI4AhXZIiFip2qOStV8V3vqeV+k0JSsCyQtKWsOaKTDsOBh/n
pAoOzXscuR97FVgbWYPAnCb/ReGssE8R+7YphKPJ+ukjwbQMHuCIJtnCdgLQu80E
LS23g2RfMl9GXMLgJasLYMIYmjPxiQp8comKNvb6Ao8a+YyeYXSX89Y11XkcW+98
NiFaBPqB0naqctn9lwdblMSyHmzNPIXOZw3vNuvurG2bEcEDA1DH/ID/lW3kKiWl
788zRQc6M6gKSNBmzKaj+00jLbcYVPOYk4mIDEOSvNsXFM8A7VWWDF5iXUdCgdcy
VtxhTPhUS0MzNbFLnZv3AZ767xaVV9cakr0FaYPcPIisAb37x7odHgm5lSOPZyX+
A+ErSj0t65rqQqDlgGZ/6r8rUZuvmzoCIc7XyOEWsjGfc8HviHYT3xgxV4Y+RWF0
fMP6levHWfBeA9Ccve/fE56tfNoZN1R5dMaSCpAgbGgqAjIqCOaLnUGPj8uqAnOi
9vBfN/qagPwnA+D6hIMExeV6BMt5ZSvly1WE0sISJGf3zOUmouo1q/JdN1KHHK8m
Z0wOTLuRNwHLCBU/q+SSvNU2TzWue8BppP6oCD7f7bWwK5omVhaKncYpqtK4qofL
2GS5GRa7QlGBTtSH5z1EEZoeije6+O/LdLY1NNbJYD8l2c3XeQ19JAro3u/LBYiF
uceg3opwRoXaNJ2Hium+iquF5kmpb8wYUzlBzslhUC9pSapzk7YI82Zta5W0UtoL
q5DsH0zOlv+zkv1R2fEwlpXAuXvuhMl8H5ikI6+FacrPq5BFMQFnkZ/ro3Biugil
PgwTbz8GNRs3qE8Z3jjW1B9tsxwVFVvVua33ABwYKful9Nxh+8kpwfnQY05mvUXG
2WW1h0VbpoYPdRo2nKBOy+0aZJrapSDQlXX+FkJoy7BB3DLgrufTUGnv6yoJAtd9
8fmDMttaptoPydRrzPc/jRix2mcTiRLxE2EwpPVoSLs2JWrjL3N6tZpLz27gQT9a
ee5yHSw2nvu/Ax9eoaSgIEvmgyHmlk0DYF0QrYhOc3J/SdJ0q+BrnTIeOioFWh67
/H82tc/z7zsz2wiBHggO51yqSRWe3m6qbVEjgzjehh6dIlN4KZOdl9tnuvoqlDud
86cQRUND908TFTpWfyrVSDbf89/OkFMA94hz1gf65HWnUy68PiCOS/8xTpuISJK2
nNgaZlsYn6s3x0QL3MOGUQBf871EeeCa7fDwDQx+Wu5SwNa/BgZ+6+8cvPQVIMUv
wsosY/0JcowT7m+vkU6WVvTnjojh59sPq0n2z+OUMQo5KKm5dxoxXg9k2t097bWo
BfIBXv3eu4wNC2FRqlyqLlT+p3hbDgejPE9oWKOcquEU5eStGxtCjHxWk+VzrtqQ
5b6hA6k+rdlVkOD6Tgd8VU9NPjZ8Ps1Dzcp1H4O+56EtK91+kgDqvFlzatkDrs6K
koc6LSlWkUWZxFFhP29SQA1TIiDN7pwAh6UR77BR14uqgKmFH7cE1HsXJEpxbRKa
EMHW1OzVm8fXlmeP1lDuK5Kx560sD/qy/8mlaXXGxEhpX6NNrqs3b9Pg5Vr2Z1Rq
N6byXjyDMBHzxQwFHA867BJ5GT0Lx6dG8NsLgm9aQloOWEouRZXzD0mGfYxReIGG
xjD0w7Ix2OHg3KE5Y28XbfA/aI9dyBqDGrhGscrH5/JzPjer3MkyiVI7y2udrKCv
dvCksZadW3mAC8QHkQ1IjSIzDDoh2WJqDp5yQSH6lMCdiDapXlgu6egVbVyxT+RH
g/hluAb6vc50hg3MLWIOYh7RJmPsWG22B5MjSHkmpvX2oqp9xDpYmImYJmFeCtDZ
16R+uBCf9ITxHnzPFXlSJOJcDwbxjTMPqFU4wsx3d5Ue7OnugbyDOoVHEmJCpbjQ
wvXtfr/SLWwjAjpbJYlHs8HAp1qCqeaUhxACJlhqBipoicE2UNJWTVBB3dcOWz5a
PjHe1FRqIfNmA6IxiHUQby7MJwaOCa07/uuJzYS48EZeo1g8cXlN9qraFVWjlYK3
W11i+v9Mei1Jv8r+T5Ng7iJc6cmq6pTGRNcTkzwRJa6WrjQbUmX1uMOv13kUXj4o
HpYGVF1QlLj4nvtVsu364kOWkc86PduwsDmOK1EhIVEKGjWD7Dvxr8x9T+8d5T1G
HiEcSlDhEmyD92LmzXdyGzwqgeESpqesHcJ+Ir3VkxXehbqNzWrJA6Q0ssZWClnx
L3XmkhMFiw7TamAkCcBcvzAX4exCqJfqEMK424IslHuBDo+dtDyUeJ6PB7NSZo0k
M27lTCXKJGYyCDdQaR4Av1iqhi2c5QBAWMk3vVaTBCgEmWJrDwT+C1Mr19KTysRd
Y8m5/DsUqpE0YHjMhCA+jSrZQL/8vGruRQRva09Bg1utfgDy5tju4ITlbz6Lsj9k
85y/Dp4oGjCSqWHQ57/SiiXJaUeJnCIjNuVQsureUFiZzGqYkvSdLr455B3bc1P7
Kz7zDAD0hMxhdlRa70l3hc2XwpXb5RiutZnKRHzLN/HrGkzrzqg3skLAQjLZLYFm
glbBMPRmZXJsFXP4leiDJTAts840SGJN6t44SQKR+K/w5nRqkXZfDjtmRPNtgUgD
7duCgrLxo4DdRKG1iBAqLB62h2k/cegpPYlNDz0tCd9ZKWZKazVX0blT2SlbhEI0
HF2PVr+P3i6AOzwKJ6teFMX3ik9SfrzODj0hLWvcbcvvTymlC2VnO1w0Fy8hmDy+
sH3TBoT4yPJodli4NUMws8vuszb8xYCdXpXtrMoz7Ttm3BbH2DSdH/tSzCOZ0187
XMV5aSP5qyhOPozpKZWMla+eF0uCFc+PNn66kFB8h1PbhJRqHh0+oykOdYEyV2Jl
uDVK7jKi85k8rARndXezZL2ygXzbpryn5jTbkHj45tSKnTihomF8Jcg1CNidcJ3H
KFG9FsXe8J21ScXzV/8RsEJqk2wEOj/JiJXH9Uth2wfoJvSq2UxNWT6EGpdUG3W2
de2foVal0WwSzi6KudqPfxM6v0Fh+OToIfNq2iZaOVsryDMsZRe3x+5AszkuT9NW
dlPnmGXcRXWTTFq+19sfGzKuLQDz/LwwcPj4lMzN2s0/5iHyer7eWT6m0Xe7c8mB
lo0T8PWffBdqscAM9o938vqvVLRdVKS2hXwlViiKXR+AEsNEKRgaRNiSW9JFTnLY
fgBwx+r+v9X+wWmq1pZZnaOfed2oTeH7hCIQMBVn56+IB9NWZLYdYg5txXrkTdmq
hBQ67IGQYceE6LTgmpDHRbS40pP7CCa6wrFYG+98dbvsMOmZ6mcvwDpxHzzdDGUe
c8rEGx/ZkS9cnE0Fy6j04SGduYLMEs/1QxNKq+51evkK5fzd0eYmlqVap9LCk4cx
dhPu8JKMu30Uhs3s12Z6fLvGBYvAp+ZYcqqq6gBgKVpY1muwI/R6ZralMV5O9zs5
CWEVAeG5HgRG7SNHXuJXegcmMC3O4iWLC4qTzJ3VZ3LsJ4ss8rhsxYQm6SWEKwhk
8gl4JJ9eN1BSQBq9lUNvduAo3lcilRzJKNEfwJvgOfITzHAXJpAsrF35J4MfZ2wC
LAxwWfVk2dyxjUcFOIieBqExSXqCiEHVV8fwxiIYTGUlP09vPBOzUMFSU+wDPDnt
8608voj4sRbEz1t35TTk4BFAtqFEnPMoflZO22PzbPA2u0eBOXBGPKzWEUtNnP/s
62UaTvgX3w8oqHuse8W/iV9B3mTgFQj1D18JuD7RjrOruChPs92sP7GZcyuhxGq+
UwQn+T8bVDr1Xk1LT25M0ZtoQZkywcH+LPRJMiOt2MRcnaQGV/j8Vlidr4BpnxkK
1FnaEkXrl3y1gnW9IPrVv3nl1RMNFO09oj5L4HeeU8FKFfkr6a54xmADq/B8QhZL
aYRUrRFC9X6EqSR7t/4XR1ZNCYuyjP/LDIPZfn9Jn8psepIXDIZmVI/+Mbl/gmIm
4hERhYJ5mQVf/3HVYAJgV2iGBISoc6rddrnUx1pM9eiHwLQk8yCL8T8uz69EmKY9
3ulLy5QvC8dPUmXze1pptyHV5SmUpdxFGVG7u3518Mr9EtkKh3z5cNvs9TBb5196
oExEVDdy/qJdN19SuNbuAvl45wuaOyVYOiZZRbdQaqQtXqQ5FbuVNZoHH8J+/SE1
UU7ebYjDjgIuyRvdX9bzq6HHgnE32/5pgCRjS6fkcmWPSmFN8ewUi/Fm95o+uanM
LVg+2tj8XLiAv2l9bJkopNJDStHCn/s9ip+5zeWUtgCkMfv2eJisIA/94Ah5D1RG
j8lFyrtu4YBba0iGWmf4CmVRNZ1t6I+GbQmF41qfZ+ZnxhPtn428f3GhfWR/TcKD
A54zRFVZcPIHUnQG+6IGyag2o6llGJqNmQfmSNh4q3k/nyslZPkwlH7GGKe+Ly9W
zDyN5tqm51CcpqSChS5Uq/dMUaBGoVsV5IhJnsIqN4/YZZwPVnOC3/Ccf+aVsUY9
vhJGS7ikToyR6HoMHD7uaq4H/Xy9US+Wo3uo50XwuVR3aAVKbWw4r34PC7eyArGt
uy419N09g2sIeIGe+SzCa+rHyvxrcUBNoYro0pNzZERLF7ns+W6eY3VZsIcKoZ3n
ID19HE3nhgUitl8FxqySj7YkMP5fcNhqXJwEKQA3hxp9eYFdcyuHhUPtebVRqDYF
af4SCECXqsA8WsbnFrUq9ltugpB8uWAO1n7kDFK50jqWoodDxcCcShfvudRtWxTp
oilfShTGtq9WSqgIjZx11JrVF4hdMgApEVPgDkA8iwtdxqcgrsLO/LGtBMo/wHLd
Y+7RXNxBMxQu+9X/69vNmtTvAmxSMoODixou626D3n3k5TpRrbWXkt+iBDg3jyJo
KCD7gwNXer9p7NljbW6kiOoGxWHFzonE6InxJDwSlPm4w4dxCwX/uXqOVWGLXlaZ
0gPSfUY8cuBCxS6y21sgW5WIk3QQ2Fzq1JJLH/ZhLL7KNYKWnOJsmiLVUCrbbq+c
yYfsWoZPEDi1xWgNdVhFK0BfkiHQ7wVnjOBrI/E7WNjmITsmyKUQViEDRJyz8aNE
yr+D/PRRuhu4rRrui4hyPn6MRuiGUO8Fg4d1IIkgCnHc7rHOzE0CqNbmyJIooM1p
Up5hn/48GsG5Bc0dQq/ZXLjh41MrEfcnREAo9sdtvlxUw4rsF6tQlhwkLW6Nze6a
Wx7oMf4h2PwtlPbTutZxHuVi+03kXsZ/Sh1SJay65Ro6yLk+BcumWbYrsQKqZHaA
JUgshWaGbenmApTIFOqrdCK01BoOOFySgqhGIv9ifYnwmSQVApPa2siCUrBWOSkJ
yyS9mRJ1qMo1w5IKNDv35YTuagILKP5oN134C0D5ko5/s6Rtdna5aIbVAEOi2gMQ
ZSE1dQNSXXFAvJip2L9I9lLWf0KJMG1FOa8+JfpWxbpSLBT1sfs7C99MoxelsBT+
e0c4nusZsSbUbq9Hah6zL8AIjl45y3o0I2LAPttTKzur6+K90NATslNFMnWpNrzM
3UrrDu5ouRG+5LALudKCkd8EJtEVwUS6K816IHWKrE0bKWm91vZm0WVS08tcyIAl
XhzuKNO8X2Sa3YHigaenvUk045+30uK6tVv5JoVxkMCMyHjiNH3rWGi5iWblEtiO
097JoDSPRyg77/8dficD190sUu4ObnmvoNviXHkx/ce9JPL1CMhmhc0wVevOHyuG
SwPq+9rwskx20LwQ0iO9RMx8DwQ23ZAfq9DmkHM5jA1cuOcyzPsACF1sz0LPG0g7
BZhw0RLNjw3+ZfEr82BuQUdklr/w1ADklr4WGESQ4Dw12tF2vRsnznojyBGybGMd
bZZWmwmRYlPyaITSheCv9W8hRcX2/wYf6Iah3Sr4Sz6LdXZif0hV5UPaN+6J9Ytd
zLd8EFR2BUt8FVZ2UFaLDgVRJP2ZWUjKp9/h0JOLjVhQWRnWhBVrYbrJSfjs7/Lv
6VcYgE0spB+4A0hYheFgGLkCGiQaJWIXnu9b39p0QXCLYnNPlJQq6B/EnWXXa6c/
qIh7DMQVdY6Py3cb3TAl8EMVZkZ9bWdT8d2fWQGEaxEcottVJ64xezScpx7nU4Ra
YqDKgZMjiNsZRA8hyU7gQPJq5hTA5sbLzDVrh18OeSCXRrzc51GFP+dG0TQuzGi3
J7jzQxhrJBaYdnFRWliHPlfVW5nCBMhiS7slL524e4xJdKHz/xq9dCgICUk9WNvO
BPtfa6Yuns3YMraGQCM5+CrquDL6Yg45RRNRQPXV7Eh68nYg5GyoqcM0sDOy6rWv
Wb6Kp49TgrmASQGVvLDtML4VFq4IZnKOOJ5V9+/cYy0tVp1/ft4r6MQW8HXdzUbB
r9TG4zi9X6RxFkusKC4FOmuSgxqmLREgqAF7+TdXBSd48/a2ZwWAbtyN3LIy0D6T
KqsovJ3czXEI94tvXyKZkBtWqJjMVD8n4NKThVavm6I7kN6C0vmHJd+GCbWJ5YZs

//pragma protect end_data_block
//pragma protect digest_block
IkMVbNFXnszwSa9acUdBKW2dGPI=
//pragma protect end_digest_block
//pragma protect end_protected
