// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CHd6iiEZYFrmXa1Qd0anGh0hWJJLImrHfyyEOAKJzrdYPUCyExM3OZB5mLTEEUnB
sjtobqfNMMQHCFwDZMkzWkmk+wTmYbPG5KX89Vii8ga3NT5nF58CadZDMpRTcfgy
pr3TrxWDYGANH1s9lKWvtoowrj8kAX9zW50ZYB0hsWXtV3PHTdnfOg==
//pragma protect end_key_block
//pragma protect digest_block
hIe1HfCxTrC8TS0P/dSEpwZ3VmU=
//pragma protect end_digest_block
//pragma protect data_block
XCnwdZdjyulBv3NTWl7ALcxz3WEBifL3si5YTdtitHLqjMIY6cEysQGoaSKvt42S
0HN0V17SW9/12CADjGf79IvbO+xAwba+JmsCVWvgCBjoM7xKLXaA4DZhxgOGBNvf
g/LsbcG0cDi6ZsOhR4vLCsGkp8Lf33kheuFhnhuDNlMSnL33NX8ub+Nxvsx9gqIa
9vPS4AZZQRbn49mjQzfTscajg9gAKUJ3GlxhnWOQl6BKrBK5TgnEWtmQhzR+TxR1
pNTNwPG2SPLgpNs0MkbsAj90HSgGbyclyPAbjyEemJAQCzf2Z2tMOdHS2NC3k5es
MAtcc4dHmnNFc3LCMKfMb+My6haBK1SEpwTR1hITdeusqQdxIjwVa6WUwPs94PJ9
E2pZDlvNY7o3PVkNb36yV9/5FLHgjZqV1+Q2AK6FZco/+stnG8z+vIeez9OnP32i
69HdxdYPwXJRoT6qfx81v4FdZOQUvSRjOoXB46IZEgEWq3nqfp6IQSFlbDHma+E/
fWoGr7sChDV+zM8olMJv5tO/XO4MeHxqCYZcymOfDeSX0R/D/60bqZKxYBZ4mPVB
kNO1AU3nLJs1gITmPxOimjhn6naIy/0XfGQwmTTMIe/sxWMh0xcIGk3Rc3X8jZoj
IVPNhlZYh4SvXf9BWH85NWjkd+WX6jumJZWvlNkm0qMlRGswMyvORv5SkV1cyT64
uknlrqzk5H9HMWvjXjcOD4ImNFHLEA/v88UavdY5/MXn4FN1cRmoLQMEQjfgN9SP
sR+ZT2HoNKX5UgvOjqZSydI/UwCtcQSZrC0GQK5h6rtB8pf+0LiChsYubOnruAaO
KAb2sHQM2EUQDs/uwum9NfekdKFTID0ZzWJtcSaDf1B/V2o2xzjmIlKtGFzwnKOM
2hbC4QZ+MbWF1D9GoSZssX+KDPNpIAfsQRMFyuVr52aYXD5/86b1v716ujgzZtrT
CLCTrn6tEYj4QK76l7rnLFooSA1+B29F+RTnLrdglhY7epfagc83IU/1I3S3Nyk9
jRCYWXKJqXRnfcAbyKUl6vaOKwHtcuZ0+zEhqZTpnAobqRkwt/eQ8UH61yVCVKGX
PkGufd4/oEeJ+xcDL0IEPogahPbytBn9VrPUIowUkJrSvLY1K7H7lP9uhT/IIGf6
nqv43lcJr7fcCPoks/RZ3KaGIi3APrYiFDPlfTGxGK6GhoaXetOx5bcxiTA40KHh
RrvAFWytVKQ/bKKRNF+nnfIzVq8uFjKBqKdUCL1PIvGwbOeYTgI8NpqTYP4YFnuf
jC2QOaVhj37hH0WEaESZrDABDAvUxDlA4K9r6oOaAk9WZMr/jZ2UHscIE8LndIaJ
YHZ5FOXqWnj7u2QsweQEXcOPuzjy33ywXHA+AdXZWI+qqhBJsI5tm+XQolkMLA1n
SAqRyHIxaPO0hnjZHuzrTvgbMBtQiyP6J0h1J0YVMteHCLhEhmoFvWDOZL/fxONE
t+XrCT0CnObugEp6LEpC8f5t+c1WTUGS1pCPunuZt/lI75leYATXI6omczIOvpIk
bz9k1n4TGa+xX3shzqzFbxNgUH520JnCi7RePN/KzkkIZyhBxtJbFyKbvykxTWNh
A8GZjUMNBisUFIA+7gVgBEo4x7l5HKDujPcwe5xxe6PcvjPh20fthTp34RhwnI7H
E4hyTXdgsdP/Js8MkIyUzDLGDyjb5WxCetpcrfgdBdvLNbDAjkCyPa0uRvoLsDBR
71EJq1Zmam1spj2qexM/m0jUbK1wLHGixiOQ++qMaYw2FkfVnc9dqpyi+KOU7B5N
phTIlSILKzjVpj0T8vr1XdPIlEfSdNh7WSIMYmHpiPn/5R4YZ5I+xlbGzsT4AwR5
VqFgBGj3o9fb4hxVXu3s9vYmvv5K+5wnFbAdUh/x12urD0NqEw1cw37YTsJ77s7Z
ZeyG6E1nRulFkGRa21HJLlLK+TFk8iQ2aNTKFehz/YeKIkfXvd56DgIke2VfR7UR
27pnmjhRRQtHmtmHD5+VoSCKHjmM4AqahQD25VGMgaCogAnCJ6PEpBHPAvLvLI5S
aU3WI10So6sxiv8Ih7j7vNetLk1cpOfLWA3KZDIAPJ97F1jgnAu/pWOsIBHuSPwg
DjiAbWre6vP7NI+82O0rntQ28Zw2TW9mfyyTtkSrSw/Q5Eaw8zkWCEdrR/zY9yjV
Agu/QPRQPBM/TdVf3l3jntlutm9VPJ2m/NVoD0gB0ufuK5cJgwISfl5ud8MNPIzH
rLRZ2Po3qeIuMenBWTgDm6QBp2l5T2kiQjVXRrSAG41QrcYyiYQzKtpSW7sS81Nh
vI+eQlIS+64Ec9BHFhtZ+utTHcgF3ZMFeK1jGREJBrEAS9eVu2IpH094FEmHsaBX
PzJXJGuho/02lRYJOzKaS6q37WXOkbHeiImDsE8rUBTZQVBPc1GvLKl45J8VfxJk
31MmK88CAid3gI7R/JHRCbMi6YDY5SQ0Ku6dMasQknsieDoKq4E5v2SlkTRcyjmw
V4A9fqjGGbmJgpdMOHKgwZ1PEVdWl4Ccfqt0atWrC2uluIQji06+9pewKuTmIpnb
jNNzOLN3jg4DOkp8kY65TjTLcyguBX3R4nhjqff1ayZ4T/wG2/QII77DHS7kP/cg
5MhiyLVRAlj/+1szvOVc/ENAKcqBpK33s3SXBbiSCAbLDKrOsNk98iwftu0np1a8
zdVd/5djvpobbxK6pSQya9Z+vmORsuqI0SD0hBQL1VyzfM+9lX/ydKMhqvPn+ylz
yPfnK97HphQD7lfNR4dpOoAvmKvh/0MbK6qTlCBFapGcpg5l0q5JQYJTsOA9goux
aJkxdRb1fkq2DNhI3g8VYg3sxMnihVWS2AOtOPKhpoD1zHSY6mJfdT5+W2GzCCSa
olDTnor0SWeFHLJTK899QQWWSgkoF7DF9IzLCu2V7/UMOk5Dq2N3/1YfWRpqnxaP
MMeJLD1CiV1H4TIXABkJ+tgbLUUcdlf86gFvriiy1msVjd1bs1FfeCPodoUZHPio
JlaWMCe1WUvZaeB82hfv+uRl7HJLAAKRiwHA6FDU1KKHxoNU4d7A4ML7XbldNJQz
kP20IxS/Si6a9Oiv78Zweilgi/spWhlF+uJ01W7PVzczLZVOEBYQJzJgCSr/BzLx
9iWgPzWb/KjQKfeXYukKdrQO3/p15MQaYGEXoO6aNJYrYjfYYy+j0eGdEuyH8iYS
bUURQYSmE8qUCCYWYxP92nShg4BpgqbCz3CVuts+SUchlA5D4QGXNZx6rxl9pLUu
MNtyfXaDkpejzEDJxFyQ0P/JydzYbmJtq14nB74J8D8o9DfOsv4Uxl/cIDceP2jl
fCS2KEPbTd/biw7csVfbXdGx4fYdK+pUbGCtlsswECigkLELMDziXZ1v6wc470QK
HBQPMUkxT3KaF/BlnA823Fp/hfSFemlFYR8DnBYYSXtXUYwgZvrddwBHq0dES8ZT
exEDjlBj7V7/Jqqhh1M3DYRAKgjvb7lJMLLpthbaFHA46QBywMTHaYlOOJe3V3Ob
l4BolZCt2lM3qzPahO6ZdzHsJu8kaCvik4zWcwxde2Ne05ue/+2TYHyEIo6WXtM2
p+12yHxZLcwf2KLrl8Sf+F/g6sfSbCnH2/jAeLNanz3dgNkF34Dvz0LB0/iXg7L7
2dECCHGNPcdk40fVnFCVJwO4yu8/Q74pcrnDqa+IlOYt/Xz6vajf0eecYi4P2+tn
6gGeUwRbHszuF833VaIVwTQe3FOgoL/LvLjYyrib0dzonv/uoBnjq3QdpYlrfkvk
1W6NVm1zPhZjpR+xK2hvEuLVqwpEKyRuWuIGR97JZ3mpLRjJu1m7/DPihL5/NfPn
u3EViHXQtbDsngyBLmkJxRHilbCkyjha2IFYRLyp3kR2/MrN9vF1EzQToL2n83A9
cKvqANJTDOx4J1+gobpN8UC5abzdgCqNi2bWqywR6CjSWegaIaJe3qh6+V6mQFd4
kdW3cKhEvyjzW7Qx/OvENyS1eqfHLhBUm4tjUUzHfm0MSUCRGGYzJQwRPPs3mC3c
q5zZ3L4PTx0A/R2fYh+qJXs8p2R2650ScG1q5Y7kNfhOQiBxdn8J56RF0Z1wzsFF
v2tcOiWoZHpIKTY2EoMRv8I+61+mM4EmSO5U4HmFbp3e2C9RHD/tMkivZsyx4dcC
I0xpLKyHL39wACFRAAWfqmyE6Q3Q67LOMNAlJTlKXG0RKWKiNHFugQnaGQL6by9R
sZjOsVNVJ1oFZXn3I7QebiV5/HzRp/5oIV7TTUe/1sgR/tUBjWiD1i02TGhEXlZe
fpVhlEM2Mfr4zXvBSQD7LodqKrcYgwr/99Iq0YYb7xoN4VyLKdw77Gw17/wiVCZ+
naZKo8DTYUmnqvfFzygu95JFuUIwGbm89qixDGzIHZQXC6Cm93NMuAPWuvhPF9af
TQLcGhQYhpgDIpJ6vC+9gv8FIr3D3tkbDaj5i41FT0GU/dKRIg9i5pTiC053CoSy
e4Zzg2QAgzqKgepJTXwSgv/3Ew7bdqsuTcHcxp8MHwJQgR6fW+w5XFOOZMzpR4mj
zlk4LtwNrYBb3vuighcdj6gXgvZrxG/+imkm/cPO68ybRczQmh27Afsb+dm6vymP
XRcsQ6iGZ2ivpAeyXkHj5vsDM41xibshGZGlyr8SBXsAniq2k7C9LN3NZX+rp3En
HMv1LT/yDSu9IBKT2pKg9olSWSUErH1cZ2rFpsPuTgwfL6H/3UGgnSUvgy+tnXY2
dasD2YleOTzw320j15FWdkpYByTRBg5liWAnN1Nee5OudR7gh+LqkDmv4EECc/PG
Iysb6UVoJa1rehJz75TI8lLQKNa64MQkkAiRiaxzMGILiI13IN7D5mNbAyAbanDg
kFCTQW4u6/p3qdnvc2azbNYgGxCjqJGgzEua5hUysfvIeKrX8lkrm5nPahNvDzdN
YIhWTsa3eo728dnt/DkLm0y4RrMLWHNJ1+3cV7MDA9qNuUYxcsCQ+yPjmko4JpYV
WHBT8/8EA/6ykc3XdxMbHzZrXUcK+BWxoljSlsxqPPHWyxgLO3NJmbQKcWEEICSR
gOLyo7k2dKf3Q62WdLjnvnfy3od7J5avcxaySqD8Muj+ztXqeljQo0D4C/+iY/Af
LKdeUfmZSy9xC55c79WqazzXrzb309kNKHue6ikCsnZ+JIyhf53l0UKaWKRL7p/W
NXzGLqeV0Gk8wxI9cr08t3SOFHWkzRvNAExG4TDsoOd4fCD9Nfc42Ch0HSUltSpT
qr3oOgaQaP6R3/SsBQxvICB7zHeQYzOhmxTMvmf6zVvgp1MBNxVdVq9kt2a2O8XG
f5Tfl4MJQhjdgRDQ42a2v9J+a7gkqVTW7ymadXYDlWeAlZpy4wmMsQ74hS+mB48s
AsFcSPuyuY/qbDhwjOIg0f+dH0kN5l49gbXsv8Ltqvc4f3flE98zii3dVmbg3JTd
wdp3n8OC+W89zZi+d0+WfMFXPFwCIfu667taM4wj/sK+z3QxRZIjjXjuiUxxYv5c
FNoaX1u+u9EXBk9qVIKSwVJulPid82mHuV4orpUu6QdEFg+hxNrIikirmxFBqUwl
11iSjA/coI4zPt2GLPNmMpe37VfgCH6bDhsdVbyax/CE9/Ek9nCtIHat0cJ67Hd3
s6/cpbAW5qHIYEw1qP8bGC8vSdB1TMc4bLqu1z1bl+7+mtQttw7C6uf0AbFjqi0A
b//Dzrxrrxy6O9Vu/nwktMFsuysKM8Q3ErS/iqPSymQv66ER9NEx6PG9iEeCcBY7
0CSaydn8KG6aJUaSq/ypRrXTGxpMRS0CRKU4NdRsUf23C9w5LV1/WzCMt0rpBjR9
o3I2I0MB9n0c0C8kmE+cdE+29r7C0Xg7XiHwg1g/5KgGYHNBucMCOnU09oEvZlJX
7Hm/Z4l6I5VpYftYNSjGML7skIj7DaIS3ZG+OD6XOvkEDa1Z6z9jPoIIuhxpupDG
M2mexwoFLmDc1WSeA0RK9r2aXuiOxCFq8mjhxXmLMfT1GzrzdoT0Rwy5iKl3Z4Z6
Dn/XIhE2RdZ3pIhqTTSSVOXgpI9mk/4bKgFpcMjdsO1MZwFHyG6zUtsFcSiQfQm7
UMRgbD1sjnRRTnA/amZgVZ+ZQ+bfRG3ZrWjpMcG+7zaoKZnbc6+T9aa1MIimv+n/
yUyVLIyC9URKE7sdJOtT5+TXu9HYBiIQ+OqFptRiaG12PeGkJNLpK665C9i1uRi8
EgzVtQ0+OVMXsLwyk1GlAw7MtsaRvRBFddZ4anMUCMSoFhKkuTOkCAw+c3vXX2pz
oQGizx5bwKxBx4hcRm0R2cfMyrRWHpPIvsazyspXUeu5pcRORioKiEpD6HENKCIt
hdrB8FPBcUHOvXTlpzjolnHarqHBm3+ozkQydb3U5Iu95vyApEwz53aX17myTobK
C+GB7OvEswlpLMySktka7uWeXF+eli0dJ8baQaJqwUbya3PHlt2N2EjMOKtZpKkS
+rV9SXUUfMjvmeYeAIPnb0VDJGEABVc6ad7k/+aHOzRn/viqF6PCOPRrKZsFaoRa
i150kdYizv0mRAxcFeQzkK+na1CIIcm0b+0LcHAi2ebqszT7XJCQMCio+EdlmUfP
knVTkRL0CgSni88P3tjWTD4ssbHrDitmXiLms3VkQy733l+G3Uc473BkdI8Xun4l
RN/EmEe4hVKYx2qfUncdMexBY8CJKPHXO7EYEx2PnCo5EiGDg3TJzu/qWUmaIfGV
aowOXJ0BYuJIYb/rGOCLEW9hlWix1H6gPGzJKIFBw6/YWaiXVHYRJQdrI8xnAeK8
sIM5U41RgpCn2iGQUtg5cyxoG2kEwTkkTiyVMfn6PJMR1n93MJP76hwVI393H44f
uxKTPPJEycZY3WR+gccppKrJaxRikKm90TBybbhYiS5tJbw+ea3CS1iSGW01xiLn
yc2/tzJl7Jo4dBOH0X8N62japapqavwyKntzY7Cf8K6MigjsqF0SEkYw9rRNO/kU
mtJBxWq8/LIT4kvP1jkWrzqMmW97BNv7t/2VzL4LPe6+tbkgmKIyNecaqEvqUEI0
pzp7+RJ9z+bj1eH3+6TWxFnl8WKJZH2ch1UkFCSN6ncjpX98H3kRD2m0gq51i6dA
0vFiTh2s7FNuMuTCLNCqtpqlbz+BbJjbdsA/0u/qphKw0FP6k2b4StiQJTtwUby/
TwO2RMb81lzis0k+f7/Pgh/Tgp3WfEmLA8PbdXsjDPkxSExujmXoNeNq8/4M6SH8
fkeVQ0zALKT5LzpoWNO7BspPrSJjYJvMiIE+6p4ntUxdrEhT6IAVgZtbZNgakGz0
lgpJr7Tj/lwQyjJwtwksaD6sevizyquxeozC1gy7VW75184QL3ZiLRZtk2fPeTGA
z2gWCYXqqxBbtUn3BE7FlqThbEsrK2l2LKyi1IkDRkj+zhdPZTZVDyJiaUCMF2km
ikbiH5MKMyCM45udCFc4REIY1rnFj+AUBOfvGW0+sXdjuCi2DoIcvuq+4yZFe6y+
3H+sdBbA59esZqVP1+6uafiUn4Qmj/iz4dK4JPC0kZOQS5MexiLa+p7pFDEuvxUp
8BiCnMxga8UzVMirg2KgapCQpMloTkF5XyTypHSS8tmrI4qLK+O+RU6Gv+zHrBnt
EnylQu0epYzo1tcFkrZ1YqMu1YvdHTN2sh7ofi8Tya5QC735d99azGhRBqrFLeHK
PQvVBstPmw77DSy12ggoMrSv+n9C/rQhc/YDMRuuUwA6sd58FVvb4Np3A8xe8mcj
R3iCdC297nOq119w5RNip3omZrc3Q2gQQlvYOk44ataEJ0ns380BJH+DUkp73Hse
EXWmHysR3H8u9Z1mRWsYQrRBey4amEKvJrzKF7bqYzfiQEtfvWOAEMz37lNTAH0q
ScKdBtugmBUDRuywa+bO4oi4zJBVmXPCeznhDBC8OXiaa02Vx3uYiaFrlEs+16m7
gQINJZV5sIrMnzMu5J5bAHhyMh7sXJowleSXBeg1AfpY+G0Sllpz46Hgjz3scYMW
Kgp1azRQ6SWG/IhMn6Nw5bE4L1vrdEqMbiFL2mGftJ3fq7ngFb7+UARyccjlElYQ
I7Udh2ubV3YU/otL2u3/YDI1HuxpxDPWmd62AsaNvha5b4p7Q8kb0DH+fwm16pNf
zjNsFHuRYo350VNJ19a8JixSLCMZ1MdsLZdRKmiqe0VpdGiPi41Xy4VoL0wD0G2N
TERgFjtKnNtYDSD8DZ8arNk7/x5m4wOd4g3Y54qC5Qkgrrd4OeZX2VRqcImnR+CO
PhN77FCX7EEOx/U7od+ntobmPlgDVtjOCJp8yOeVAmBVFAKAtmGQZLdO7XfeLB9k
D8555x2HMeDTrh3cDzbZfDBOV6QXw0TUlVRjK0zsuxV+wK2LEcJVi8WAhKLqOGgI
3H1RuCjhI48hlGRliRTMlYY61yo8RL5XR4b1XA/8vVX4XZTQ5eZFbtKzwiTbbwWy
BecCdTlYOm6EO2kbIDOLWp9xGapUIZSgama6EQ86TeZDYzhHD5xJjTorP8hfGCR+
4Mb7WTZx/z8flhnbbiWlKnecHirnrXh2Ny+DqrN9efc9tAV6jTfZJ1hExoUboCws
l3CRFeWb/8gE1y15Z0yW+mvOciNQdqUjcK5r2bkzhoGv5s7YwAxEq0f1c/GtJZU6
Cn+IPWEnKQJI7/AU3H/skusthXrRTsTnmR3/saTn+ke4iLmZdhQLP8EQV4+9tK58
iVBFyZri8te4+L5jdeU4gttt1vx0rQvebN/ToNW9YXZ+4kfPaeYUypKIerU3z0i2
0hKhjaquRflD596QjFd72LJejMCvWiWZUGvMaxtYp+04DwcHOPwyrIWIMNyc3ZYY
ealLHnSKiSIVK4PEvcoBYYfkxETY5MMsheAhu1oR2LiDk8P5+9AdLjaStF7Vq3W+
QMHSJfBqKYBlOiWlGNjfnHZpM7iQS4kRx1xZydO2lX74/6rV17Ppnw7le6vRT5VT
UrDG3H3Wj6dadljLfF7guZcDKvXj9ZfFAbBk+3GTLDtPh9FIeYGJRY3+wTtqSIEQ
MwntxCVb23BncU30Eqsh/bMRk+bTvxf0QZwwF2bosHaIlFCbEYtRI3Y0vbaO84rG
hnJFvkUEPCBsqltENOG018GZMoxaktv2XUK+avg0+X6NL1aL/DMbK3lyQyWlVHlj
eDL4cpP1Rz2SkvAujZBtoeX81wNbjzrIxM0Yz6RDymYT9Lo5AmsFPx9EKNTmjUIc
aCKUk1FmCkWAfecw4wfs8/vLDl0XrdRHny5aPfZ5Vcb90WxFgL8jEapUVpXxyn9B
fntAL06eBZAOr/I06OA6Uoa67gbUBpZM9sY7NK/Qolxn+incZOHCYpR3+AF/C6vJ
msO+0kGmXhQLONHmas5D3SLXNCNOd/c3jkr379ObLXwDs6D5SIizBSh2jKx4f3em
TgsFHfxmNNczfcEQE2hwX/Zd022mHXwUTmqqtv1SS2zyoSj1vBcTYD9Tx2F1Wly2
FSjImIyKzKN0YAwREsIfopuFT0rgelK/RXs7GuxjTe6toApEjnFPVc54VSGgvATp
zgPNfhtYwsAsD/GfYcJ7wIsaGrUzWVTLjfV4sx6F7LYNXYKEliBZ2tWkoQ/kJRUG
sy7NTswYowWwDE+/BsVSitqt6ebZhNdRbSEVGlPsxC08fyRBlDUB7G6llWfClbtZ
BJ8WUtDbBY6dTPr/SfAIItKJvkfLTKueF4rtXyN2MI2gEWkSufuQVebPR7ah8Vut
xp+12ZyhFNV+6ERDSfLKMVVCOQhp53nHZF/BUoDAIp6qZCDT/842RFBQbuwxfQgu
iyuRVfZ4PRyC+ECjBIbvGZqPPC+TV64g3PNWY1zJQ6/mTPG51wdT5okqb8HI8Hbb
8eyeDcE/N0enZDA/YEuqveBemv3kJoABjfxhdxJjbDD3C0u1dSvL9JbGlYAcW7RG
3P+K/0xv8oEup40q2097TZhKQOXcnmZVGrGXhg642wGW6jYyCMKbuSpXTo7iGgti
SDeenMm/EBrwgamfSuRmKvWs+WzxwhwEkmtoBS0xi7WloHwOjMlE/MO+JH9FsBd/
Z/eGyvrdTI+qKSUq4XAuYc64kAp4qDWs6qXbNyDHlkPV1j1Dn3dFH/rv1x+UKxDF
RwtsJsNEcZ0fIyVlC4gFTU47iUyY5l2iYWjwgMeG9nZPpQW8chge61q9FV26+Ldf
WfqZBtpoW1XJSAIudK1j/2lGjR9swtI59GPStCy0/TDcParxlGk1H8jlBAPmRMHa
lLXwW2BX08Q1wqbnJK9lGkpFshaiOCJCLyIaVkGM2oRrPXsnWMcNqDEVLH9CVuXI
hNpHXDUW5acXzcV2TUnbs1qy86fIo2IXaQKmHd8TKolsIlN7zxo89QfOGF9tiWPa
B8iBBFx/g15Eq7OFTr7Ws+55bra+2O6Tqu3RglRqaXBpFIiwZq2tc/it8wEp6mTP
jjYIxG5Qluc/y+ihMY3gCHPR5IiF+tCgGUyCn7MtLOL+ES0vZG7No4P5gCui5pDp
gf/yFNNbi962riBlWds9A/5uBgOted4ouBN9WocuSZdI1mvXqcdhQfgx8SQOujpG
Z/hcP12VOyy2KvzPHUNNADAAyt/UO+sBRj2zAQUNJPfGteWDuWIaHCPHYnaN8ugk
0oJDMqv4ueV7BvnECrTFybFrcn8uAIytaPA9oxlrZ0hu2TWpIkUmFtCDtl5lZDJ4
TM/fe94EQfzhgKyytHN0dWYx9e0snoVz9WejODalakBDDwRFbIefL4M5kyT4vaQC
v4YT0+5Qr2ggCwHyEnWOe1WLw626UcpG/7t6is7yv3l+r3QBUQyQrR0GMGGkb58f
v/Wb2kIxxRFUj9guLCX/D5ela2ho8+rKoTqIT5j899BdhSWe34/qgsWdqGgF5T1d
cajxsMEXEc8bvBkc32+ZJAWRcG59JXYlO8tYaTKwTP1sWfx5bf9/ejsqQYqtrq5E
URQbI8BcWHH+zUutG3TgManHRAIOAbOGZ7QAOvQ3CiS5bz3tZG2mIvhspPyysjd2
5LRk00+uutyaxf9aI+aLBbmpQFAtDIDxN+Lp3JyruB8DlKuZhD75oEDhM+EBmHQ7
gENlJEcHgyTKiVG/UkExTFUK5wp3iFfVSe2jJUCS8DCDS2RykcAdS1gC1u+JZ3Fs
4VuM95EWUOF1plxh7Ln8tRgsH4vsH2Q7elREx1vI46EZ2jevlCjrZzXZ9GfSZvfi
TllbE8JqR80vNUy/5PzpZ4OgjSiH0BQvZLyeQW5Caet3rR3m32l5uUdOk3Wb6THh
OD1fyj2XmB/GV+7hNre0trUMc/MY9fBz/Apo9H0AOvv4GEgJ5NhdSeSxobZxdceA
ZmXuZsb1CihOKdscvbbmY3r3zWUJTOQpuhBXJ9pk0IK37Khpka5iNYArEWiJoPrY
EqLbXb6clT5eweFl4gC04/VKbn4ywE26ZR0FMD1ABnRlNS6OELHPtpGt5N1sjBHI
RMlsTVeX0Z28mPb4BXjZja8FQuaJlO4ZqB44A+hni1RV+CblighwRcsicM1ZXT0I
tykMsjJUzxSIs8YdoYC+qitinMCiRszOa2LsIR0SseoU3IFZ8reI6D2TFn/2xSN9
8UwFOib+3bnA6fkkv7z8bShHIAYkUaskLcMcZ0wvUPJfqm9laWLObWSK/uSeE/D/
LUeoJi21DdsLkggUctPzAOSFlBwS1GxFN+0NUECw845vUQJUUu8TICCyNcGc9oD0
+/M/g+63ibu0OyqmSPWbSHMCcOS1UE9696ge7o3ZWrXLQqVunyk5hmCC4GC4+BW5
gRze/c3xhjpelRoyotEWtc7J0FQhZPJbCUL4Kqn959BhhO6SDe6rOc3/GyXaBLBQ
U/41LAxy2qvZigQjW+/dRztJnnkPgXDAn70FzQGFG0ye6fv1kEHiRbJHhp1vlDw+
Rp5WANlQQolUDaqhCT0s/kE+ytsZZ80ErnAptQK/XFdrOG+0dOgEF8l+qxg6IIQy
kuD3IFHYxhUx6ltPIUDyQFxi7RWJLEAgaj7BQTO2n59s+A0118vggRt6b2S+qFLR
0LvNWsNcddWvvIH4iALGTmAzOtLVfjLQrVlaRjokgRacKZWnBLUqOB4Lt7OCodDN
s4G4MBE4kAnuwQnJHrhmef4RBAGFKoqCzWrzyIzroe63xcYQlb7M0enm01USWURO
VEiDJ4w9TQjf2A4amzMG1zJWJ2C4olKcOC79XnjDSDbcAJmmsE9dB9qtAAqUiAEQ
5/jjgvcpF8XR+EqnxNEOdXsowWIUlbws7f5rz1HeI1FYJWk+WwbKAXPPh2gTqDaJ
3C4zqo9MjvZEXJBjM9N/6yF68nE9Ebtz8lou+SXQOu/cMMc3MPJZzgcelOM9bbuk
CeDzQCRDoSo7Lc7Z+lnyidD6fZY8GVwU1wUb+XQsZsH9vszgiAfEjA/Zw3lEkbvS
9BQzLS9EEP8zti2YK2JNb8a9b2HVL4X8ruotxW4eODpjzwUVTSiFvgjYkUgYmQK7
VhoTkkTYD9P032oBAzKF0qCog2XzKJnE/rHZ1jvxktuWsrgyRQ+HpFckuczH/Dfj
DcJenCIGT/piMLh/lSeIJs07oWyG+QxVXvPpfwTLefv8pBdxp2wC1hMyMzjAYBVS
TjWYmHtS5P4oQbDbAWh4RjQGKz7STh6DYK3YG4uXucwK9d/7GnDvpcvODb25d1Gg
FZyL8Gawx+XFHRmEp/pbk6EravSM98CW7TcepGXt/VeUi32LZsPMPN1QGPTco/oE
FCTnUhK1Q1DPa6i1WTdn7ZX+8qhUQHFQcj5T4tv7oTard7Qzz2hPUdBZqbOuxXmj
8mM7MqO0a44wDxC9UqTrtEeYypmpIGRcv/ZtyqG6LBu5GiFT4EMT30CLva0Zf2oR
0VY3GA3Q2gg0zRXgSN4Dg4pqk/anLZlfUfu2fnW69w4gfRAzOu2/drBukT9/tO3D
gRQprMeIUz/nVgJJYL7X5JqUJXzxi+pZDsSQgfIbRUyiDhXykuAha5NasRt5Edg0
l3Qmcz9x6cFH979WpcsECI9g4VzS3W6cYJEnsvuR/q/nWcqUvYSNWdobRXxmB769
QpPYpVptZXFn+YtNRkdfcDN5suRBFACKj9tpA/0bcEoZwc41vBgl9ezwXhXQfTQC
HdRkNZV8nVxuS7EeHhi0bsaIhStgnZGwTJ4aFTQxNJYmzdntLSQXknaoxyFEgCAn
F0dFzF5UBJ+zGXVTubTMsnSiNvqrUwVvipV+HI9L0W3lP4qIhVmpM2MsmzTDiiIr
KxxSCevMXbHc08L0yT7dmgfcHStrLEODatsugk2U10emQRSaOIP4XoOoSMITvrab
EP3W0PuSTqoluUrEtmLi3yCofKMv/lxXnGA+inggxE5FoGlmV3Xuo8Q0qc7/TUeH
suNx/LsmBvQWgtGqA7J9FR01NEyNyjrmiKy9i6Q/PqI4VwEcWOwXeLuAyKcD/eR0
jf8meHKmoDNxOku0IJcm5NJ+vJMrn58wCVd/d1Kj3MaERJnEDbMLslvxBx11OcHw
G+3unvo4FC1WS27dza8gM/RBmE1j4iZDcYQiCVt2efjgaSYQ4Jc86Q/DOD7Ck48z
tALmq6cvgqYPia/FdGpKEFNDhr3YHuk41/RvubrQW9iirJhHRd6tTwxOa4xJKAnK
utkPMmn2b5ho6MoUnU+2oodwB75bFNJFpZzzbrrAXI8lYmBQWtfS60vrie8Qyvbt
dFsS8U8XeCLzbayE9N1XnncgCyzOTbCeU9UBE++xmILSbDPVM4B48kED9STva75X
ofAjibqeNfZo3XRUeUgROEKRYjnAUmDBsmRbYfC8ilpcIe7Ij/h/IuKwB+7k08JH
o6eyxP+4QxIe4lOtpeVE3t46VDGghEmc++aFw8nSNBp+qP21F67dPaETdY1wgvIJ
F3lOO2v/TFloFGQ7ZDx8vw+QydGqvtYG0wKgubJNSOsJJ5CdSq2ClP5yB1FHmCDR
WRyH+gpSxAezVjkdlw29ntR9gK1Wxw+ulXkhkUeDAv0GvskrABTup+dGOX8AfX1p
i3wLlSot/PPaBfGtQnQuhk/Fg4lWhl2os9LBGKkQm2QDHdo0tvplOlcBsYGueuaT
S42kgIdAjx+sfB66egCgPNwJWnH863Wr8IEAZuI9YBVbupfP3S3bdpNuH/3qwRyA
5r23S1UuXeoZR9UQ5P7h1U3uJvce9BtvBLMJ6cD23lABtkiUtBwLJv7tfpD24yyE
WWNaWsDhNpp9DwNDhRW4x+d+ZVcdrlwSYEJ82DOHteCkEVhFjYLSg884TITQxGCA
q2XBLu4CjQ1XmmhsafKAOoQMRxuXu19vm13ggzzqjt336UDvPBy+WYBMZEwdLj+s
FIaAad+dL+f0Twa40SEZFUCydSRmmcW1scerZfJnlSS33N5LFfphUK2TCBCyiPIm
WjAEo7elNMgRb4d9tTGYqzo3VRmvK+e8loHQAhEbySNNQt9Ne5SS+i7HH6pD9CY/
AuH0175LT574cM3nZziSaldFCarZ1iMRI2usbM/iLilNPgiFNIRwFb6M17t6K4m1
nkeGjg/1zACAN5cu2tzS+wWzAooEYp14zA1ym6sSja9pf7Vfv4rROoLNVPB0Mf+g
WIEOZ/LC6LWP90b7wd/9lgIoHYOVjvm/RyhypSLX1lzsaVKi1MBpeaHC37rfzze2
hlLmgEJN8y/nzSYTYLPaMFLbDV7Nv0Qo0zwRNlyG3kFDD+LSUpeBkS93W0vTCKeG
IkJRGWllRKwELsqfSbTFmVyx6Pk04jy5gThEMwBqXIOK0brLoQcRlkBz2u6XOpr0
vrDrgp9fVQwuIDrzMi2D/m1DQYDhI/FP2H1XB7/nZ1i6ezLF1hHsFDUXzYK6wbUO
fW4PLf1udULmQWb3fDmRLC+IBYDHtueJiJfhP+T4pQE0qPSXMZwgyHhr9wsZRdb3
8PrZXPcpIUQNOv5azV9aHFWvMu3KJq+IM6NyP2ETkzoPUOwJwJmJwPQCz1hPUb/f
eYf0OKejguqAQQpf23ATkZhX78nYVriz3IM1YKwZF0qUBeI3NTZQFV5rEZfTETKc
ohKQDboiLrniCpNxip81uCgbtvZShNzr0IbI8Q2jFw8mAzCHEpUTCKdpRxvnu4yN

//pragma protect end_data_block
//pragma protect digest_block
ShQSdh06NWtTUICnS+Y8k1lBKg8=
//pragma protect end_digest_block
//pragma protect end_protected
