// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:06 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EsGMQK/zddvSOLlxLpDxzVwUPWH4+C/8F2PV4Mvc44jXl2itW0RJfJQHr47Q/tQM
rYxpobXs6qkH31tx8JVVd/MdmCWuwsM0dps76rVaDQ+u1JwzdcCvi92ufl/wT2Qg
xz5yuS+EIDmhDp3XsiVn7cMt2Rvc+Bp1XrAAed2cl/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29488)
VxHII+vDCX3T/CpVZmhR9IJxqZ5DdexFIQ8e7pbBvEXMXv+Omkqj4m1uJXYuPppS
VNvrNdlmnyTn1v80RshgdaTS32/89B/pX0o36t7uuExvcaSRUx0KRBuAwstEAvXH
NJELm7+KMf0h0ytDazCuWdBNJWvqEpL+Lk+srG95zKOOXuDuxdyOBx0V4lwMG+Pd
4WLheA+Owv7P+HslrjfpeX17LOKSPp28J3dqzqh8yiJxwFN86JsmmFO7+UkZP4u1
WSY9qNNhtA8RreId1Dy5UF+Xq4WpseJ26qBPloUIOf/xvLcvQGM1tc7of9ACnkaS
imHyiogfMf+zzhcr2ocbMZzI2JqsmmUcSa7IN6Waoa/+srnnAEhx6+wyWpXncZzH
5ZeZzFcgkpzTJT6OIGTmfhf4TL1W21+YyKV3UkSA4ch+GpgVPjvJO/VUxs4nNJ1g
KTmolSzBijOjFa0Dvlgtnx1BUDL+cKJMMT7DV8QlxkGT7S95BZ5TqhnGRHfIAG54
TK1a9knx4eYDOZSY0Qmru0E6A97y4wiT4mtONRXcaC7F/Y5Lxy8ImXYQILwe/Rr4
NpEfxqHEOuUIljtqMV/IgQuM58I9sutB4dJGdKe8UlY5jtTNYTGCBe2X7sKWia8E
vOEZnuu3gBxtPYSqpn4Zg2hR6JYRpdUw+b3+zQsIHz7R4A7vsYi39hLGtZeNlNd7
4k0MX+pXbBp0pKB1Ib34fg0v6PL3nec16u8T9kpDFEsFkTsCuwbr3I8CCDO17XdT
YHBwMCYELQCHmys6qfJ07dzDCjr8Jwmiqtzr2qMtLP+VAZrKpDNNVzzgdD80fxst
+VrHBCUNRePW9igJFp9hXRiLuFxBZS/q10FyKCKaZ58bAlLw1IT5kfdP344W/yDA
RKj2LdS78m8+2wO1nXh3M5iWfVkncYoY3qeoTAhkIkvMWN9+vzhN9zwFPCZ66qeX
kydy2GrMMLFAOeskK4Mqr5X5/4WWhlXV4CuTEeAbkDQObi01QpSzwAg4C3YIsXHE
i+pPUzeTOeCMySTYpl08EjXVw3iWHfqCxgcKYnKb21BqUxipIAVBWaWdDWKxQF+I
Bx7vTV9in/LH/eR2sH1iFtMx1XkAxu0vJ9k7TvzRJzEibmRz++hqWmyuIZVwxA1U
pUAekWUDIWE/ELfi0SYPx1hz4iMNmURkLt3rePQn3U3Eo0WYp/yNGhPPGMxCOdQG
Id7mWMEJKZD8p2D4aWPL92qBQmqUz8k1kVBL+ZqOwsSmszd71wyR0MQ7Z/oTHhxP
FV9xaNaXk1iRtkWP0uTg/jL2cfh+V0SUkYop6Gz6ii4lHm5bIDCMDFfQ/mAwaYla
sKfJJUN7u5OIA8TKqFCKXk8RvEcUSJwO46HUxSUPqAxc5EHiSh5zlpwzeENvfXAD
CoLbPydDndH3L1zYbRaRHlSxwntdlGPzfIenZYp9JyWl7nJPasm7bi8pePZkKQgT
chVVDnnAqFB+JWnrfJz/O7ZEXOIaOD0dGII71no7K4p2vtE4VR/0jQUkmCldXqF7
cZNtX0DtfBwbYSFQtgmbsFmMPRIPAdBL3Qhobck1p99iEo69w3TCUDuBHgk+nv07
yVj13wYITyOve1FyIEc1j2aZe2z0QCKOFGs1DjjEMh03JfUHnC6jtfjXSrZxbLQr
ppifJVnUMbljZBrx2aC7XGyelpb+P4FZa5v/7ficj1FhG4gauLKhHpFaT3TcP6qJ
ZYBvZ8wsUX2aWBG53VCu9lCSWmEXMa3lx26X8920LxSq/2nSM/jxefV/YvBIerwJ
YUVyNv5prrrf1FMml/+JKPM5uztVFvTuN8rkhMDvD5k0vqNEAeoqxpCnjxge+ekB
zLgNXxthZKeMdqM2en5g2w989A1OFFIgjrtfOZc55lzpsbW+h861+Ikq5wYTmEqg
qkyOEuhDUXOeKU6dJYPrGW8bTMO29TEZPpWPjg7cXafmXyx50I/O2aR9+8fZ6chB
Tm6OhyW1FIOqU2STa/vWFiWDIMEbT7l2UwZHDZjvoQEFY3qlWVZrP3E+GIccTL+U
aVUl7tdEmcRel/Dg5mzb2HYuTdcqaEwMtIw5eUGPJkInjEErfuw+SWXKhx1Kd0pO
Zau1jMmgLpQJANTJ+GaEcpEcgkdo2+mkIkDsrFA1e4HiNaHfL2ABje5LGWAxtgiL
Wwqq2vC/+tc97+8bZA6VqQYPgWkWb4z6IU4s9unXUHIHL3vmStgWfibZSgq0TgSm
AGPnHZ5PE/p6eh7DxG+4+A0aZF5ObnYa4okgQimbOZbphcXbGiJ9I7p0cCbPnx3v
S5S3Jc1i1/WuQ+I0buKh2ay9IQk1lyf4GMFrtNqeg2UZLXbORWFo78vhjVwJIVPt
nqS4g2SPxwKH+k317JkmYWKrfFKEdpuTK8hwhwQ7blG0rk+/ZXpoe6IwDrP5xnEE
jVTlulrbeFgdDAMcCP2+kw7T9lSf7jVh4+nxSCPECZhXlyXNUWc6LLzTy4i6cfx2
WqOlAHcsygt2nMkxtTcv+7cxBpp9PMXNTEIEb7G+ysf6uU+s6QA5hDw2iYwl5jW0
wh/lQfoNQ2h0V3PIfrEDM7N3IMIsMApJ0WL0SJS6vISl+LUQWRcb3F2RZxhHVToh
Q/eAaKKU/ftcRDvXyeEvSYSdlBXV0PBrzedg8Sy98O6prpflJP3/Dtd7n7wnT5V2
V2ZjEWveushyetJ+vndzKTNUwpnpfPmF7BUDpQohDPLzc8qcJ/SoKohe5tFROrsT
cW38v1TE+W6GAtIVOWndTEJWwrQiE5pcDZxdOFdwB+/1dRCbYY54HKqnfAmHZQBc
/31C2qiOUHk6qUeI2bPt0mmYNkEokhRh/kKLCp+UY5dY7wiYGDzRwhl2yHkT8+3u
nTWZbrzIWNWHd/LmnVKE3NTrPZ3im+2EP9d9EcXiCpzAwRpVpXcMd6Gb56qiE3Ja
LployUCBss9qJSQVbnenhJ+jGEss5b3qkOSvnTtq5HsHoUZdfdnXD7sp2WzhX+GL
lxS3aMsFNgKCyE6Lg149goxkTlPobjfsBWmfFKLQrzwcS8wFYAGJvP58f4q7QmZj
mjjjKYUH+MF4oPKDK6XE0Iox/rkleXEJIBtsDsHHYDRqH/ZuYKwRw3SI4rkOgA8P
hlFjIEMhPIhl/bCZzTqSEs4BhGMQCkRcj87KIf1r2ir9VwdxanXjvKB2U67O8y5I
Ig254aUIMsNlBKt/54dGMcR/ukxdBCu5yE8BZcKSbVhnbwJ2z7aHe974t4nS1ryT
c0bhESFW2b4jPRLTPM7Moui3uXb0h0b+7gw3bUY/ejzCo0uzV5vzpGTkrYTpnbJB
Xn020wZd2PKDUTuES3o+E12O5zxwhejivyghNaxjRDip7GdQNtqzMnwtoMSpRTjt
GBJ+W7rJKF+ods1p87e6P+sCZCglTrIU+ElAEsxcIjCXL+VTryJjE1nRXLBhE50g
TAkFZm0YmjeQsHu4WvlC+FXRq2kHhSLv/C2/BCPMZHbl4RQbC5wPVTt/+T4o2+3Q
EC/hb9dt62JBSG0YPLMBnJctXI7LUgyMYHaU3tyoxa9z8dRBIC/2qjmadhy7X4Kg
xQxf6/PgOlc4zQ9DuzY+MSHXan+UMWTNLg2/DeFkcQcn1kk9UG+fh9ssDgTDnsL6
yiXPr+ARlCHuIsIzr5qXD6jq96xWZ8C9vyRLf7cHJPi8bkY9lzLBoUr+k0NFltIU
JLAcnv81meEVCXBi6u+clls9neyoE6VdSS71n+wSbgDwXkZVHd4MxMJ8nZHeJoTr
TCLXbw4HoCKkVvtmW8F8SrQ3sOjRDTZwSVrNhn3nnu1I18PKCyEdiYvo6M+15kEd
xnysvLKSSu7PCk2eXYuIIgqqUs8WsCH35I0ZdppwHfGAilDswNtIKutoBSTsb9SW
KxqH/xxtqQob3c1Gbgp1KPFsCYWz+BLCbDQ6gZOSnuejkSDwdotuhk6Dn+ARvUxv
NPlUmQ+xzbw/4jrQoJmAlOZPIV6233S06ZlrjpHtRKJA8DvNQECj3zFN8xDuQ67r
Cs1i4yW9ZCTZOd0wefZ6uOsZPZc3KsJZuDqALc/WwZO8pK1GJIwYR5grCQQC3r3j
B5r3tLJeu2DpbFME79LbGmX5zBuFb4TMlm/2TLphETvVw2Alci3tBJ0KLfkELulh
UFMmTCxDgl2UX1sE+mts2F1CrEf60vBAmBbNZnvrZ15oIW7v+BK2zqcgQyZULU6U
2WtymTtaQHZkcyqTo2t0yXgMFocDSgf44MyCM0Wu1dKtvtALIeyr8EXWfLxBuUCD
ZDALqp36gnTtIMRRlNT/2/FW6zMI0L1yASHgo5uagEGvLtRvpcajTyIxmDCMT5BH
HJsMxK2iFLcRtDOJwj5qMazdbLhOz0L5E6jFUen3sWplsIf8o09f74UhEjt3ntLk
nhWXHJm9raDjnEnl9T/ZWcY6+ulh/CtYtxcaEwEbCM/bA+sK9LEq5MAQ4GSi/Kxt
7YY3dFgH6jxN854u7CPuwOpR3iRovfXN9Ll7j74JpVQSjzoCImMSofNfYbHY7CjO
at5qLrPMJdYuMJmqNHw8JcONKBzEZ4WuOKssFKRMrDorZcLRZ1Y4XSbk1UE96DJL
ePEvmYW7RR1lnd58DpLJ9mWvUsbr4zUuAYbD5Tv7+I+GR2b7n9AVULcythtoyWTX
aLA7NlOSkju9v7qJr/WaLW9RDM0E+DOMMWeNOXVcWan/s6YltZz3t6Bqr0QWs9hh
kyBhRrvsSn31YqbpSqwo95QaUfbsg1NVReEy1YcM6ANTjF7F+Ne3uzF9SVD8vSy7
1WAV21WLUnIM+BZX+HjEGuNNpcwp86JFbXhig49IxQ0bXyIialBI0F6+bfxLRjq2
pR826SLpG6P0x1GcSXH1azql3EMpWepiHmY66p4nhYWp893nrKY8Lsaack9Nqc8v
rTl/BSA2JnraNvOAD4j+SqTe/+okJ/HBpscAdvKuzy6sJbhm07Aggl0s6S5zIqPB
SOcUncGt4Y+wbdw59ezLopp9a/YUbCGK8ZlLC2RU6Q9CftRbYWs7D56Z5a23wLJp
eRqB/YuOi6aktz2n9rmkJheOSRDC7JsMi4S4LTHSqfqZ6oRoBHYfKS7n6e3FTqiu
+6e518MrQhaqni1W3Hj+Kdttn+D2xoDt160MHAYALgGaa//YO/tSBwkUeQoUetik
/LxHIvv4rxwtNsHA55owwdhkC4/NKs7k54ykHdyN6UxxDgaj9jP5Znp08YCdodTx
kuhIA1j0IK0ZS4Fd6m4Rf3YxE+yBOBKtnUyog245wwZZqi5CaqYC2j0cFwr4l+KI
4WvDoyhrQ+Gu/xRl1q9GW6vJhwJMs3taMEN0S/sGbLoRPxDlh1IilkPxc7UduWm4
/R9f5P18rJOoeomCgYVDGD76LjGs2miZrIJuMWV3cV1ADvGkcpEyQUs5iUwR3l/h
XRvnSotDIWIsc94aMdH2dcy/aYORtQHNA40MJpM8a1DPvgs5J5ajX0iWbO2kTh8I
GhmGtYLHFLoYfXDpMCx1qlP7ohDizlPJ6mUh57wGS6ZSS64kacw9BBM5WWHisS7Y
hHK7m5NGCHFvFii9rTIxIj+DlkAIX6AiTj2lEqjofitBw2KPBhMqvFOMh0ed8GWj
6FOV7Ld3qCTUw8gYiWRNqQU8VlUCMhMlI+Kzb6H0VjID/quZ7t3E1r+HQjGfJxHU
rTdUuCjONZYYD6vvLj6PfYX+VvlKpra8lc2tzjZyrjsqZkeyddWW71jsmKNedh6y
v0uG0JpYl/fOdSqcyLHB+/cDxdy013JNS8NUhacGoqO5rUrViZW8eB84UrJdox/M
LN5c7ht9kvIc64NGCG8cVnrsFHrEplyxMHzRTPngvtb0BBANgPAvzC2dosGbQw36
/OfiCEiZLEnqJTbyFbMICTYlDv7fs6T3LdxmoBidumtUhe6Q8xc3RMlJnfi+TmtO
HhEZZuF7Cma038tgfx5Lt8XOA8k8Gk5RG8Pgd22ry3l5Cs65lA6y0RTxxO7Ek6KH
Zm3zPAqY3f8FqQl1SnW2RdPO2TcKQnXzShd9KVKRmqq5DNDW+RNNegrk8stj2KwS
Bnzt40MQmoW7Jk+8JQdeuaiz6oWVeCvPvmbS7N2cldVeqFNYpTa0ID3MI6VWCufa
UQmvjHp4BaTjfo38JZ5vxs0d+yk+Iavju3r8Xr5dANyNxx8SZhN9NES4wLvjgUU4
V27lt3bKJYu1H4q9TIqGjzEK80ypVHL7/I/iWDd+5nauGPmRfHoJGRV3t1ctte1X
oHNPYk8eIhNMW6NOAsS3fIEytqPohDZMFqGsm5CV73Y2yNWavWyhbN0NhbMfKlSm
y+dETKNqv+L6MhC1RN2YIe6vC8j09g29eMtJH054HJbZBmaZ5TrQezNAM9gLUxHN
3czPWQtEuiy2qRZUDkSrZZTZpt42RRje8P5mg75Ev1g99P0/JMRu+fJyhVm0D4BG
tLB50ncQu5gSmY1VCYluLg0BhZe/04woOtLRuJzfEQ9je+QHI2R49o5XzoKn9khg
w11X922tVII72g+vvdlrRddR+/kQBDmX++VMtypSu52qmCac0eEyuKz4UrpikOLN
f170CmCEq1BxEnriO7aWFCO9oR2rLCwTAMZRrPDX6zRwIn6k9HtpyiJ+zoHm9GVh
fWoPYvHS4T+Oer4mr7cwgpGUCQYEZdj0i8wKd0vyf3bV5n5S8y5Codq3WjhN9GOz
ggIOt1FAKzdFqwxHtUV+ExEQ6Z+ZAmQEEPAfrWzmqcAt+yXQAJaSbGNJIUZcZrnR
okZWR7dp5t6JwN+ndkVo7VZ9KY0K9shZcAA+QDM1rZAJcTFF1okAzWA1zvbuZFIK
8Zuvi9qwn4bmHRcyVfcECfQmx+dCP9yH/pOiQtJabC+k9rE9ovNy4HmOpNDLQTxB
cMU3yjsAY/d6TrsFXafLMKST9X7eKKlrtHvb9kiSpkSc0bYJsSBRk+sfNHADZzxk
4HhxOjWAq19ejilMxnOdtIhMs4p81uwqCYIWP/l0FDxpUYu8EidQdQ+udbRywLjW
c/mHv5f50iB/4owwBCCHB/VPdnukrZUAb8FJUUQj+zHX38G6YwVkL7zXbv51WQxp
U9EkjSl6264Nzc/6GDpwu+TX4NOT8FHYPdinMdvmz2tTNHN2EiO8b3M+o71t3vMX
Uv9uhujYg0xXRBG5sBVXF8E5h2v8gDl/qZM1Vh2DVFe2tGyyNhmKLykyWP9SxqtR
jye1xvVlGmReLOghSMobZsl5I3+0QTdUFVTgQ+dqPnsQSCiMD6w3NvDRNZrve7sE
6riRV1xhHo9kOKnIRiBakcO9QUJ0XyOhAjyJVwBXdx6UjbPyRxLDPR4p+JKV/Z8J
SZgUpQlhHd/Rl1ELfzGpHRIdzifJfBzrtuP9JSgsv8UsnJqnQGZLTNIzm2NMQ6WT
9MdqxWinZMNDOG/TDa98iH9lSPRJihw0Tn3NxanSRFPoKJ6QaqBEH9sj7tiDlamn
cFSJDI8NXEkUtE/+cAbdD8OhmYpiYh09FzriVt1hoMxulxsXPn7IDmLejgVNYU5+
so6cjPv2tKPzvxdY7WwlyJEBcR1CpieO3/yN5WC7yf4jA2Sd173WOmWFIStoHOq4
jL+i1kWFzPDf88ToZG6g9w4KgbBPGSHipPa9kIIqVwn6Xbn0PHKPsVxwqGprwHJc
y5mqhtenThipD9TDkwwrIuHSYKulpiRzHq5NfMn2i3M1t7m+hURfb7GdxyPCRin7
tmArzWtUvrwwWsW36a0j4mOFwLb5bv77xf21CQe3gkc8WJPs4y+KXBt5PK/7L1SN
C3FukHf+TVhOZQzAcz/zGPvxZrosbg7UF3QYqwAerwS7VzVRlATAhwzFnkW+6Yhc
Y7Gfx+XTvPYhy4f1BaEbdrDytz9lgQr2nwQqO8Bcz69tOv0Ke0vUeJGrBFSNyqen
u2HuWD1uvqNzfiaf7JxmgEpiuZPWz1UQ1ztI/qZdSP/A/r3m6av7Hl6HCZVCPn4P
9eKPg7Zgj3VqWrmlKoOU33toOmy/lmPRA2MzLBjCwclsiPlFUJu5dBSt8HugmIxT
TS47ad/bvGG5ZJSARe1AZPn+TXlw+iH7e3qXKEXmVslksKxdgSMSB5Xg82NGd8zo
4GInMBC9o8WtH6wHs3ogG/VOnwA7ia2jWbT9ByNcGj++y9ZT5qLQJMFVsy2GwyYx
ES2R07DfS0wHPajcWbP+Y42dQxM/p0OnpNSg1bmVA8v22Rbeg1FXZL/RMqB0/S+D
bDooz34lQUbNJal9+HdryuR4t3FPVWIpuijZmDFhhvtbtHQndtPA3MG5/nIMvE4X
l+ZD3e9pBrkOYzuspDw2tQ/WTH6ToQ1GkY3kbatL2IaaG+UNLyitxqKR9PO/g4ro
87dnHcF/4aKNnAK8djSq869NwzIAeSqCYQdW/MxWKLLc1oC/tbiP54UYaISvi6nW
LzoTjFLRwdPQmYLfsAnyxBCH6Jj8/FM98YZfyPcCbMStAmyVkfYht3VleJFueOUg
E4eMZLLPLbN8ZbEHT2z+GxAQZqiY9DSKk/ri3uMALlGSyYggsCr3G6EQ0bhA3+wS
8YrAd7c/z9q+FXWZYOnRyUh8LJeA6NBcyRLcZ2MO4/G1jLdQPEWRZFzrqp6AK526
1IDrunQ6VkZhMm3RDDTDgAI4Cyzf6avurvLYmtNXxN6v/l+J8g1HdwMOc0mGmv6s
VwUniO/bxbzPBZu7/OwtwIbIasKqH9rnEEq7p2k/+2l9upJ8DKJdq/XQvmC3wy3Q
+b7gkWsPxu7P8UbyExVVpdNbU/pdl9Q0Yi5lBXm1pWAnyqNIWjniUc8h/ZXtdG2a
S7Im29sqM9HeyhwfSGf2I9u11FOcgQz5WhWo61cS0T3QGTvz7r3IK0eKiHQOUY3M
EDBoYH3wjk4n8tgLt1W14Sr1ukJw6pdHCp9uirpjqFGsHsaWQwAAPaA8rEi8SVsh
NuEAeSHmCCq6cm7VsvB9GQRZl6fvuDk7Ov6Z9vBxUfWvwYdxDW9ombTACWi57ToX
2aAH9g/8oa9CUZK8OkGCNB1oLtUEyE7kQEmbxxB34h1EAjyzXD0Qehz81AeQfOJN
Fcwfv9fOJfpw79f0LSPytluYNhdqEZAPqVv/aAYmTghv7blWTZnIiQF9vRao8jHI
Eii2qXUDJCMuy1y04EgD8zEFFPnUYG09IfshVQRROdFfmNsItqNUR4hvDXZl5VRG
gfcjVYap+c85/4rPoxcBdq/whKfxq5xXLvFDKPYvc0uhX2uZapPQOdfPzHG9T8Y5
jABEuX49WzRucSfZT4WBf+pOrSFTHRgvGj9wVeZ/oG4eES+r7nGOcjRZL92kb+Hz
a5In8trYiLYvdHmHmuwf6lC98ERswpLcNBpdvCW17/lD9tJgQzRSskwiPY2wr/XR
NJ4h/nF7r94AVcVvCxczRs2qm3FoLGXSyB+MGtMQF0KoFmYdaJfqmd2avzOAmdmi
XrnurIccz73efMaRAbYJliUjvCW5O3aRzTYMGfiN94lXjWBg/gF0QU2PrrD4Bdp5
sjGSRbtoxenNbkzdAezheQs74pJmQzMT30+uFbPwr2WflTOZCOl4e9ur0nTaKn/I
qZmoyYeqeeQ0SNRrpUrXhun/LZpN7CYxTsM2FZMMYU8FJm2ivu29Xa3h1gCJ605F
v5rnTQi1fRNJAmFbzaIv54KeCHTHInE3jpmJvVtllRDDxqs/nHootHoR3w+7sPma
3vgviRw/AvrGtOhvhSz817D6uC8oRB7ECGGG5hBnyoPreLxhxdDi8/daHU5X4xeB
DYdzgd/B1iOfZPmyU9XNg76hEN012DelZYxBbD0dCuf7sugNgqc/j+uiz1n/5qis
2aMmzEpfbdtGKa7xxkjENn6cwnf4BZlxvGwhOYsx02U1zZevcWsw7ALQa4pLweBL
Aur/OljArZM/M0fhg2E3ScsXhxjIxh8ny/5Ran1wtKLKuYIQVDRs/ujnY5h2ey3e
cj1WjKY08OedUWYGlbr1fZT6pBY7YIcvkIsPkQvKRMILaZZL1cTRn4Yf1ZalpFNO
BNp1e4rtdgDXqG5lREnCULnIutky/ZZHiijvH4WXaI3cr2vJB0ViFgQ8TwN9UU0c
1+BOPH012ETAWka2UlK+Z75GKxFo+mHpqtPrHTw0C7yq6Pefgu3w+gNOLRxIubZv
9eOv9kSEigGyVFCXzItTiCbhjv3qsPbaO6yt1cVJVQmXVeOHpwu902sUU76p5/nf
zsi/VKr7HL0xjOSzi4aAJWU4Puw/aZbhXGaPUS/Vw+/S8otC/jrASphfq8aCbNdM
0MlEbLIhMi8pBGHHPrAY25R4azJiUKCDgNJ/KEgx0P3Co8yKt3qfN87hlcv8kFIF
nKPpAnpAaWklb8X3QFtIklbku6s49zrIBZXK/CqmtQ4rL57C+ZODYSClRDGY7h15
c1FBaG+lxzMs95qrMxi3gvoaJ53nCCqwRw93NgQylz5AMhQrUpfcmbfeTN0wirNq
bZfH9MO8xQNjVKj2VD0LcLzjEYQytV5O9sDT8BiWKrTm6lCc/a195P8KGlvGhLnT
NzSfc95aZFiCxY1oEHjlWzfuKIyMfX4Kn/3okyL18ZYEESGdXSlOyAOYXxIU5w6c
mrLexeDu0G6jCbqpjwhC/K8H884CUMicy7kZtj2Uq0ncjkvTJ3yd16WCdEoKXEzU
Mp54/DK/ZgMezHBqRV/dVjiDToSzYy/solP7+RLIdA7wNVgXELnb6wFBTAfO96Wl
PbD+sS3dCohinl5qvU+3/G+mqG7+7IcEOtrqYWIuZoOMNzbjXL9mArhIxnjQkhVC
c0V8awX2ZeueoZfdvu6wFlWqs/tXhS+3yeXr0qClap+B44WSt3lUF1LFaZa9DfSM
e4e5fxE0gFTRX62dN4eJQST+VuhhwvyEQ2446hgAqLoJtf6cogONK84FuI8/AHY1
rHIEg0C4xkBC38DXL63lTFZt0/r1Tx8vVV7YaAuCVt1Gwi4rtv1VKMcvREEjkZL1
NrWvPDf2rNTySivshLiTzSFwTdSICQzwMwTvxcKUlHsiJb/MfWxeFnL8p6YaJw2S
moX0WWg7sPaCr8t6uK9c6P05klHi1Tvv/HhiVsHqbOj1MJnnPBcp42GU7DrdSoS+
Ht6AzSZj5fl173E9p8EThWPINZ9rVGPW+3asCxu5DEgZjtOmW8gbRK6ZDQdopCLe
vCQ85BeOEAz4evlb4APreGAvfYg0I8YUk/7Bx//vtfvJKVe4xYJeCaRzxftdfnnT
JQVxUkegHZcXo1M/Zo+847OROG/0uzhRiHovEb5WGkYFcVpLO57jmSuKTKdj/YSQ
Stu5hinQs1fdag4VfQaWzGsb/8pRMKKOt42s8djCk0LwlyAEttj9RH+v6/Jtm+hO
jO2R7th9tfhKPdFy2dp1347rXV5rn56P8lh2R3GsaDdaT///7MVIuXG+gpDS4DKA
ZG0YxZyEKtX8PydgRpsUOPSOBTuciStUg1N9/4zjqnHQebBMi/OfwV4gb3typ+FE
pQ6z2u9RBPPYL4dJfKLkwivn2KJNmMFXPNbEipCHbiUTsbAJ3+8BjWm7d5mhCjCk
kZl19JEDRF4xl4pw7g5kcbqzXSPyDtVjsJS34plC8hK0b+NbtWaouSqPOg9qN7yA
svuTqULtXNMQhqUGQX+l4HWib1uvDdFjSK3mbPRvj+c3fvTllXm1ot4rY/ZdBcEm
BwjIp+OALaDkHGdLOHvZyTNV/PI3xiguX9hRYJsDMFP9SPgjzJpiDpqDrbdRe7eU
x9/UunD2+vlgYxSAknm32JnY0kX/tekBUO1OSHXoYjE9w+bGch9kUPAnFJlcZx28
4HPL2/z3ShgyBluuEYPgEucYrDCIMKrH+AGFh/T2GZERFaqwA/j7Db61Crhwz6IC
zzygbQFZTemLyUPc9r78xPlDGkHpvsx2DGmIeIWPli6OXDADxt+ZtY7gWIzP9fvz
icEQJYcOMsqe3rG8a2kqUDhyJi0fkl8VbIXgoZAzefOdXiyWGo/LdFt3xdDYIT26
yVV58bYgFkLyUpvHlF1bMhXv2KluSFMYFCxUbjc9nv0ZhIHoaffnCjk5WtywwcZ3
Z2hb3Psxvbfh03zq0rre9qo7qZ6hFjCIgsMNoWaGmABRDPR7bEk6QqqQRIaJaU8I
xDqs6zaGsWx0+8xhLk7hOKWqokZ95wl+jssiwS6PaACNHhuU0EXKlzMmRXXKE7j/
Yyg75qMShdZaBxjAyvPBpM0kGYHs4tW5ne/M5A6vjmrhRii2AUU7Kk/uwNqnpn1w
qCetJ/AXEkNS7y3Ni25y0m0RN5mdcdoIF7fxXQbq9mr4uKanAJ7gIYuqJFXzYyVP
OkudOiupN7FgSsvvv3bPMVJqC4ANmVremSJpGFQ3PpXphRnUP177ue10CayGRUsk
rsBrgjYEAxuogcglYq74AxsmoHBZ4i6jsCa2SfUKpCLDHIa0YnC651A3dzVtuzfD
0y9qrmB+eEk86jHpVK21+YcDo8r8hM+yC9tJgbVnsp0Y0K2egEfChF5qTTwfJlqD
ncx7wAZjzdOp+/+WaFsYf2Q9WoM6w5RuglRxpwNBUyGtdc7Dy2DyusFw/mkzxxc0
dd+/NY28SyuZH9UZ2bBDFPT3l6h+TzbJGiIbU5ZErrnUXWPrE2zPk7yu3q5wD7LO
GZEWWknm+ThEI+KCtfBwUp3Td+og7PQQAGnhI1DJ30heuh7hBoDBJYx5bVSQ03tR
0fSpEL/Knwr6J6Y4ZMGmbUrxBKRH6A0oE72Kh++d2Nee18QFvhzi6ByDKK/CdjLQ
/wntP/IH7LFbfJ6krIOb1msltfE9sMkXax65OTxMyVnhcCVoqyQuIgqcHrGsiCmP
FH7ir0/8I+w4Avw+pzgij00I3lm8pBKplKLq2pKj1YhOsAisokbM2Kxc7vW22oLG
MRLFZcSzTV+VkrK7fHil5EkhanunH26AlTH+3S91One4R4QYY1NMkhjYfHM6fp/m
k/VestDt6en9+edJb5GodjVS/QQmGj+HITEsqcVzVJNGQSb9M2w6XKzWsonuXEDR
PmzNXWIAEjV00TmmR/lKha8m0AdMELE8iwHmx0MzgvYl3AVnto4ICmHibqM58lyh
BNQi3XPTP9Sl8fpvP3dIss024wSdBc5c/cvs3gpivtd8J5MIpKRmEmmufsS8z380
hN4PdoWffAyAXaRrLh8+Rqqx3cNISS9T5hzRsFK959GRRbep2/xMmeAkswJM2VlV
NsFf+5sR0HtLq0uYrchvJxrJ/+9YpRIUF+caom8s4+ewsCX2w6mTEY9n9NvzPWru
HUzyXu0GMD9fCxak6qisivLxs8G7hGROXEduTpb59E6hCaFqUn2qbf1Gt0KTc5/f
/A1eOFrlc/9F3siha+dRm/iPsPyfUAEd+CiBwZpMhviZdRq3/Z6h6sjPNXYtIgcQ
7WBHYB/JyGbX4untK/D+iMRpprxc4O9qxOY4I9wAgMpaWbh5ICDmP3CvbqijGuUG
itZoIdmmpvA6hfD3DD0VNIdFhKN1/fQ4ExNe8FvYC2nDFcHPR+fbw74X+G0/BVZE
Vb7I+7bOETnNnqMZTS+mXUTdFLJOX3+vJAQnFdnK0/EeqdUN3Idvzsj9vpyTag0M
OcwSjkUPgnvCtm1PR/nNQLMzaZYLnsw07aZFTfT2O+ypsAG/ot5rYLUYnWvOKInP
N59vB6i79Rpi35Ab9c/zUcdZSF19oUQSadc1AjnmlO+ta6QGlAAhpA1Hc/39au2T
M1SH6z8k9+KsxDmzHuU5dTknvtpwN4yzLgSQs/HfPJ7sLiK4k3gQNPHe8nqgwBtB
aHprG7L8tJS24Y6s6kr0y4hknFR7Sfywe81BPk3PGVp5u2wPTbqi/ifT+BD1G/Lh
/SPFkwDa4GT0GUyPFWOPZBLNBPqNnZ1PtYG6IUwtkXOMzC0bwtYvobVDTp7nao8q
jrdsZ7NMk08+/GmNto27UI13GOZYHPASTN5BiY0HWzGynJwsIegmi0eynXgP0VEs
Wq6PUurjX5wS592znEpWm96RpPs0W81jdbZfuUxNR1Z8DuH55QXMZeoCHoNPlHiI
Dt2EueS/HNKa41/94anjhzC+DGN5px6/BRF6DVXrcKBE1s3A0jTlXVsAkTIrG4tk
nNaVhJ/wDaClwx0zwrz4BlhCtl0HYrhvvmekL5m9APq3RAQySCdSPo3VIfLoObq/
Hh43q8cgg8/2KhgFH2yMzVjZd2gRF1JwGr2nukhHppNCNxwVxk+CEefBV/ftBY8l
tm9QK3i8ltXMQJCeMXcw8OZQ6A6Pg42tssaTV51wjpIYNN9XQJjvuviyiLjuO506
SdDjEQIOREu8D90ZB8TU46D32STwjGyzwuy4JLu7RrbOq6JasCi/5QSLajPK0AgZ
tJdm7yAS1ybyKmsQ8PdvrF/01g/dZpJESoCSjmMgVnPckzU1J2pbDRbjGyPLeIDT
ULJUWstAnpdaNSR4mveuwVITBhtLmzlVdmjk229H+VECCUDganiiH/3zK+B7wV23
gzulebeeo1qSQMe+8Q/Yxy6Wq+WZG8fYoKalTxF+f1KOE8tGxuj5JT2PbFCW04pb
75lKSoWUdOJ54RsPNJi/jz95OGe7r47OnYdpzWsvHIJ2VgqHUXdrNu5LjzHy63zB
Qqfqap8agUXIX3l4KBUVC1iaPZlAx/y7ONHPe2cWl4QkOFs/DFmVqo5DHbaYYW3c
rWvgeCO6onKtRqce6dT+m9pWrUPjs6+V1WM3dXpbWhmo9vfoFnZNhY65weZ5Swqf
/xwhwn1uHDiORuVQnCEfj+jGT6ceIGwPXaJ0cVkM7M7zNd0uVQq39g8Zxv9EBCMP
Y/3wFjTD1n/2l0boJyaGcwMMrzgWcvcCv0kOG7OUJ34IPVWn1EYmFUSCZHWM+gFW
yPKK8v9zVoXyj7SMnv3+mixoMF77BsuWfOFrzzNnOwFqjEt/kEDBtJmqeB0I56Wj
BGaHRpB2DO763OrKmU4CTu8ChfDwX/zECsN7L3o6voOJdLIbmqFaBvH6FRbwTQYP
mvKA5inFX5e6i5fxBj6UvTEOmUZcHGu404+6q63FUd8TnEj5Vt0cqszvahCWTBKm
UuxaqNMEMOtB9Lj6b3s/jH+7TY5IucRM1oVeB2/i3EEMudcyLxZDpJJat9fWrm/L
/wiU0OTchrRVTpIXQNmjzK4wIlb+V5B6LCuHz0Zc++0QPpRagGgk6+Wu3Aw+MzGZ
H4fYQAJLaXxsh4MVJTl7aNbLm52PWmNr3gWN3Zh0oItQ8+wfdP5Go+yoQizMqO9u
UTv8+yrnI8p4UYs1k1WtGi5dU6npGyhy7L9F6gwiaA2QVLmT+lB2i5d3xdkRf57D
tKpKUXRjorDCkAMyRBZkCbkN3+b6KuH5Oyj13lIC3dFWMJgOdFrLNfEDG0AEwZhF
oCcnp9mlmer0sJJHGnjzk/TklUgahYi0RBWqFqBLEnWuEo59pTS21tI9daM9vvph
XJ/p5Wj0XjIeoM//Wk+4ni1pOQRaCs9hm2QWHbmpEA0xuwjPsXoWHl6Re6/cuKG+
zlR81dWNiSvTlpv4m3UECQKoMnNc7tvBTfWCFC2s6/DAXC2TcesgE9L8voyKX16N
Txb8WScIbk0xpEKqZHdNELCZvGZtF+w3kwL2I5gUZmeLpndtA+l4EpuYM3aQa7Vf
Toq6qBJzU8vORYXBhzHFQ+JvQfviI+GRPTVIMSQuB7B/CmMp3fKEJ/RzwCWiZu5+
vVXRJ4TFbEeXBOW5OTSrFx0gAgXUGxiXDpsrDaqIZOywY/SPRBZo33c5ZyaXLoI7
1K2fHlV5bFiqotS2f2ptP+4Z3OTdxRX/+HVisPy3ogwYiAuVcSmyFHBLCHJRSQyM
nsS+yHAyuurBqrd4h10BtvtIPU1cgPrs0GsYtVxMhqXAWB8pNdaiHh/XVbXRhXrO
dR4LbSAn7Q5ExNmCmJSM2lUZRDTJ27i228XnQfISFKuAWH49sIv6Levkt+6hSfHn
uT3NfzFKDeO+dkUNK9pki+abh6umCJmMQmbqaRL+If0e1R9P2v1iQ/ja4CzLQsRw
UdRTFQz6cb1yZNGvcH3ObxWzQYHgMPlkrHs9E5AXeiiAfS3oBFFp7ari5JeTKv87
gN7m5mxJOPukUcYkdUE0kPvfLPU8iUo90WraX5bSMGh0v4dDYxIfVl58udVrk/C7
qsfQhiHV7EoHHWDfrTVhdgcUw5BrwhXWx2jsqPL6e8Wj234OcrRN1oiPbzZZWX+T
LmLImpPBQdZPk03KzpFpLfc0Yb9icCa6En0EEuaoAyE89OqHeNTjgzqgrvWQ/NKp
f0FABuxQ9VXX031jiAYES8nxnaxDHxk5j2P0ZJUVDynvo8PA/skzYUVcWFs2pZV7
Hd/Hw37+/DzPQlCnExm0pLIXC8Q0WT8pACd+WJlKnwZu2MhLTqgCruuLfdRPHcSN
m9So1Vsi/ZW5CuuXQasJGnYsmturbGMKlTlo8cbZFFFNyigzS6A4KQEpS8qGzqmc
7S8iQ6nlj9cqotvwEPuTBgiAuBGMQu43fhWTe7snshwY8ioO5ahv137qSCC/0Ruo
ZJJhKqj/cmbHFOQBcjGu7DgHn2ivhZXHereIWZRQef84C28pBoP+CKBDgdCeZrfS
S4qVbOvYOCitUw6cfq0CL8Gkk20Tog4JZjR/gGWeB0cFRB5LLt7lNhr7zLVgrkB6
f9Bt7mj/Xoivx5pzCgjHFGf9l9F579alrluFo527C7Al1hqDfhppRfCDIi/xezX+
5Og5+VSIPwQWODneUedWE4dZeYJqukHOHSunLQav9DDKir5y/Ee0zV/CEDe0txXA
luZtnePbI8tmrkhTcGpNN+wyG13JJd0NVVogIDxCWzVB6cam17ic6vnuVSFd7AN4
jlKUJ2zFHRqOH36gitlXc2AkH06kRHdYwOcn45W5/s0vwdc2Q0CHqYLBXbcAYHqB
zuHhSQqqSG+4qm/Gx8GOA85EQX/qh1e0ot2MRG8XFNrmOM36Hpy9zOLZM5pVVSdG
VsBr3K5/G8DTYdLzVo+/cylLmuY0cHxuriqlCw4NbVFx0u2xiwgyaxi5ejVNVZUs
0nVyj72aa/uBZn0mYylv7WF67WV9ufptNFC1T+BXiuwaxhPW+AcrhgHopv1s3i5C
FP9TU1W/NwRAKsry9eyKshgUMOpAikKie00m2Ldq2krf+zcdjiLmHow0xdE3lqOY
NF3Qlijp0eMyS8S9ZYZYrPW1Kl7DZLrvv28Y2MuXLhO49jOQsK0d4QEff6x3PxS0
VKvx0gZRuhcDAwaR4rpp9g47BeRH9bs0KlKTlAlg21/+Ct5j9R3+Dox5sKNdRE80
am1L3/+En78oSlY6K5sIeZqUEQahfc8kasYt7r9e2IioI2aR2e05WhOs3zGfjZyO
B3KTcgGalbPceumvy5Ja+ZFYc81Rq9lDsrybYV9F+YniddOWnjsmNYNqgmk3K+Gw
90PTC3REREfaSB0Fx/JA/g+O8iXDeErG9ucE6C0Gk48LcS0e5QImSzJT2GpEIllR
Zme1kZ+A3573muprFWdivFPB8P1ZJ7jWG5SSXoNtsKCRH1I405mzp+LjMbdw27Lt
CkXUjY5sxTpghJrj4tCdTftUtcBdCxZX7JU8C9oyyeljLD1luBSYbPpaW+yEw5w5
Totj0/ltCG1SR+3dGj/GunG61vtiCmTnzaZA36kqoolppNOf7UynaY6nUeJAEIs4
JsX/eCTI+2k5fYDweYQTfVkLBoN3heFbtxYjbE4KlfIO76NNLk0IfWctqzg+5AMB
PEozlHmUwKz6zxufuP/nNeXwELqGOnvq8dbYkEZ/GIdlphU+kvMJ9TzoLiBqC0g/
8lFWEZU2ndWaw9P/74djsBtt3GiKXmK9tN7fSWhzn4vX8t/ietGE6Ac7lq7hGrc6
6ZtuZqUMqcK5EhTMlUPY2ZIFxTxX8Pt/vf9eaSyhgtGXsZDu5P88RqwfQ8szyYvs
e42gNTDVopbQ0r61WQpNwp94JZnzvV8NDLr7/sCs7LskwpV5ubLvsdun/VprvX73
ptM11MUVkXXsXKLJeNXnSWi8KC9qLIAWZ0LE6uQYl+C7wFIhA8P0l9+VTrxgrOEn
xadUgSeNTuE8H7BZJDilF4ZGS0LWPp4Orq62F8QBErDRTN69iwcDNmnt/MqEZ/UZ
g+vHch6zZmqPOADj/o/u7uNZlpGbOYrPlBXvfuPWMjNlJhic9RytrkVuUBOwOXu2
9ANLGk/UJ9euI3ymyo8qLRXTyxmTKYhiCI/dCvBWqluNOUGDI6BMK3mRtIDz2adZ
+3ChQQ8YABr+LOkEsOc87alI/wN6g1fobBZO6cWyMfLYTS3oYSNLe1pWEDXzCH1n
Uamuxk3RU5oU599esDPXnNWl5VEF9UR7SyP0g3pMsHvXkfZN6yDzkk4xHP5llWgD
0QBjaxCZBOU1+1DpVGTxKRH/H8gvpd2RZGDuctYlWthlwugFRDI7rjMiR5b+8iN5
iCqmqlO24LRP/kbxg1V5V1wBtewHmuT0pDBVFMzzC+fq9W5XTxnXlg9f5ZzjJD1J
duFJlzJTQjysMme7gxZQiJ+nkiHGMUKlOMVRilkMaLrvwt8HZCtgHxzEHr6Rgt9N
czJHMjfe88WB1LMK0ZW55dx0vdbC7XyHQJihpUlqjkhOmb2nEcMMO/YcAOoOxlsl
I29Nh3S46Qt4xcC3gwqPIryFVIUbBm8cU9P4r/ULIsPC0bDWLfVbTs58+pFJo8/K
dMle127x42nSAh19ZesYAGjMhCfO/C9Bz3P41UfkpvPNZoHznfPnw/bZN/j7QED9
Q6R5EoQbVuywKh4HKt/OQU3eT2A4wq7RmybjYjIXPao2XhJ+fsJQkwvSzB2aUaCE
G8T5S/6SSkHxuRD8Gd9AHL6GlLia6AhE1l4ts5NClBBnlZ4vkD2flFGls/Xbn++F
aoi84jYeG9gi0luda+6DiSLxmrtHKfflRzY8tSO0ERYVTa6XYpMX7OlpapMKwg3G
202dUmuUL/CdqbD34l6sFYmwheC2kyEQr9MGeOTdzcXnqxpOx8gxDeESodCGDhNN
Fcwu25xJEBD1yQvDUVbQfZm9je/W0opI2j1bakJKy0+nEmbo94DVVAL4n8q35k9Q
WK33hrtr+jlzAgInfHvDkztP1nF8mN9YzbI+q3SfMo0T13k+WxNxbcpBSq8rQTCd
qHZc2C28l8uvtpfgKg0VDVKsGOLJx8YxOtBugkaGjLA6FQEpGRvcMeCrL9r/GGkc
rI7h9A6UpzAG+B3nef1AChxcBd3m+mXKtf47lAs1eJuVT0/Grsrtk9Yl2VIjpbFA
ddCbpvRreHKbk7bhQfeLUbsupgFJUWi3YzU8pjNdSAGNmhCefxRfvqfIZA5TJKq9
YPE+2D38M4otQixGJ4xf+Kc87BIaLW9CBXQqgK0wQrYa+tKLq9awyRGoHkysPvTv
JRnftk9ZYNJAbFzXgD/1+C4DnVfAA8r3i6yOniwD/EgKZlBIKf1Hif3M2oHSPwXf
ebq1wnDZRUChWr3UZAFBpBT7GxBIObi1mmHD3ENubpvPivIVn+MAiM5cbjBgviOv
A0G4FKbNtw1TcYHZdWLb8olJhNNjX9R8GzwPyn33JabAd1BCZADwDB9Pmxh0tDwy
Jx2ZTV1oxog5RY13vCFcPiOcxVnL1ieXNbklBuzX+7A30X0swzYIZP89xaMa1Kq4
lcz+TUJl9fOvH4VcXRWP4gT8THHhvDYpAHW15icybDLaeSholtjwrrRKhQ60qn3X
1xAdw1gm6vQHf66Srw7JFQRMN+ALc1uZ/R8t8Ro4sGHlWiyYsJR/qToglnyDQPii
dt35eimy0qG9VyGlzCj/vXDFyDacZzO9hY1G+8wcS8p8xnGlduC1oKNpJQ5KNAuF
hqwGEAYBrPcIHWOyXtj+DMah72Cw3GTFryVWQ2M7sHv4whlOAtMeUpzJ6NryRumf
VCaolHuJJZqxBTYw4dWBZWWaI3BJmAlRpocpqorRObuURqfvIlv4a6wbWriMUpc2
UCydL0yeSvJkOEVU8bi4GtEa9iSsa+FaaY7TcDgLbR583uUU1q2wMrLrWmEV9cRy
0nSTpoja4Oul1QISSP+IQaVl5iTQQ3HvYtOBNKPyEgrMqU16HMB8hS/DDPMgG1Jx
ecr4jnkqpNHSuMiP4wnXse1ppx19/XPVl7YrCwt7kLLC4wokj/Miqri3HIgub8Sw
zhW43rNg698mB54qPt062H+Q7jAu10uwW0JFxtELJeCB6bMZVhCwl68wW4zeBTx7
wIPr42iQPBOsGu66Y0EFCHvFF4ujpxH2xlkzryU+VV3V5KosECpMuCgj+hf4lWxC
KNW4WyJQugoatxYoz2TnSw5TVuh71Zy2EXGGxC+Urx9LjCtOE726413ZhAWXeI5E
shH3esR75onV/Jm7JUsa/ETKqUg/WlDYkis0V61Dnf01aaXmQaKn/5BuBkr3EIrA
9l2AADPvslo158HnGolDzz4LASIiEF+UO8dxtWx2py1OXEyFrj9deOEzExDCSKaZ
41cuaOpbrX61I92SrVTHxx/t1OUoNWrHgZZucLJi3nz5+wOuk6j+l/1vQAJwJAoA
cKDLnTOP6eZVeptRFSrjyio3V3IxYPjCoVB50veL7K7OqvCY27KVh6pXIIroN/cj
vi/R4mLupeQ2SiACTUF3c2Qb+AG6Nu8oXs4/xz6KU6C955FkeeEyRa2vPZaJZ7wo
JL5LFsK9I/eTp25ChXjj2wwEfvsHIrIufI9ZYOrLk3seQ9OwtXxDBa4lm1MwU+hc
29r05LQD4mBoGQl2v+krR2AUbA+C+RoDoCA9HIgh7e/iS54MtM9NQ+BJ6wd+F47i
5Z7/0R0zZw1I+Df9ZZniTSjOVmUzH+aRAKDG6ca2eIqR7EfUcmDeCpIVhrn7hr40
rlv0188uPQTB5U6O7bJKEwZ0iLh9KUpoojjRVDeIvzs2wCVP6R7FJT76nyf8Dil2
U1VYDh+AG4D6yQDyKxT/GeJNUZcla4xcdbaWjB3I7MFNpiRI7gKrNAtGkspt5Woh
ARSyY/Hd4hzjoPGqb15Kexq1vu3KzCA9vYCSVH8MMsZMYKD42zimeUohMSgKB/59
nswDc17TLEaNH6ikZotyQi0rRFPLZ9pVlvbJxMtedzESNO9wVsVeRASsi3wG0io2
ELOufcYnb7+nORY+wFa0n8xCHklZdgDepFQf8YZQZQmGnMl0IBk224MhiDouSNQU
dZnDH/Dm9MGftIvYiUSVHfZP9Dhp1OEl07c068Gm0DpIC0AqdIzGpfnDDeBScxJ0
ttopA1KN8/BQEDQEybQtiinYFvyqZorNqIQCeGxwYZqno90snLB63h5/5CvoCmBx
ucC1n74jBuoOLLtotki3zVYn1xS86rBeVQVRTQt5yH0NNHRL8El5D8QeGgZ8mAck
TiI36nvyKZq9MlNn/mOwxAKqYQhSHGcmu4yq95s00NNL1bI+7U+ePu8jMEZ72FzI
CbflzgoCMqA591jrauRVKORoAHSHs5PdRabD4ZDOH4j/aD5ejyTRkkDoIRyE8WJa
uTcXIKj7rsF7OtBCGZJakf5CGgno2+XH81dXvS/v2+qzH+UEH4VEwz/rBx/na9Vp
Xzvy5Ks4oYP5+Mj+TmjWdSLFfJNobUB56zADAbhW812TipW+pxLlkuFumlbHD5WZ
E0xgahGOAzD4LTY+h+u3SWvpWPRedImAog71UbgLBeGu7Zh9zW800iXQeU7kJs2n
A0/RUsruzWispD5KyKOY9SOG7YiB/nf+5AOZI81z1KYsSDK2FOaxaMh9sDdqsjb8
gi4MKYGJVbOx7XcsEKVH9qS1cTFoX7fsZAqt2DY1u1TSd730htNUHeOAdtehs2T6
+9d4dWr+c7REqiYhMWa4Wlw6UWwsahDF76iB1P1TZadFVBkJzoQZk+NQ9BtTohL9
uSOgrHemGwm+8zvoVkI3U6DUZWXv1QrXCkQFGQH4TSxPRVrWqhf/lUoDMlTFscMq
AcnreFUntk6FarZ6OGIpBJHlhi6XTNDkYLg96X3bghZRCulfr9lvwLqPOU95XeUH
YkeQiClvQw5ZnK/ASggdw31zyGpLjAFzNEzqsv1oTz4pQiE7G9L9b2oIInRwO6tw
/6tf64rsTN0voR4A68PjotcDkQ0kvP/QoZCGbAOtFzjx0EusnoG6bU+suxGTTHhs
lBlPLIcHfaYQndhjqPx/lCyGtNCaQhgbcktMocs4Zr5hxFq0ERMDEgqtcCC0ZSwr
r6UCB0+XjKrobVUsNdcdkFqa0VUXpt9VhQItFIbrwp5UnYQj2cih8nn8e4pgRBmz
5oaBig3iRr76wnv0tiITPmsSnovja0bZBAQKgNAPtQjPmAEYAHOShVl4VTXtL93W
I1jtwzkv8Aa3TlxYcDO6hBdos0F9NxXNGqP8q3ZWz8XXxEdRf02W1d9nfaU2EdAH
8+Ib7gmlIU0owppIm0r7XrGVeaj37JX1hXE4IMvfvGHDgMBGLK3MLvHjcGoekt8Q
3ims3tC+QBaEX/rIN9vrYu9Qj2P0wt8UJh8TM5Ue0DLD2fs894coPr8YE9UJgH5O
E+0ZU6HSkPU2HRVPnRW7pQIz83iGt2H8weN7WB+3i/O5HUiRYw2UHTx0+RVY4Ra+
2QoRYRaNAldyMju4kojDQt88U7ud6QjU4mcRxVojAykX/G11TxVRnokQeF5G+LSz
VsyjHm2e90BdpUB9IyZpln72BuFHdVYaoHfzAgZf4ZrNSDntVBxtyRHidcOQ7ohI
CzLkZzSkJle7mt8+8YgNJjRNoOWx6xAe1Z5dvIRICQIX/vq5M2mHohMq2y9SCiQI
yNTJYlp3R+UhNQR/VfT3Ee2S5YkDpTVb+F7RWtIFJzZnRzHYgf4AIqs0wp1armay
dRhubWASBGNhYha+1LPm/LeKegFPW+Lgu4cALAJWs3mpJGcOdRTg2CSh4I0BlNtl
LalkAhFUdmOngjXWfPaKFU+6ATr+xgGKtcLIS7ZM9K+wK7vfFwBOR5GN+Oc5mlKt
ovyRt6UbLdIee5xbzzNCZWjnbFBLseogJ3cOnK8PrWpT0xfibT7IczIrgdIyW4mh
+GPZrdjPk28VKv3mH+hTG07EuhlxolsXFsAoQ3QvyOr7Rn7sLjIOhCTCoB5uqoTX
SsR20wfA5ot93+wy23WoBl2FuMnYSTiNKxPejgxKAWhpa4WAdjl1cvEE5ozqm3bS
nmTLSLbxfutM9DfHW+oM7H6GsBqI2fq3cSKMKfD6YLPWtcw3LRI+3h1Z4O3A+oBl
5kyKKxITaQ3jQEhhssc3J2vkpXJXN5R/uL3VaEzp2rvnysMCH0zp+4JcZL91SSnx
UeuWnLW/E0E1wX5G472p6TMgRzKDLgFbToryNjlQxKIjUfKmJWGkCCqmxwLGXeI3
r3bvf76OtYyZL8d+EDHJ5eEIgikZddLbQqvpqcjVDaqvA0CNmItd1YTOoWEOd8j7
/YAK+BwZ97Q6cgAslNFzYYlM2BlGZWBy4RBJ40Peptf4WtH6ZboM5rtQBEQMiaeV
MvD9ZASEN6/9/VlvkZGw2x7yf+/S3QHiOtYkMJoLVqRW8SXR9j/qZhZPd+z2HROH
42/iwfUZAgzN9LhfR2kGp+YAd/lr5TniGTU25yVt7Fd1uYQx+rrNZ+ub71Lqfqi/
0gMnbm+rWi/7mpuhue4yThOCZsGDXfNICrL7IvOQZYgvpQUxZRfAlL45SIHsNsKz
P8yzXvK3FQx3lbBpXB8saex1lfLfUs6823SusH4EuN+TMYqIeGlpxAyqbi3tWUun
OrsCHVAwhvl29yrNsEX4wb897TbRfWdzNrjvUWjBKJ/E4m4qkbstUVfOq9ThjCgZ
kbTTMBQD3jsspa8oUDIvnPZDScyk6qt3YjEkjqZW3U1BdFmPixxtburRJB6q9DGq
bemsMwakLhmlClo11ctb8/sbUJS4vs6O9SGNbk/WdIeqX4kLmoucsoj64L25sUKX
DsHR+WZKUBMPfrDV1csyzJiuZhX0p3x9mQkvTaVOlEvnLgyhhlUGb0jYLvayjZbn
sVrDUkHD+CvpMy6Tr9gTiFPkZkFH/iw41XhY1RvZLsOYP2kGQIL7fFk5pecmtKSL
az8Zhbq87h0z7tkBpeOEUC3/NeM/KOhy+q3gAzrr43za/k/OuY4JBywpY5Vx9SeR
7KAoGJYFI81eZP0XbuLTG69dfW58uVLImcrTFWhkdhfiQWxYAgplrueixRIFFD2r
mQY2ICrmSKaSk12bkXYsYHgxQv2wLpsy18pOpD8ufGAWBDcPm0tljNZaPNyewRsZ
S/zr2PlxEOhl3VcVTLVrLvx/N83Q23cOIc/AyTLR6ET9E7J+Pz7SMqEAomhM/jW4
UB84K7CL6UXpbTVA5/NVs9f1FVaTPVp6o0mdhyWy1N/rnBo8luJ3VpQrJZaPe8It
VMVnEE1N99odVyNQQL+TFkw+CG4T2M5LGkSwnHfP0/1102XnZ5W5fbRYH3TZrfEx
z+p841LoO+LIiSif8XRR3p6RoHiGcccYI+1UWYBnMw5HlN0IHWcFmZ/V5xo8YC0I
mYA7rervuF9dsu5J2Ios7A8OUvS4sqD2Phg9zR4AB06wkTorT0b83ABi353U8g/L
jg27icmOX191am71gIk51Lziu8CpybTdkySpYhwU3GrBNLWQePhxapOhm1AFnXB7
2oQz1iPD5X5aZx7PaUxf7+8mXdIyjkE9SpXBoyAgLiCK7F7SfY9a5WelZFvZFUj1
bUZPQDqFJjHrk8KoAQft5JIcftqMS6wdL+Ddagw8hYGs40V46No1nHNJdsKOo610
Q7UMYOt5ioADr9xV2lF6OZfYcnNzLt1ZAmt/6aRERTeq8LLv55vt8JFU/PHvPoN9
eeZS0OY1iYdffsA6kig4AfxhDBjNUmSxwWxAtw5OiECTwewkBWXmXgkZLFVmWyE/
1AJiHoohJPjkxZF/L9sCXfehGm23BQUmWfMFu9L4HhxmU/NUj+W2PhppS/DO6Skv
OlPpij3sr7hp7M0btpfxA3KA/IuqzHGH2UO1kA6DW9mOrLuGAvDbUEN9KSzizVVk
UC/TDkJMq3da0WQHOCcR5fnT2mKOfRn7RMU+3Cu82rvNAp8AnMHiyq5Woh8rzvt3
+aHhuxwQCEaEj0jNpPViqfZ5L6NbiZqtMkA2s8OWqw6/TOFs2l3WmuocvO7cmNKF
dxSWieBgeaclPxsnN0BGciTIGvuHKeJztmEM99RmKYxpkFe1LjDMe8PNWVr7QVrF
DKepXZGIz1g0Y4RiHo7vbnI6TNBVHkFWB3zTsHINe8t0HGRiSG406h7au+0qQpvs
D5ItipJH30gdmIUOIWdZB/HWnxxr4j+Cr8ihUM1ExTuPpLn3TvfrlHEI9AEaOYK5
ReXSYRbOuTAAwE1cshRqGKfLLOkGnptyPLJVyNd2XPFEnJV6qg7a52LLP1C4b/UI
FE34x5FfW1FJ5O9oknI0rxTMyDgT4v+FkDJ1KLETXXU4z7/XQuWD5irdVq/sEbzD
7mPpd/c7DzQs1flNXY/P6FGzRK4cByyJH6CU+biIHikl9GsZIEVwgMTAlHK9uZ0q
ylXZA+2We/gzULkFvNbsmKnVJb52D8W7320bd1lrjRIyyYm4uf7G3ZuFMe/0/N2n
t6XAGwzi64bqrWAoeNPc19Td1IMZuicK3k29w2NZfY4+rCqPNW+Y+JXEQjIxdvGW
isgTRg6p/sfI7s7ztQqJCyqTY2v3RMzirMFXaCn8t2NbPaoThSj+6xwRmq03c/+O
bruSA+q5tc2lHj/Zq3L+IkBS+Bhsb5mbPuVaUtxhh7tsPEcU5wh61Olp6NmpcThN
tJzTHrsOMwDOrDGfMdAtsrA4bbTNcezR+dMtryDeqw4e+DSufDlo8VqJhF2+yNxh
MKIrSU4ZyvYOc8bPIEzJhji9gO2zJugHLDHHWYz7q+qC3lUouncRTObo+lV7u472
lOYHnZBQuLXyz0YQOx91ElRZNqBRuQHwxDKFiyZOpGSBHQ2qVeqPVUDfPvjXn2pd
aiXh1fgyzTSdjjX+ntx6Epx8IFosM9nE+OiOqeHTii7okW5neWEMwoHfvYoTdEiW
8/0jJQ8Bk4ZnAo9pfGjF7+2vVSm1XCpZqwoZ+NE5Tpmf6PpE053LMF5vg6Cywd1p
WsEt50pmzCmPAqtNczzeo2EaIMrfmLTkWS96DKlpR0ZHHXiLUG8ot/OP9fq2HZmH
GGtobmfQrIBgksf/KYkEhKm90wvhmvmz/swchMNgflIeGSiaOAcHYE8FXyNd4e89
LQqrdz2chji3FcKqWIb8d8uq6td9vyknFX/JRHg6tNwDSy++ZSAxWd5SKPHoej2L
iSjc4RE8FYlsBCa/xoeJDs2L9+KmkO8p9HXwGoEFkcB6LJjmDC+tIqJfHwwWpFp7
MBlqCPDIQtcUKETa4tiyivpUG4iElgrzosGQcx1RNvGk80msNkxXfDhSJ0F92UqJ
+WWc2nOsS+h8dalo6beLJRDvfSGS8F5R9SP59BjR0Wez/eAxB3ix5Dw8pN/dpud7
YB6FWw8V60Dru7W3oRqZgo8iDfgoMkfp/eux9frYoFbq1Dz6qRn418xdgcYAc2+K
HBWTclWN06r1EDj6LUERSaSvJcH3n4mqlBAZqb/FnBzLoqzskk6Xy2iUPM3sk8Cu
6BqrEBhYXWTka0LPX2iczLNVkU9pVXDKOCZ9YM2rBCpeAQloy/XJvSq4tacuDK5Y
5DWH2kTWqsu2TOYwZZvE2r4b1OU6KhoHS0367zrXwP+RS3B0PJap6Z/NKsGtYABY
8FKfKFGIZufA6rqXgm8bBqTEAoyeLhZ+lt2hIqMrdVCajeoAtAVqFWyjRAcDLeOw
VgLvyRo/Rq/u9L6mh6q3h+YgHy+syB4m1C2xvQMqApQXe7/xoeflp5AIjpv9CC/T
mNuNf+6DyjjzabPNr7uQ+FPOkCVb453/Lhe/+RcJD9NRCfqahQsLGz9uvMeTGxgK
9JT94Onuc4Wgsr+UqzgvsStVvOJq6BewYx+84rxFP9uRDwov7Njd+j/8RjM4+HYv
43LYizMK1Kjg8TVo4V4BnV7jCCMdrWioICY9v7DAtVKdTck0RhWAoSC4FNfbQSKN
n+GXX4VwX7daMzYm7Ac6zq75tg6u5g/oQpTTEeGYX0qTc0Rw52llCm1CkBY+XHK3
BO+8cqtZ4S+Lgpw9Z1QoGlIoDo1Y7Pjmj+4GOw7OIRHpcEPwW4FRMDRjR+WrkRdi
/+sDB+PIYyYVzBtUL4RR9iUeZjXIMjhTJJfD8PYNV8Nrfxq0B9IeaKWRmaJ/2GaD
rv2ig/0Unm7Nmxi4O03Kmo8sEMlVBWZrkR0uv0d+BW66GlhTxyHgLB4aF2xD2iv3
84XR705gmGc88s5aE3CgcYyhhczPrv/meXj6ZyI31u5lKpPslTfnI4RMVg2ZRgVg
Xh1kKJ+98VUgKqDS5MPisLjweTU0pflDhHtvDiJKtyNnvcRfDQa0+ekfuVKeZCzD
Z9RtvGeueh4a2hOIspcNlWqlkfnRop7REcktrFE9zfrN3F8QnXHP51qVWtj9++9C
cshLTW49Zz0n7zRj4ap5P+3Cbj7HAh9o498Va0GyjmOpzIWudkHBhJgc1dbVAHsp
uKGG79UlO68HsxGahJUHq0SUF41DyzGgEv4n6YVR1FX2zJ/Qasx4hRbfsRSdzAx4
NfBxeBP13TDXiTKwxkDo0eKlbgvoqkp0iNbEijjYaRsXs76sgGAn4gB+RDDLGfJ0
2kgzsGtavq5JuUWmbT0Ps1fzAaBUJl6aWdQj1GOcn+ygfjqXziWEduS/jT1F602A
A/bEWuz/iVax5HhpVt84h4AJCPO5QGTLhIZSMc745Mfg71T1yZydCLRX/g3NOgrE
LneiLWu5OK3pvCMNnY+hQeFEpuiVpdLg6K0oKFUflST3hdyHCdhKf4gzpHzM9kEx
BltOHckiQg01E0HwcVh2oJY477Sjg1GavZgz3JvIFS4t7LAkm1j1dqflrOcLDURk
4lMtuTH/TPMpDJ6RKfDsEXdf2qPQv3ALyC6BpX3E1X7QGod33Q0sUFAIiKTb4yat
cFm2dYovoOrmmInfRDKw7E5gVTrs1Wqo483dPCWZ00XRsJLYHRWi4Vf1wZyqVcIx
iz+zcSPbGjtaZqjacLilMkzeL0QQL4maR9WkIx8KqU7rQGjOrIUTFG6FbcZi/mL8
FX4Qy1Zs6sVB0WehONhj+86RzHvSMTnuMsnjInOyVYXy0DWtJaPy9raIxLqD3b4X
GlrMmcnJ9JzDwMlO6elBsX4KsplwK9Td95ZWBUzPT0Yh5pQugeMJ3xqHSkNJRCat
rslaExWv4/+UTv6wHgaO+wBT5sIkq6+XJ9+RYch1mo1ksa46Avc2voTn2K1r9e4l
ZpXi80kwJheOTiiX10+FLfR0wOjG1Pf8B8J4TWZPcSashojUtytsvFcUfy7ikgyg
1//tc8am7QQbKXAxbR61uoCCCl4I2hpHg3waRot8b4WwowWF+pkFgfDTKUEVUuw9
DIEu+bg7oYrN4JflbtoXHqoyWPVzxRrIHZLUmY2ZsyCzXDkwbqVI0blFf1Qlw8TR
0DRKQLlB24l5uZq5bVySxhRg320JqgMB6kZeIjvSxUJh3TSJI5V9DJu64FMudxN9
XmkZrFkQ3l5kLuHPUeIsD69GpEvTkHJa0uhYKHlZtyt/keIXkTBtUUZZYnw7cTrD
lKn1sjP0sDzCUJ5MqFW+/fEcTT8S9fuHu5+8i3zz3SNZO+SSAtf7VujKKqOxO3VP
3yTomt6RsG2SrEpspTy4duEeUNuRfn03QnZK0xexhR5YkuSvi6rjMd1e22d+QPMh
3tJ00dsBOtA8dGKsAlvzAVFYk+7BiXlsjy1yQZgtzWPKUth9LcvRQBl45s4jQm7U
heZ6GGKcfCg+oxOurKIhcuzoLKvADGQNup1ZYXoQd9b2Oq2IzsnAWY8pkb1qrlK/
irT2c5AzrtWbCOx1SQ15x2O8r8dI4Duq3QSzKqcrD1ok9D4F5h+nxWNCO4PAy7ks
VhAu8OQz7FOwbwycJAUZnV+m2ZicI91mg22sdeqQPIDJ3b2+F51HYqMAkLNBmwPz
OnUy2ehmPMVMM22fMMLsNoJN77MB2baRkp0ubpcpe0JS4eDh5HfRrYo+XoSpWXYJ
QoPPRgD/ZJ0fVVRNImFxlCHXUHP6NyU0+p5hvpcACxLXRVn5O3dnZ3MR/cs2oaII
yEi1vsf4dzX+0M3OIaeGfqUBv6G8fsWfzAStuYr6TPaq3XJLgTx1FWrWELWw3wEA
RjWfzncw/1TNkA7p2yTC57H1QteARIv309GM7xOt/DfZJSQIejPzEl8vgqn03aN0
iP7V1Y1UFds70V6vUEj8IiMDwf7yyZpXsckONNCw4KyDJB2wZxDkCf+wIuEZn3Hi
LGBVn1wmy3PGZw3ayv3e8/T69AvAw73itM7SsLjmDFHhBXEM/e66IEOAi5IpWoDn
CgrpDlucsoyWIScEI21yfpuyO+kj17JlxfsfiMnsiCgh7iVMPH7fTTEQ0DdfOUJT
ONyAwTFRO1KzeklbSBeS2MSQHGhw9V+/WPhFbuc9+loE9WaTzlLeLTv17Ca+/0j3
3neHu2rPlZ+ECiLdUsSmKNqnbblD44Cs406qdH1oXHAMRHzLCxCkFmn+EXxgNfCi
B/no6+3AfnVO6kVfKL9wEbj2Tf40t1z1NpZ2o1fid1ba/ESoyQ2GglC7DeFs8HiW
VraZNWF4WUqs/N5QewV1PVCj4VdHS9qbW9bagjG0nTgwYxHNi7anG1ZXQwgiAUda
/ALWKoPlZoNzq5X8qiNk7iqhp+gc0hP/RoTvn9fWghpwWbLSw/hntOUs/MK0+9KB
LSqh3kSb+ifGgutr0w5KE19rOZa9GyChNoHLvc2sElSrOCbfwVyF59003+u5UL5B
Qub16lOKSbvz0yHtRa4WfOdFq4tTb7RuBJlUFwmnGkV26gquJmn+15fa7G9TSUiH
gIejk95Kn7XGivFMwYbwXVNv2h4dnRMqh3XBBnu6qNUHu+Apz4Ou6ofEQ5kO/J5a
Z1Xh+ntSAxQ3QgwDoh82I/sQNK1kxUjCr+nWcHz+P6kKUrQfwzbsSxX1w74SfcKl
1n0Z1ucY/eW+cbg4daWewX5vzbg0sF/JiDwM/8mK07WryeECYu++MNCPqJU7NzlN
Epf7uDnAdrxUcrwHpgaOyXn+3fPTSEcuMNnXGnyXLb//D/BtLT9s0/3B/kK3dTTI
n2ec6uA1dJwBAxG5ZindvhFhGFezp3ayTtKgdzkG5udGUZ+wKSZ5BhiAxubN9Q9M
+JWa6B4q2lRItdqqxsB8UTVWcu1rRP+ASPvIpZUPwUXRZp3nyHHrWYDTdwSajUmU
HQVxVhuTtHulJ2VNaeRhWjrRa0r70yKwzcmFOKnoYpiXe8LK7o63N2U49nA1G0f4
zp19S9p9q9ZO6fiH0truVSO30rfuvwfN19fpRW2yOHSF21bkcM44HwAkQ3ChKCss
psTKWEEhDamkoSdwDF6JbDu3LOYSO0joC68T6s8efKlsYYLzJcmLKNgE70EXzZcR
2sb9r//ovmEby7xIvGxIiKIGrq+URaKvtlxHtIlB1GXL7d9hReWDGv4Tfw2dBvuQ
tGUPmsu8Unhcw92a9T6sUmMHRMKkihqyVZc7VEw1mUJOj0Crr5wiByVmL/DBWra8
ZiDRq7Q0DwxWeT2Til8uAqdjsz/r5xkzR9K6TOz0dK1TtQL4wu/O6t8LvtV7bOWb
t5Qns/ofF8xr2kaRYA8R+BebPPbkpvIEcKg1sUcovHSqHr+k5W8SDDPS6Wm7FaDd
oMAWP28mSDxd60wu4THmV4BF8Wu3er1H7qCuN9Q62OwAknJCNM9shZS80DG45DRP
rkVpcTx4/CxvZLifsBND9LeufCXR6bRoskSnAKgN+SIoV1FRXKEWAkLpzDWpuesv
5Cl3ujJRGuHba+/P4LbcvCg9T1e8nwhbgXcj1AJDIPyu6KqO3wn85YZDAOmautnT
Gs6Feg9bu5ZhZCiiECv+MvksHCzdkxFhrbgw7E2FbwAb8UrhPVGC8KFC+CCigyhZ
8RsSiLm1wuzvhJluS8CDiBDgXCTc6rGX42NdBzdF9pPs56VyBvksxh2m0n7pOiRe
ZlY2lxGi8266W1ZohmBxHSZ/BeVicE9nxp7SlD5aDTF6yhx6sI2MI6WmESEfZ1GS
U0OmfY1tyJgCXZkoE/Bb+ZwRVtdAXU4+zfbijy4C4twSVNl7QHanvhbE6T7OEuhL
i5nuBSeWaqPyLjAV2XtogCgTz+8PTX4ogPRhMTUOucMST1JHKq7cFrm8uG62zAs9
ueZ+v35H0x+YpGuDp1MkxcALv+mBhMdW69QGg8dIR+Alq930oQKEem56+eZJIkSS
AKy/WhsqxUT3nsKivXOIyeJEbc3KVBjgEEyPVjoaDqsn8dI1355YdJN3b+7P4iza
lbVhZ1qA1PnLVFbWGTDtHET4+yg519Uwu+dOKh4ilP3D9B57y7hqtofGKDAM7WMU
dKTaAAkC2uijlrjvEQN7Ialp68XjTO0g2K2JDiwMZhvypXe2HKtqCQkSDZUHy0iV
tSfKWKChDrRtByVeDJ5PsdNOEwCiHAYyF5oL30y65YbhF9xJGrKC1OkCvheBOpgB
omQDGucWQXjzGYJj7CPV9S9wl6DrIaLNSQBKXcwwzyUaXGlrV4wMJ/uY/LDlSYL1
I6ggaub5Nb4ztaU9HacJKzbnWm6I3QmtYlz1wv3KicQvC6EmrEuYLIrgu6DCS63h
qh7Xt53odVC18OM0rJs0/QlX+HxFqgaytSv109+z/prFkkMJaj4LCZx8WQlV5HmX
1ZN/2XFINan+h4pl7TLRdejUcppnPVuANqtTZH1Q5BNTRS4C0WmIYbEaZh4RUrU8
deZLbuzpNwj7zamVsWcGUnM9CL6kLKc7mQwCR+UMBuPPEM9C6zUd5BtaCp0C+Lv1
Ve2+AFwltb8D+StMP7gCMwvXi9cLS+h7Cp0x0xa4B6BVOisiie0Mo6vHwsxokDd7
g6SCPKG/3VgRS+gDh3SY82GVNcgp/kZPnthQVySqM9bwgc9eu8K4c+ey9Uejpjtp
Sfho64mizYDDY4MM97UjLLGF01zFqZaohQNxfP5Ktose/yBg8RvTVBRTMg+2BKWv
du8RH5nZrgbh2/X6mVcigPc1bncI6W8a3vK1xlUKnZtuJ+qJ2lFR0VuZGIMu1xXq
MvwJB0hFMwSobuuTidugi8quZSaktH4g7e5SpwD40lsJPmhdOSjRro/KkCFDPi7V
TffEX0mlJ4fMHi+0F7pTUkzNET9cAH+1em+yBHCECPTTnxaRXr4NAdXvTrQu5mNr
NqSJE5lvT6PgITyGWgmEGOg5B/4sXj2DiZtS+YulOhUAK2/VyB8nVs1O5a+d4AjM
sMKGAdauaWNERksEeTYw76HLOmenU42Ex2gjlYSD+geA7A2qskCmTN4JloWBUccJ
Cfrxc0L/DvHvMx/Gp0dO9vE1mvPK1Jm4Kl6P61WCQ4FqjaN2+3Fr6JVUaQf+3JWw
Ok9h9pNqttOGlH/2MeFooeL0wsHwKfIHZr2anpnQcLwHZQX5NnEpWzTplJu5hANq
cXIKHo0CE7nNG7FCMgPDXl9GYgjFHGrVdUm7COI3BdtiGZk9I35eUVwixCm2vXQ/
jmwvsDx0l0pGt1PYmixLATo+olflhKaFRqyNClgSn+g0mhG89EUWU7Fvepj9ORY8
PejGw+YPnkQGBpOhbGTxvWa9rKiETQe/E7f/XMT15wkX3Il3RJ3ZOj4jIcvsJ9II
LM7tWN1pTjYCoFrmkGzryCmxjX85A5gD/PUQrAF6Y/Q12zfSUcdmZpMOnXH5fg9r
96//vO7tEbJ6H7oMg5xqLQ//ACW4jKlZyPeIBf6luCbVVyTMWP26hQ20W6mu8oc5
DZeVuho27Bee89SvCdNdb4z9ZMmoGLbJSELVRSz1ZxZ7SttSpzmVAeXGXcnCEsnG
BkzTFpOegFAUb2RP3f4mzguO251gDDyo/Ym2F7SahxKCvtT3fU9dY50i8SkpAX2F
SRx5Ajfd4ytcwPGjp1HtrMDFgGtH/Dtw6852yNbjaSaM/tbxjOLqY1qd1DfekzCW
5WmBKqvF7Fb+IPi4KYhM49XIv3EE3qNOG4fqxvy/mpvELkZKqLwzB7HSX5JXQwDa
3sGhed4LQPx37SQBgHrGRsHVaU86ojeXeKqJktpljfNJ+Radcbw1XQJeMg41SLcw
/v+7Liz9BchCyi4FNw1CCTw6szgbzdFh/CGb9wvX/fOmdikepp/rvrxbwTkh8y3g
XRs+rHCvW29bDwISJAnuI00qbm3D+kMvnrkB27xlmh/ykR3Q6I1WjNd9dJoYWBW/
NTdsLV/PLVA2OSZPUt7rml3XkZN1wa6kKnaP4m+K3lcdaFbl8S05oWahq9vnDJxK
sizFbhcn5zT55q78e93IOEYRs62W5pVGeIOk22dXSI0Lmt/moQJjz1aMDVGNH8VS
ND6gWUt5bWBC3CmwZAR3EE5MgbHKlIeKZoCqkQydbOEowsqrMixar5UPZ3ETL6m7
jEkPeGP17+eIIZV0Ggf36N71pKxrGp02O5zoyQei/j+by4JBFwx5/L5yTMMNc3XV
nB4xL6FIPF85QQlShELOtz7fa/cx7Njj3iKJlPgL/3zsWQ7owqTzvCtWTp3UIrKu
yaWYVtNX+b/Vc1GTIdx8rtLs2ZNCSclx7b4cmjPa+twwMeVGPtrO8t0/xiCQe6DY
q38qORo6QLWtwwALwBLnanxqKDqRXqDRSmuEABmCx2pThusTsRdB+taitu0BuoJk
wQ4cBhQxKHCiAOKfyrfYbnhJyVMixwzhJNQq3nmYBuzWcY9ZT9QBChswRcX3PAfs
IAhrfJ0RKjzvIT7QDEV3Ajj5i5Eul1wXyQ8L4YMy4QjoitczbzAhkQsA4LQCk/Oh
eVevO1caAiLv/pnDXdjequgYvfQZQ1QjMOd33ri48Cw3nfcmzJuu0EOOEuBfL02I
fXTlY+lOii1yp98kXrMU9pVXSW9J6TnRxYbuFrh4SOyhx4GpAb33zDnD9/Rof9sN
ER/sOUdiN8uvmZIP0F1U6IMRXdK8Loj/i/JYcN6hOcr6L5qg2Bcr3LgMTSQAFuk6
7JnfiXw5mGt9Jld3xwUHxcTCtIgyolwDSyvIuyHzWNz9idoJYcludAbcyQxvr5IF
BHhnlEFD7bYgKXvjnklbfq1QxiUjqCrp8EKsiwgF/9z8gsXbK0Q84s8s7UID5DVG
GjAWfyp2pJbRIvPNRLgahozLXpYjhjI+9ToUrTJeKixQGxPa14RKtw1uAqMEeF59
AzRIShZMXOSBuwbdeU8m9cPEwjsnfb3C5k5V200vbU/SBgWNbL4FyyAOYicbzfk5
WPVb9l1TT158rMEmMt5I+u/43jFOiox5xVRuKQY01NmZwqxRBeKg9TeuOEm1q6HQ
r6TPRi5fTmhmTZGgar+UwRcQL6Fq8Ki1JdCzdV+QDZRzN6mE2NWW/xIInQGtQhSI
0l1ni2/veobyjcAj2Kb683ilcE0gIfGM+jnTTiv0bFyvZKcfVakMi8NudYBgbYPz
xACWascqeX6ebKg3gPsnbJRdsy1gQHsqZRBZk3LScsxGlizaIVGhee9qgKenotle
chztExivwP/++BtPFKvUTR3KTm5wRjGyrIg3hUjNfEpYdgAgkugdCNGmhqVtVYxo
kjs0YzG3F8bEJAlfToAGRjUiRzHvBw0jXiKuvQoPDIC3vQIeJptcH6gYCfvnYTbx
HNg2uiT0znul7MApE5cBst/Fqo5sJsXoo0v64TbYnS8vygqPpS38yakPNUAz4xg3
ECu4+5dgQ8TIbiti5dwWDFHECnFvWW26GFHT0jNkoAobaef/8hUFJ30WX+Udeh0N
sCl4Nc0HIGgYRgc/t+woN1AQVwBGfWHxH++Aa6GEu7snXurGyWn3Spqu2hzB45me
oOxN7761oL5uENnwgiSI94vkcpmkNJHHZjBnfPnBbLKyXdOL843cpBRHyTyW+95k
8hUvppGXdGrHOemJczvTn9U1r/lOu8AdchzJDFrXz6eGOm2shuk2D3Ial368BVe8
upNhy1nXbBGTf/+fl27xbvf/YD08gLRHDtrkc1n6P13oWzq0NAXhHTz7a/e44fW4
MevDVfr/jbTtszdIOVrt4rXAE5kYkEZ+aO2qcFvnreBJEGL3OhQBIbGQpPFnMhds
sC3DQNWwEayM1/FHNb6r2FiEX01z4gGiN76KRBRR5H1Ex/mrOQeFV3fKYZxUpS9t
TpY8PK7KVVVcBLFoLByXL9WUrJkZUY4QFvFE/TMbsl8IeQiF4lt2Fv6u74MSVLB0
9ACGH6EEoTtq6ujur+JlLGR37rD8r4BmpqtGeWOlVAgQg0GwbwiSnhrQT/b2a+95
bX8WvpAJgYTP19OGPLI81sAQJ817+uGCiU/8+dtK9JvgmNU9AeoMfYhSRzjf+JoL
rAT/Q/InDOjaNzfp/MRmJgUFwCDFVH1UjMG5XFNnjcuV5+zpVO8J9PJqvTD7d4bg
U/G8upX9EYzAXbvVeDi+N5CA2ckwbEBIuiPikmZs/XeAsGPXEsSmDBHXBng5kNgQ
gjpXR9P8MCKEaz2vD5h1frXlD4sDS0eqbolsXsQzx7sCquk5VY/RE8IZQQuhlYUm
SQ2l3vSL/mvR2RU9QLDiKsiPjIg2bTEVghFY4g23jFN++8ZCAODCOxb7rcYVG/ki
vgQK34aHq0Cux501a2tE4Q08IqM825volDsR4C/IW4cpxpKEZynEEdJmcK051+bI
R4uqiJ5ncR+bcWBydx1UL5oLd/S8xwSZeEVI6A1gujUGBnS6S4KjqEMae5hKOn27
bIFChJQzXg03Dllpg1v7k/L1uLAxHXmW5+JN9Kcjk18ez64rBmOBZKXmBcn3wfSK
Gq718vjw5kGqHypuli33ZtEIXLlv3IzRcLcSL6TtM5kkCQEfObXl6VV7rDjG6/D8
oH0wPHRuue0U100qr4PmX3qgNRsITPDa/RXyvUjg72fqGSKh+lRm3Otu0l5/QJHX
Z/v1uMKFUEgjSsbCznFEXzjvytGylPisuo/D9JAg4QmRHct3uBNGYzMTA9fHyU+T
Zo13jF1n6K1eSeQy4sJy6NSbN/5zHk8C3F91oGHJstfbuZ34GwtriDYdIfA9S/xC
NXp4wmz8MyIUbBTDAAQHEOrvyOGcL3B1/a9p+GD1nJgBQhCROvgoKUQ/gr4vTyQQ
QhG4WtkY69ohE8SGE4KLova/0d0VRBXN2oIMwCzdLIdhsksG0wtnKJ4ERcPyQBIv
61JsMYZIWDQuARZjz+NNMwRL6Iar62t/qNnzQbbL+2LDbNEbnXuU1XsF/kz7AwEy
y0Df6fJLIP65mPjj4qiIgIlPyQ99YeVfvtH4nbYii71vIq5HwpeWGwzMAhbextXz
4nYl4UXOkU0k9P29H+VftzDrIahxaGStra3Z7yzEz8C6Ht8EBb7Mrd+3kmdXrM5N
fIVA3dSpy+j01gPdP7yN3sYNPQNUuP7+tVWNLj7YGhByL47vdMxfrl5P7qMe4kqk
y0FNCKSkb+SxAW9D4ZR1n1RAzq6vm132UEXGr2eIc3xf4DlxcZHsiTFM95tUFDfv
u+dZ5NHykxEb2S3YRRgT/ISpj/VgbMOj8oXO1OZ7B3FoI3tE2W/Xg5L3LWrL/1Bh
Bx09wCndy6AhEGx7BH9SoampChcPvmdRG54sJkc8bgYRQXT1ALVy5aUoIgy5MvD7
tUf80PCL53/W83dTJ1w37qQ3MlrulKzP+ql4Hrv1vJWMJsZyzQjFAitZ2HSgbZlr
7gcFReMB8j9KXyTXRvrBm5FBsd+xAegcDkfFYtsLwmWDXVIY6+YeyD70wyDWw53J
UP/A2Ed5l16mt1ma9SkLRs19oVw+4kM0ECU4ZZiyx8PJRrz+jnmuXOzUCTDD2bjy
pv0G62AL4qIIDQ5FD5Dih0d1yDj7iz7lPjzPhTwKsrsNF8WRMgYpV7E7yujNUhVG
Q9QnLvRtx6ZdOURmx9vBEWS3/ASfus53TMPCXtMZNYVweIKd7QuS6quS5ikMv8Sh
RtymuyOg8mTB41+fnOwByRB2tTnOhXRpaifZzNvgKHqHpkrpiiuQuSXUjtYVq0jA
LrGcrVi6eLsubaJ5t9BvNhmXVWEXJW5jIZxi6iKBgFO7w4bg6U+ivZF9vpUc/JMM
oSQHWtQVPiukAugIzBasMP6Uh3ZOFzZCzKPSjX/bjjZzIcgl9IU6QsyeK38z7OBr
NSRyPcx8GpZj5zH/4Ic1kcyAK4uNhLrpyqIldEVj36tcAIZKcf4Z8VMlyvBTut+L
mIK8efR+sdFV48O0DBIrC7AAdcqH4E3zGkNSaWn2uXnyxu6XGL8YjuRGvLovoiwk
qsegGM0ES6EMkKL8H+9iA1nAmSApeFvWBYzHJtGSMn8KwOV+veGaltOsF2KQg+M6
0A9eZi3hV8O/JLpOJZbT2SIlcZ8axDSlihejbAqjq3KoodYpptXdriZGfu6u7fA4
xMs0OOeCPBZEva9arw1h6vlo1SMdsze8oIjMrirXeF+VVau8N+XgPC3CrCz+Zvdt
2VGxxCUwKCdoWsVGuc+lAr0zpAMWcJNjI+BGW+0ADyD5Pd+1aOUI9kTOLlNQoj/W
0L1E2WNYko9YHUTBipW8ShL7FbFWa2N7G6f/nRqk9moCN6S0Wc8ntor1ktm6UDD/
yKdeQ2MyzgkMwv5cVJxs//nDVSKR7d8iOg2i6aOFEtn/kZGubALlkB2+9s9gj4xR
aTeFSlSC20kiOeYUxh0YrVqr3vOYRvOGC4DngJms7MsKcYjj1YHaNIZAHuJky8ia
YRoIrjiefkBpULRTp+OTRzudwchl4Rpv/nLu7pEQC5DRJHVeX66pG5xdyglKq71w
8lysQ5SqU2ex0soPvxPSQ8vjhvLznYtqWDTndNnTky2NNjsrngNLP5qsZ/s8A8bF
Y3r7J0v9VafAyTIA0PgFTOyDt0O2D8HM6+t3jkQs1/LNTQ8CPXHBbKszFGw/BMEq
NKJgYsfs4rUDE2s2CSHF3igGp7YJ3zPTd40tl0Ze+71l+QWEnIsxyKwBGMpJ+AD4
fG5+n6x77bPhNTt898po0f4DjCsIMuJeatNm3gSVxu90Pzqq9aLrjF3oiZPbfuwS
bhDWKKG3ohxvu/wwAk02le/dXjpUu7b/Hcy9j1ZmocG0g7ts9PL7BDe6fcIqQrNT
uMAO7boWm42A4Z6t18bZpkR5A7rnE3KE8L0D/hiFHpDZGplyBEKEFq/ecILo+Rz2
QPKbQUhMl+gBTq3LwFcmv+KefR7qBKrblKz2MgG+uo1WaMJFWzOPdCV5Eyz3EbqD
yIeyiLgwg0yH5BQ6bCZJfOqHFyjQ3sWMuFZiOopDoqY4Csa8lFZu3RujxG1OWH86
2QNeVcEUzXVXCGZ+YnlVZQZutbAOgy4pGjCE+HGFqj6YOjSgDQhEKEIsVELIqW5G
YtnsVwTg9AUEmBX8PlOWf3Wbz+kccDkA3lGL7Jbkpy2av2250xqYlbroPuWOHuy6
bHJ4mSaEDPzZ0eGSZa2ruZsgfF2iSIeg9a/A9C6yJSRxY50RYKdgsRjdUMqEQLsQ
5AvTI1NQpU41cRcBzQPjPbqTG3kRdWg8f4zzyx5/ZsYTKbUh+LC71283KvRKMcSJ
551YIcYHU0x4F1uOyVbf/vW31JjvcSO+SvTae7dSxTfILNK1vVIovh3Uax+bN9vs
H68VyYSEK9zkyc7sOP4J+Zzz5xrHw+uuDxt/TZhxLXd87VzWi0NbgHAMDhWshjkU
XB2zN3Ji7HDPZDbCnOPGL1ETI5JL6SM98Z/QM+eu0vlrfp/f011NGZSn/E8ji/kT
+jHbC/9rErQuLl4/Is/0u6/WX6zlBGWpnYErYncXaGKVKnDUOjGMQIuaTy8ytom1
7lz8gTAylx8V5WlhOE11YDa8sSQnjb20coqCEMoTJVQ/hK9uAxxDnAvibOsKU9uf
qY2x39eMGs4rr3hw+r6YaY7CjuEJeYAL2/BG/8Ez9zQ4rCPk3dvbXRKs0LrkzUBX
k2XcoTNQO3h4UFFt2i+rzU+ywbW/3kUw7SH5+971UoJOwwyf1foXly7wl2efSrsw
6lq9Ijj+0RNRx8uZGA7nSzQDY1VQltWPseWkXw3NEY+Op3rUuLBvU8vTt0fQCPSz
XGad+DNoPX2XDhIQqAfF+7vs/nxUjnLIDW/RfIfXAfkihBv8NlEOarUDiWsT86uI
EWAA+pd845XVY0YHR5pX7A==
`pragma protect end_protected
