// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:13 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tlPJCH0DyyNrWv292ZGVIMUhawD6YlXuivNyOoIJ5pHi0aso+GxFktcFZ4MK29Q0
zJBQxcSdYRjyDuJcNyF9rOKL3CCRMQxS0qUz6CUa7myDcAYQNP0quEC/BeShYoJz
97tm7UtH6CIqEBby/DDp07Zg8Dzb1pJEBlY0RGuNHN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29488)
VBEEOS6S3bhJ6ohMmGSPIJklBp1i4HkkNxWn/yTemjfi+HTq0eDN4zMqfwHk1gxX
yJparn8yMz3+yvjKtkz5inHwU7B3VFYQfncQI7SFArLeGBRaUl19Vt9TDFb7Kevd
XFxscp35aS0fm6pFm2PQ1+HvrhlkHS7XcV30weE23ZO9buoLEbfv3WBhe1rMLpjC
etGqPoCTjvWHaH4hZkCb81LoLKYEUDnK5nosF8ug/Ps8JVhKUbzEQ/4i8677P1ei
zpRBXkBdbrIXMh00pmJD+QMIp7T1TgFP1DgJ6bQ/8mBFfxjZ7wdZ998eWAC2ZzA/
Jy1Svnjmx+srOlhRs7/8HWGMiRtIIedC8J7005R6KW35ioltAMvP01UPTLyFchs5
sujXX2BInEt19ZKqMElgBEqVSN1UIHbEkvUti6s7m7c9EsX/spD47b5bjKKfYK6l
XA5cV1VM+t7kz136DXzM2WrXfxD3Vhe1T9dch39cbZ5hHqQGNYTW/XX3x/qHApNe
8js0V9h6pKZIlavgFbAB8mB0FKIuth5f0cXrtz0BaOZpgBjMRQ3YOevhDcTo9pzz
9MU/Nquwc7c+MenJ0TgqRGsUXHh4I8TkUcDV1B6C2nxfOkz0QGuMCogAXuTdmNmx
UjwfdHvHyMgPVOgR17jkyRK1m34Fvprrjji8zP9S0f9jog8rXU+H8SCPMcO53a9a
UNSZ4cn+7ylRuB/BTwF1aFMABLjL8z1Ty27s9csGHZyuE3S49SOVGsonmKEus9aS
Har0rBG8NbMRkxHpOSSntWbTKoK3QJTLQUdHh84AEISm9mEvesJ+qXkbkWuCa8tq
F22NdoQn2oBjvUbajV9umDwAIdthI3Vaw2R1iq/uNbcqC982VA/K/H3wgrf7n31F
hr7fEdVrlaiJ78gATyXR4lSUjoKld733/ueon7aQAu6YbQAP2Mtz+YsEqW2flcvu
lr7WV/VqbHK6bjrXSXyE1/xsbBIACGbNkxH9SkPHd4HZ/6u3qfWgiUW9m09E41f+
6m7+9lqUCu0LccMwMN4BMJh7+U4PBkjZuMN/WAA70kXxBaO9G5O3KQtokYwFujx0
mPFeWpyXrYzyEIVXHC56iLmEwBlhkOhYuNG1zxtx6IQ+BEfBn95OyhNkU6FV6ouH
gcm1RANnw0edY71yKjHOPHjC9pjvICNV/okv0eNV9AtONSueltZLy3Vc5gnRsec0
Yh1bxKBAVwYqxYsTgYfCagZXAVa2nWra26lTlvB9LDWHHDqw0zzBxC1oHCCzstr1
evsFoQZu8yZVBZdo8uiNUNKsmfy8wMUBJGhHDleRivRg25pdgWhjFLz8ioUICk40
LrT8T47esaUeQ7b0imaSwcYg07PqjKC+9R91GmLLzMC87+5Nkv0hZ9C3wTzVkGY5
AGguQ4z+QbMg1fD/lggJ6p1U9HnvOnDhEGqQqqZlYnrERm2B3Ehb1GvkGvBump6X
6iNQ+Yq+PdK1iyaY72TlSrX8jqQcdmOh1GzZSK+ZKFdWe029ju6h3m1wtWxw2ppP
cOhVKSjyjlhUsiiUTT2XZFQBWXxz+sYN9srSU0ddjp0F9FX5MVXpakGDjXYhuTXg
LUe6Jflo/MLiTIRvjXWQw+TOJWBn0mQJUz1FuUKzGhHORgUO85N1tGiGftV91xYG
H7qiXA8ZtjZPxjuVg2Q1od3ESqVK2hyPAAv3vRY+jMk7eDacXMpDXrzaFS8SvDYV
TFz4EWXrMClshwlWZpMkuqYGR1QifsS4voHQ3IkcARaj3G6okuZiRv+hfUE2YKY4
avGWvNEdd3Nn+I2iDDI1SBRI5ixkxFXHUEXP3YxiFt8zaZDlWlAtOK66FVnQA5jH
J2ZIYelymKwqjYArXWavdK9HEEVhoTHumCbPPtkp9w+XM7eqCckDXOl0aAasxKBQ
9eB9rOiahpmsUMVjAUjiMBITAsXJa4WcBZSi41VONcNsPWWZYv77uI2OZ4DIqD47
xrQDG2/NQuHdZH0yNxgvjw583rcGVp+JgZphidJaPSw/xhYnoidxKOuAKO3xPKgP
b2soqXF6XD5A2//OceyXdryrSVEqZ+H0ApvWwSRUKxNanYnIAaC6ZgjrO34FGYLc
+UvYKYiskOHAtq7fZ3REKGM09nHFd8qL01D+MOY7uc0XwSx/ONl+BGdKMm33UqlE
tfo0UZyQXOyfPPc0qLcpBpys0Rgt5BhGWaRJvdL3u1Cb2iRds3okBdjDCjAVtpFI
nMYjeA5m8Vjo2UDm5oT3WZ/J4jtzxxQU5FKupdS3MnGQFsnn1Zkz39357Ylvqoqa
dbcjnI8WY+Y/48f9f6yW1tyMWr93Bh/TqQvVKXYtiwGlLNE3U6V86hXyafAjDBbs
CL7zCYsVdnghINqh4jM5wpcu06sOF8p0+Y1RvLzHttGwvJi3JbjlkgSJ9rDjnCBC
qQvG35TzUduPx2XJZ1A5BR9FA7jmViMORj+h7ULE8hwlYBcqhvSvVFNOXMqkaXCY
KRukSkd4IRRCXyl3osrFR4fELUDJ/y1FoXH9tQt5QHMOehak3uICb/YWUv/uXoCr
9DlDj2DGcsFH+yLG0yHLmmmRdFwrg2gcCusXJWaZ20SkQjPkkMjeuzjCosmaZzLG
dcc4Rb8CaNJCRADqUAKFTkUb0JWDwYiNoDYF0ZOMGj5f50DvYjrk84BWOaG9vnpw
agBAaBaN430WAdiZ9MvNJfKWHvkAbzOosGyPfno+35isfcoBn+QeMuz9uXF841US
sOtO5BYBXhPk9VR2L3Eb9Xx8UA2eIhXiq7wfQwwGCVGHxdXpq+ChOBPokc+7Ofqz
rrYZcJvTWBOJ+a2jex+q7QtJuxnd8sxin/s0nnhZJKNvHbPGKy06L1ws9lUyKTVR
0SD8qEhmbtRitA+nUZtKt6tK7P4534kw6ZUzR2OqWrRcFwhJBomHR2lXq26Oaw0p
izOSkn3jRS+/zlj6j0EbUPe7xCifDKAVtp/3o0U9b1UTvlcdlmj8wwFsVExQx1nu
l6KdRcnHZaMS/3Gz558TVRbnPwABA8Gekhp/cBcHjJDSLprmxmPoxJnA9vP1lYCw
mlO980FjYXM/p8rclG1dxX7NgrvpJAuFtn+3DEYTg7yJwubKFCew7ikTq+kC32zp
qvVB3aB2MXZPp1rJyZENBRWOyoA3Neeb+Z1muCK5ARew0CUlAB0MrmOdXP130zsW
1ZUmHkVSFsFYGbr9cskOdeos55GwmJinDZwOSCwHosc80BdFyvW+XkQiyhLQs9MV
C0mBJO7Pkc3aneHhHQCEDGJpn1OSOzX380BuXUACMgSOBHGTdOyCyDeT54EWlSEr
nej6VLDMBeTN5Dtyi5JZkVXNiyL+rom8KtKJgQEKA9dROotlf5JSwBXJriUbl6kl
NXcpcVUt/OlbMdTnWlZv8tqbNFvk+lkoW8ykzYegfEAgOdPV5wgSe88bEn2QxfG1
2yBAt4cS9QPW2cHjZjJSnrM8XLXuWCbvaUJNm1wD2SG0JPKM5PDvuIOHO+oNcRjZ
8IsslJ7yJyK+i7SZgDGAcktajtaixnkxGuOAl9dEl5ncsNWafrdPdswtMorxdaCY
4S0p8fbfP4ZmH7slcZYGBcbIUUwQVYg5HnJ9HmetJdPfqCGloG9cpfzvTvMqfBYZ
0Nv2cVU3rezg55ZGqzxTwKdHaQJ65Z9JjETWTdOXQ7Ls5IaWk2IbWbFoJWpxux4k
F1E8Od/slXBXGEWhBE45bw6I+s36Z7zDxtinKv1vnsv+v0d4Lu3aWAvy1IteB1mX
tIij23CtEy8AI+3baVplKGlFCR8Lgvh/qsauxu5zzmVMWwU0eZD1NRQCI5Ukml0D
LYkLRgn0ONn6C4qrQHPXrue2gZej1rOUHs9POP8w+dpoVRobm4cKYYaBmEqul07I
mGP6Q/zQoSS4Xm5/qYAtIa1TYXKSnbG1E1i3z8WDQdORRG/XNPBtodYXcMW6BhcQ
FmM2vWASXILHVkUsCmU5kZfRwMb31/pBu4oQhwO1o+7l0DjgZaXhREn6lvuNTuEU
M/Twyq9tPpH52YsOXMaTaI7KOGlZvV+sdOJNDm8ozlU51Ejsv4bp5B6Ww+OXInE4
sH6ARk22uygJ75SPGgWeTv5SczZv5auGG+T4mxL3/94AR2Gm46KsIP0yr1EbIoHb
aNLW1NVI72JZTCgnE1bSLJybXKFrzL32xDwXVMlrWcJ0wFGZeezqe4bEYy4WD5WT
Qj6EwsE9n/i0Di0e8LztHJYAZEXRU8Xm2gynHJRrw9Kqphli2IC8ufuxJDLybaIF
qWMrFDsJ4OKUJd0ERD4GdOYPmG9fW5ohLMTbyjhsKbpaZbzNRWOapneT8tZcv9xe
NhPBoj8bnKHexHmXBwxi686ja+QpsNegire4EGqQwhjzQMR0oi+d4uFf9ZLVur0+
jVo+xcGXhZcZ+Tcb2aCgiyZ04hG7D8H9FUau8DqZtF4MMOIm2up2DiLSKQHnbLU4
+Asvs9UJwg5Uf47N+9j8eE/sogbcCbDGKnUbwNaL0oTVdrkKWJ30wLAK6mGgEsHR
KJ9iYDKebMdhMmHTyK+jYwQS763ubWjggFMsgZ7VjlyKlon2RkhYtGdF4mS+dbvi
NqFpmnjCgG1wL0QggDpLgd5g/RsjYuM+oQI9xXqffB15CjBnCMr/VQM4xlROrlZe
t4bRLRaKpU+0Q5cQGoC1njbGS4Hosiey22LDbYs7S3WB+eN+0dnX1dW2CMWLyL1m
26NJDtv9HuHFlh2F+KcBCV7f7HM9rYo7x0GZ4P/AWVzYWzcepjVPGrkgNYs2KbYb
VeivSEHza0hoqIPV26q6bYDI3dgNcwBGSTePx/oSfauFf80Y9pZ+hYlGW6fVZA3z
4452X5wWnAPR3MK4xWJNKVSla7Fxl83dEjussftOdi9KO+Kp/U21jwKCriKJwCy0
XyE1cUDXUZx4BXW/Pdat7ORoHl/jbRDUlJtj1lWmEDSpVVWk/KixVgK5sNr79aC8
nhfD61ORZesW0+KuXlnbJvXb0wyDfW5IOGV1xiahfeXP2fyAIWlYZnvoUX0KQllc
fm0B5kxRp0K5m1QASu8VXLmKdeFyIsi41LtGpLXp+7fjEIOEt/93xPHgrTGY4qj1
t3SDp1aq0l3wFEmp2aqwKId22fYu4UoB0QH0WWVLvWcpu+cn0Sg2QHVA5hWN9z7I
tG4X1CYoLoptXYWJvKV/I/s8EMTcrg+ybb4DxkLbwU7mVkfJ8gLvVEFd4wnU5KWI
8bCJv4IMvDD5IxnqLr0IiE4XiucrVBa6/vcpwtgIm/1JUC3lah+6sWkDj4wsRP6M
8/Kg94TO+2VopDCoAL36vxA1mJsCope1qG9Isz7pQW7IxQuDZbIrRyWWKO9dcTn9
O8BcQiotoer0YUYXaiKP5SWU11rrcaZGM+GkYlRmKZFvHdyGW6xyfOaVATzoPyr3
j5F4GHnCl3A8vv3IAi1jYcbOiq7uHri7BB97o+plPWdR+PR7auExO94YM47EpRG1
IE6mK/4cMn0T7BKyMq2znNRxQae4c84/4ZEVSviXOQofI1nudfnCYTRB33CA+yUY
C5mK7ETCdUML8xBDnSx2i7hSHXCpgdDC9SdGqR65/OSP2wBkCcZb/JTdN3fEQcwQ
d3Vg2ZqJVK2Trl6yJoAPh7wJZFydBRI+jb9R3259kozGEUiJr98mawhbnjxdY8ka
M97ca2WTXcf+GiuhntyH7u+0mg1pEF1zcJPhvG3NBC7UrsK+mMtH+VJJTOFRqVAe
72ECldKKFspdx+IJkdwNpkajKm9SA1rPSwy0j9nmHgujK9ScqZpOVVxpnNAOLPSa
QHTAJ635iW1OPx/s2ceo8K41x121j36166Yq/npESCxgSpzhf2NPI9+OoUip8spN
SRn/0GVG2Kp9EQz6UuuWM09+nnfrAzKgBHFPvpJMrT7ZR4UuRzewq04l2IC811QF
O8zrGLp0y8ib2kj+9f3QlZS4wdJgxARzmuu5+utQ/gp+07lM5RQgZsgy0OLejNH9
kP4uelPwnW8+NYQGwol+PqtfqlBwprzPnvdqYRaBgH+PjU3RpG57NDANO3vHn/R2
ZB4HbMVzZ7n/pNHhli1L3dZ39NQ9m9Id/dIkb7nwRcJl6cxYyZuVKw775Lxz5G/7
Fb8zgrJ8V8QzKiGNA36/JUAB95+tbWTBmbUH2HjJhcFMP7ca/A/nAL8aQIUjow21
wfKqwimZ0xazZhHH+wYB6tY3JRHPQq7D0lVQLOLckFGd1lo/gHKryLaS+Xz+QZO8
6YN33xJDu1t4HPQ4lAer8hM+L8GDfogif8/1DSxyX4O9iz8mlylvSurxEwKKqtdt
khwVy5kLgErTcL8wZ1x+DUG49+RlAl6/cZVBKireXs+dYVaPiX5oyYixcibcVAGR
xX8UvvLD50Bck5W3nGSl/KDKl/nyM1/RnlwJSBGZFYY9YHHEs5RvFrNglqy3mwWJ
ZsqlAjMuYxDAMI3bwM+ufMDB93qEeuh6LEWsGrIfmUw9Yxx4Z60sFAu6Ei6v7+3e
SaUwzImOW/kSLW8vBNFOjNGke3xt4zaWhgJJomBBKnZh7G0WHLL1Ti21kZh70prX
BIts7XAAdlIjxPnhYfUeSuRPv9qv38wL38Sr69BVe/tK1MXwxK8bnujhbTcUNkjS
b03Bhhgosn6k+Yvaeq7mzjaCAV7eZNFTEYLsOMYN6+yr4IVE15jd4AWfDbdgLXXH
awOZbgnQKPPjf73jEAqZcg6lSFStmExTW1ZSx/n1EK4XN6YL93iAGrfLN+1n6cnY
Z20tn7eV/egdBSlL+nb6IKriGIkQDSugniPf/snsrY9pUYNkEyWHwI6vceJn4ttX
Je8XXal+jg1uNFAZ7HFYA1sDtFMryf8yxmYcssGjE7CvrsmVm5pXO94/1qMeL+Q5
GezWWQFmWtHFmKdtp9QhA+b1i5QQpTHV1EBff9WgoWXsUMVE6srKFKQUZmz+6U1j
uls4BEJDxU+ppm0NGmRSdwep3juAlmq6lU+OK3HWayzYPkZRAiLLPvsmRSOcYCzr
5nmZDsb2R/akYS8rs70A0UXHKwOe+O7frJUTLYjQ6RwHEEOstUt1UaSRGO2CzugA
HHMZRXWUk7Fti19fDnJ6xii5QkZsaGED5QaYl+6Fe9u41jkDNQ59n4p7rM8j8RLA
5kouKvl+BuWnRdsCV+0Lvyg2+WXs05trqfk5oOkXDG69cAmpoHnXoGelvhu97cVv
KMEb/LS+/YfFN8gOIIhr2CHnRMluSCU9K1JHbycVQ88Ds/yhZu/lGIy8J5yilzET
SApyWXYRVMMv3ziUIM1rusoCJB5Hy5SJ0h/ipznO8V9nAMYGvkNeq3Macv3Nkmfc
1zJBHOClKO3I5DQD3fv1BlV7mT01uIW762WtKgt2eb6AkqxteOqZhfA2plkHUzy0
Ip5PH97EkdznJrUPzYyj8kDAK8uFWyWwTHM5u1ostOkspC/1PolOtexTZv/ofrvP
91JEqmq23pCznBuF0C5uapwd8D9Rz+WHV6C/MlSnQWQYFV9ZO4XXBpm85GjIZ+iJ
UvH1T7eYwkwYGQm58SKeBuuWZU+bChcghkQdPSQIYeJeiNgndUrc/l3n6Une/I5/
E2J1Lk/1H1mqtYHqtQ5hUUq8Ao6O4ZLzsSrgyZNkRQFsleaD/cARFn5cJR6hmpm5
Q+ISo6iBtRQUAAL05UTR4Tq/Gu9xFeBiH1ZYbrnIRUQEMiJSv+w9t73b7wxfA4D6
6TdaLgeePZE527H804zEbbkB4DrabQ4/lIty+QFLDZtrJ+9ARneDeOzkWvNw5u5N
Kk0kqN7JqxipdAXBODODozFKVlXAziiQu+SqP9fV2r8nw5EivUSFN1mw21+10N0B
eNpL35crhjA64DgU23EImB7pNzSHAoUHkjZTsKZa5qUAKjFVmdiEUbIFHznQokHY
cJLooHbwd3XvzbUmINag4+B7iN0cXNj4dc4Nw2K5IZooi/Kq/hZJTZ7KUMRudeiA
txSgXgnFhuXo6GvqytaqOd7zjdDLT64O0RMH5YaZs2jj8rymSLLHm1X8uwe0rTsw
gXAem/NiMgH5GbXCi1bxjQ0bVG7peif/R8xfEIIXkpJJQM09Rp1pfiPG1TUGwbcL
DF4pDKffZpE4eTwtYXcORX9sWt5CgrViJ6+VLPYivoSE2+KTMzzSSOX6+uPA2aJs
gFe9fSxmpYpoiyQ8uMAb/WWD4P5vPHMjdwHlMjuXcan5pzTHYwPlQEp94VEJqCyC
Zgpc3oH/UVY60iEAsCGicRj9wdJdhEIv70Kmp5sQuHP/ZHc0qypPDMwfTpRiLu/l
e5+PxpVQ+hPdFZeAfneuQj/B+/dvbY3WV3yy3UrnL/Qbiw/ibkx6W7iuzSq3UI8+
5eGYKWQ/ctqW4zowCrJibyw7PuzzDFAy3qvVhM/R1zJMeEqqEdIFgMFqGzKsZbvK
vxHunZfw7Dm2QdohpK0nmXBESHwcgqhhk8pippxU887nkMs1qOlAAhCjocQ6Gj5D
UO54MaSB8VMyLGAjTyALp9eVBHv+VHVuhCf5t5ubhsI6OYKR+0qZqZWiEYJlHa2g
bmUj1z4mv4ICpLvIvv/XFLuxo2Zbbyol+NSvC4xybtbJL6CrLXWay/3DGPkIEN0m
BjC9EQC93DFXtnd+A+U8onsQL5SZlryHKVR253XYxxSg1MCJld6cZ9TlAm/HhdqW
EkjmdHy2t6rHL+Bm4gep0vn+jx8Gc6g1Le4GxOpTNNTzGLzL97CU5judu+kSD1Fp
tLa5kt/8zPc9TVOAeq16yoAdq2kSOEuBtzTWO3fkJ4h74Yvxh7RCCMtxtYl11/CO
iPDb5Ewr6uqQJcyWeLiOJazH+Uni3bsZalZt1Tp7d/uoJMntio+9LB4HqbVrz/Pw
LdFceUolhVMsSgSAgQ9nMmv2pqM1vSXUtKOxZIPzfBxcWBr0fqp9/vhfDVKYoFq6
Xjm1bKbcA6S8FV+t0hodk4j7r+3zlK6tyY3uqThuIOF5W9Tx6hu4dmjrzI/kViAi
Oumk+X4SRqXGKWcATyXT2YexWeB9yBy0u0rf9bBZFvlFszpAPotQQfcKz/BM6s9r
OjqxIgfgYDcbq31lG1vuY6k1hhPIIQFJ4iLuycMauP0vR6vbKF34vzz+rWwAQbfg
Jn5UBt80SnIMMsfVMtx75XLlhSzsecL5rXUcT8rTpl09DckiolgGpxEM9jwHiaQi
ZHGCvFLfJBm9dkJMBaDf5EPS0cAnmxC50SGOZla+16XI5lJT5HjP3ECnUYU9bn/m
CYQs8Kb5Mzqxo71fmsdgtWtaSQhwwuwugAsR+Zx6HaII1PEFIxd8ZtWmPT7P/LmL
rLWzotUwsTX8nmNS2PVQQv9II257bcKibaVPxkbQGeDt1PbbpP+nNaqc4fTfBYDO
8wITkpVnseEinCbdvASrTx2W7e99VMFi91tYvCJR20JpF9tkyuBNyg/kBVYhx+j+
/6g5GaLBgYlRCiSxUPKols2jpJ6s+AhK9d/zya7Datw+4kspg3SWqTum3XSHMxbk
g2JFnKIn5DJGwZkbswij0+heke/j5DCxQNqmxZ4sC0KMuO0Yc2ef2es+/1cA5Qyi
LhyaxEepAE0n+flqvblQOJMlQTWryaTnDP3XRY4ncL2dHH9+MY78zd4CPtIYQpYs
gAzc8m3ZoDPxDpfwTM35vtPiinO2wFtE1uazA96fn1f5RfTavSXdSy0yjFpKaM/r
i8TTOxRNYGUbo5k2U8aoGvEEH7DDeASIYRhfI1Kx6OtUYcnhgPYv8+8/V0AHRkcj
gdGir4STcIzW3+FUY0t15o3Gnc49So8NoyN4gLicHvDXMroXPsQysFpKQB7FiH6S
uKdosBf2RCQpaj84A9blw8cqchMRbM8EbOiw3k/GHcD/nl5iXvZucuUCJJa6Tp5V
tp0Hn9ywAhqmQoYrlpnFelcRQuWcjhO2u/0BmQavJ+SWXU2RIDqbQW7olLFkR0vx
HzBk1Z0RB2kkP/vsBFuJEHriYKekeREACYg9JDWmbskSbdBaxIxthGdId3BM5yI/
Ah0iPlFKCDGvXZIxpgid/tF0rs5/W/rWO3Gf0fn5IuQSL3vfKcGPtbdDAfHLLp8f
198Op29eKxq3ZGAF4XIaAz3bbTMZaHINuY1dyjn/uzrcQRH1R2nXBpv6wkzhB8Yi
LQSu/mWFcLc+ddHZ3vS/eflZyTWgufRcszCF/MJKtYDRaJ1YHMwOVqgS7PAI0CJi
jLzjgPVri72BUEqy28mDxTzUxJ9Fl+C66SJq62+cizQvL8/Lq6AVf/o6Z1dsiA30
O6/KHAVdwtQVCtPPNmcxua9lE+z9z83SEOB9mGanYSm64UuQF+qhrI8XbXU9sXDa
J5ZKbHcAyMhGGAl8HFaz5eDL/PT8RepNvuVJz3+gnFApgsG9eQ+/CErWCvg30zqG
qJcL4lBtmMkfcyaFkA682Gg6rz+JbsZuXzaGi34wClF/L2Co4UO6EHEfCFNV31CP
pa6qO5GpYAa/K8G2gXOsGhbMzZdVdDDGi0+8hONpuswtL6BDtB42toMvh+KSXiLv
kK6Ws8FPsKIXvvgy69WlCrySWnfCjv5iYk1ksstC8myVX4D4fSl6cYq2RjTNhXZ5
UpzRO5e7WCJmc6IONZQx9jrYIElQeS+FCU71sMojt32o9E2vGJC1umLI21MSlgFW
trs0rOuHcXGeUE/CmouoiujPs48XZ/eCjAsvMMr90WvHjHRbN27mL1qPnmaJeaEY
yh0ZqlzHQiJLerjocUhSpocdk/OTWSgdw/J0PfeTu0v1G34R0yavhbljrMf4CvJO
Blf2t4yY0Re+EjbNqMpc3MHw8QwcfJpo3JZu+FOuc5iecGlsc9lAkSpyJyBqwK36
yBYtFbHuqCGD6bZeFoFj85CRvDrRbimPm2pviCRk86q8rKBaj9TdCeMFaj9xVMlu
DXPc6iEWBhzfNgXxfl4Iv0boAyaABk7MCFKRVnP/P9d223/S7MLd+pPAh+od42wT
unEpVASP8KLiDy2J8YQGrrEoagl26Troob7Tg8D/jFB5hKKRw6B4ASc500t6t5zU
k/ZlS4RTwIx1Mb3IR9afjPlq9moFsGjLnXliJgELDDvKbwZQL7ZluIY2i3ZUXNip
tx+qtfHBQdfYNmg2r8fzR0ONLyPZ8ZymkJ9pFC8RFsZz9/idutXdg4QqfW3RIHuF
9iPz763clcyyHVaYJi7ctugVWdpD+Sact0zcVkLhP4CTgxB1qlAAjH10SmUcFfkM
vvfICiiCzB5i2WPxuYJH24n5RV3KXbP+Q2/aGChuHp9sNVw7tuC35pNjc9KrzatW
GNBVNJB9NOyGdDDHW3Ty8KnXwLrz/OTg49OrfveK8vU0VY7TMMiyS6FGyRryPO4D
IbfXTroH3yESazON2wzK0RX7rEH5mtS95Pac18oLaxeBulOvzatv6MonE9sRV0b/
D5CdeIZrTuL6ZRRo87KxANbrvlb442cyMK2kQjdY+dHBt3kzPdN1TZSJpfios/pk
BMWDJvSnxUckdKokWq5K2TN2kD+lTHObj7pxn4z3h1KWuK0nsEN9URELIgx5Gr+R
tt5rP3Pb9yacreif1DCv88rKg/y4nzHV1jb4vZwNM0t3aLIroBzDIruGiwX0IelS
QozpyifmaXODd1VJ2MdCsS+zZ3VsZ/KkX8GJaS2NCwduykYVVe7A4Uve+wryTXRy
Dba/bttqKn6pf4zxd7JuzsAI+T5x0X+ooBXf6QLd0Mc1h4rfofYrgUSQ0JJxQAEm
NicZx1qRB6LjICZpkVnYkQP7Xsf8tQQsA4tSFKYVQx2ayc3NRVSve6wgsj/2pvdB
PyzVUd1JA25I2Ad8WGEB/qL5k9iI18xZQ4rEpsnFxqZhLG9mJQoRK4sFeNhIm2db
jhDXbRGxLzLE9qzP9yzXMCq2XoMD+A42lYjTHkRvCnTS4Qtm1mV9qXYA8hYikQsg
E0fEC6hGovTSerBQLswtbAr5oa255uOHzyp107dG5sheIcOZBjblOPL/WehGvCda
O2Zr58dmz7exUemgRwHz0GCEALIca1J4+sspwduJHOih9kCm815VaiF2b5B/Vz2S
rOHtX3ZNMgG1eOiXideLUyk/0m64K2iJfusKp8fTDxC3JPkLvmoMhTGVuff2WGZW
7FX88p+moT108FkU/NQ2VJOUMq5tEIxYZU/ZYdmHJU7iBth60lz8FfF0DYi1Pt1b
h+rl3Ui46B3tOEeWS8SJJnW8Mudy8WG+Hdt3MUatzsEp4bXyN2pBqGHfy6idYzDA
/2B5W53A9qz4gQH7aQ4W+3uriMCCM6B77PC2hzlYhrQIjKPmbSYsgnOFxrBjNlHe
/jsuVdsOQiQFwHeeKYp/yTYFFbvEMgPYlFjFZ1eFddl7wSt6ko4BvoYUK+UJdZ6v
M7XeSS8Hxd42wLnV4hghQxnPqYvMn5w50MormH4XoGsjsAadKfCxVruk1NlFvRi+
/sVgrsk4YkUvhe2rDQn/nnpB2xdH25zIOu5uuBJXv0PEVgPpsm4mpqP5qpyGMtEm
5Dk6ebYccpUDyL4qw1xVjOpC2yckgmhCRFbp/UvBhhsAaQjUGxk1wCtaJ7TX7+FW
OcDRr95Ak+kbChTzcxBwN3LeDj1YnMSt2hcKrD2tqSEsOZHQ/rF8oV+EkFqd0DVh
6mr5ZV+8Hbjk00wQC2gYi4Wg9RjwBlaOGGuW7g95WqTn4V308yG/b0czWNGCoi3P
fNaU+IUPboMoHnxcD1tXli/M6kOr2RVhAhi0ZGYScVb00ANGsgsLZMI3djOQN/Xx
gxKJn8qOzWFRZu9/tAgmJ4udC4dUru4thVgPFJryvd2mUf0xAkwTGsVQeYL5LAkM
nJDD8iEHQSEo8IxsyxbS/uyDSXc8INqqDQ2r072Gukb6euRteLiAHByKqplmzOIy
WnTTFqQ0eU1ZH4rPXgbVg+VqvoulXA9E0jombpFz6ts9udUh89Lm6pDmZ+UYWezX
Wzpyakhd3jfy/eOe/p0MkDuLv923Bb9jsHlueGGgTNA5L5MGvRqpVHyvRlIRTRql
fNqnd8aD3ww1D9wKJTAnf12mD4egiO75S3VhRRYAeNp/fsDVP+m1V9LThQEnS8bQ
DMBPaoN1Zh0VFKs0pxYDzCamV6p77w+TZaEwWf3ozp/jLApwCg6SFlO/hgJb63JN
Sr3VwfqOWPDzKvkXOiIC/C/4wKUiBku/EYequLJqDLZ4S/ghQIqIbzG5jjPclvAU
3nMY8yF4omZA8jkk8Olo1cLlOO9eqZIzPk3HUV7F6D6n2Q9L4HqnIkYu76hEaFW/
YH1ITOaZIvwGo1yWO5EfnTl2Oe+vhx8IMvZspv0LQVdCs92ibIttwdcjX1FpVdBO
1z6HC8KmmXCSqO+cfuHOHufnH0ke+gci0hFkoN+mm7OvEvyvnfkD4MaoiLXv9LKk
8bsjjRsY7HkYOz83613l9N3vflHFhUEnyq5BuCTmNi2INopFlFfaPS6/ZwFPxL0b
DcTIafltyQJS3+XUW1Hq7lNgqQj4lP7YcZzawochQ9P/XkOaJoUJr5+AehAFT8QN
gMIPV0IiceB+jKLsT9gM9n9GBMaKhC+ZKo0O+S/JshTMa9sgGjerNHDGGR6EHh4y
36gPKG2pmpcyEI8Op0dd9ln0E4ykWH7qaqujbNL9w2YMtZRYOTsyzb5U830HbHPB
SJE0YGWxJ9ncj4zD0hsB/fbd+4a9C2w+I8s8lsbCQ0Qqh2KtLzHpCWttzkq6N9SL
KBXSvx/f3qbawOuYGw2Jk9DBimzeJ1JKKTgHZZ6LOU2XtxiEI6ORzoYuQIMfKRyX
QP70E1/9MPDyY1u1wlLxA+Vs9AYXMyNbu/Y6eFHan+n7OQdswGpF39yoy5ZRb092
7GKWC7oe1m1YWeCMK95uHf0XTxwlbed9A6yDyBAP9csbcQjx6p4k2y4//Dw2DE6i
2cveWSVrYs8LP0gWYiyLpCqtRc1pmkuWapuoqL0KazbUpjpLWN5OwzpBcnaHpDXu
Dvg16Z6s9K3TWWa0PxJZGqOd0Ri97TNFBO/uwJHGDHPkP49M9Dl9DJBSqtjwvs9n
xl7NqKl8QeJ39ut7dtjctsrQwtAl8W/jl07xB5AjnkdHQxGtUxwmrBMo7Hxqhj+f
Zinm4RNFWt+8azak2uvBmNagYzEkBv9nA/gwp1tUGilarxsWhvjtfyL+00kzVMrL
MjpeHpkQnLBJ2BmtoYhaRlYcIdINY3gnXLeLyqlo05H1nxO844Bx8cjln5DnBCqL
I/bQ8EZZsXoLXBEp1OuVe6Cuh2JiS6h4e2WfHw9pDe9sJH4POSvmK2khq2wZPTmE
MWSY1tKptqWK+VOhOHluos7HJs4dEb/MmL4YDH7nBOfeCcwVcH/xAHNe0CWElQtT
gEz8aUrtQek9CwTFWA2182Ck+eL3Ml81gSj8Q+p5mb3Eyy/M6Q9RWyV29Ecx04GM
EmndDDbpvF7CjiUT8kAj572p8CK97DZwdq8/Vv96Ka2WpKqwyYP6u9S0j8L+BrSz
c86c+mVnQm8yM1KEXBWJKVynW2LKLB147TqrLcQ3OfIdAay6TKINli1Uc2mBQQTL
ltaD+97rovs4oC0nvizJo6egaa9biMzF3+ysu/JI++qVBAksHYUVZTqjGYkz92Q7
AVn0dl58XOtrVeVCPgMERuAsARJnl7Xk+hwY85DDRMj48FEY93G0Cti7QaFZvCXW
BcnOkoNxBy/FdanMOhxXcg5ElelcXpMD8wCQxJs2Ocb+8t0Pek0Iok0NWbbRxOFl
9nYNwms8oyx2GoXm+CUqMGtbmlDIwgzWdF6GGVbVNxER3AU2ZE0IfAnnc40Gws+W
1O7YIAdDXy+PzXQh+/LBG2wGX1uw2GFywbHCgq8fXfANXz4OTix/EUGuP7U5n/yw
9AR5HqNajJREjvT7ewmhI5sOyPO3cy3djKJyWHf3A07ydMb8Y0mYdCcq86OmyK0Z
uJQjYG9WxxRENUynk4q4F4AbLptey8LK9FQe8QrhE6gr2gJtmUmOJNosDThAHo7d
4aZZcB34MqG/9223+tFJBNxnZFN14XlRyaZBkNxuKSu9ePI1kKDU1zXN2r111zCP
D2akysQ/CQnY3Fqm+gIXsLw7YlrkOfsfl4gRqCAJbo1k0ueAR2ILSFOyBKZI2Iw9
i4+Zq+gNJd2uo1AupaZcuYLGavIajTnYI4p39wh7bZlMyrenj5AOU4Ytqw36ju+l
DYn9gsZEQykc/a1/RURQ24VX33R/4SvH3l3qamUS35H19TCjCMS5cOEGHF6g3PEj
1IsbDTkHF/vk4NIPv+J6Ud5QU3dUbfBLjo8GwC9agD3VIZJ8ntRz9+8ih4GKrEOI
EieJHc6ueNtUNaFUDToz6bTIOffzg/7lCfSyQyei+vnCJ26H6tiVYv6DhWv2Hbya
WdwdxcjtqsNx1h6B/ozEp/b4sd9kC+Ro052/jkSesJ4EnGLT5Gtaky9QCbdCHxy5
gvL8YUqjCedPp5YcCAf6yKF3S8KHjXQ5FXxlJc+/rn3ZQF/T759V/4fXqOSI5b1s
Lhlw6yWqD7FnatdSRPs8tZJ57sMJpDtV7651k7Mrv40r7b8EVTIlRum/P11KaR3N
EbC6o+XTkvnnQRgpKRXBxDhQnVHRjvJbhsVqRqOjHJY6BxlOKwanVpGmxumJhpxN
9BqPH1ovGN2VqShkM1f40B7zxb4i2nWlUBeTIwnXDjtUJIWocJfHZ2IdoZxMtWoi
SiFV8vQfveYPOxWKyFm025fH5LZ3l71ydxDsksAeq0NfBq2vJMlLlNu2jRrfHc2Z
WG9a/omBEMkjwIlc4vJ9xlE5MAKqPotbLoGlf5vh4uTSrb4MDUSisucLaNtsp3Bk
N/M28jqW7McA5YNUSJ97G0hSmvGUFIS9Erv7TeKdoHMrR0ulxblQm9yibK/vMIY7
v5nw584jpLGq74j50XR6YdYeD6pdMEpsQazPCvDBpHnYVRVwHFAsLq9XcWZUDDGQ
v4CB9DSDu9NLND2zH0g6zKYF23poB66LA+JGmTPtbsoFpNITerVF366fX+8bmqH8
YQnM/+OHmZY/wPG6rWNoRavnHnqrtXGdt7Uc2rjpYYkxbxSmadCXkMg6wnK0P/2A
7WausMz+KO0WmJAaPpdG89h/R1RRrDXuyHQ9xkB5cq7EAgIwaa1Yx7Hp6WjwncLd
pl/EiZafnFZ3o48BQifnhOChNINWsHQhCQ2tCpq0NfK5ZraMEPQ2VfpfABbmJXDK
VMQqUp8aIJvRPE3i633FHxOOV24ZDdigHzBasAZEISihkBHQix9X25InuwwKlcmS
XIkvUHtQZPnBL3EoG15BsGw6CCYxD/5YEvLX61l8J/b1p5+Buk62EbgZrr5zfZoi
Fu5q37wrpnp3ExanGK3S56m3MdY9TOhakL4z8w38vlaBvdl4+D1KQOqDyHrQDYwa
B8O7L4nEpbQicFqYueDXZh5iDhNNYw4nYFk8F2gnsLJYTh/PKKfGAKtvlu64zOZ7
1KO6C9naJwqpPdVm0tvlpDR6G85HaH16Unrp5zMvTK1njedxrb0fJC78nad2V3sd
DtJv793SD17wYytraMNgSwqkJQRBWqNVV3t8XC2yMHZWW/nVWd6pyUkOmgiPPkgQ
ofsd7Br3tPYnp7LUlfaxa7UgkKcUfEiIy8w/uILW4QFvdb3dMTKmq7DE9e4tlNnN
gkMpBoTAh2dywhybP+Ontc3Do3DhEig6/ylYs/+d33Gd9hPtraAtY+5RJWWAPMzQ
yfyieOPiwL0MWWLVEtNBf47E9ks40gP53Ybq0sJ58IUH+dLZlKSxgIf/iiR5rCWA
8cUG+7d50AKwPTRsD2vjVgenM5r6cY3Oa0UCYga9ghTuLCuOUJZ3wiIvnazg2Csr
ZSj9kYKjPYBmE+mJLaMysMrvZc9mSbQ+dh1oktqEAZXjoXznLpDycxohpEddDX9m
oPT8W3HPLELQQtfn3tIFj4EFDYC0HibJj35Q6NbpZ9/5AgrAsl1dkYJGj0jhOtQe
n/Wk/Rq8dKISEh7xPjr9A+HtMQweIbbrXGCulKGnJb9CD22sBd7/QQoe+yF1+Drn
E/89rouKJK4p/5RH3aV2hMB0ChKvlyL3RqnhQMEQgBfT5MZYcmM9vTPVM8QilwL3
8fsF27LANouEq+0EFGe1fAEF9vbV0rRz/QAj/vDKZ1GU1ceH35LthkkxoJjxM7tG
vOZPGuaPzDOvoUZaOeMmlFJBIn6a6qxVpGUFWPLEQU2/9PD0FTZvQDNVU5qzmruC
eZk/3niu553s8alML3LsVT+jLnQh5NT9USXL2J7sk381O0ZEwj2rrqryPCswNO07
LkoMv++ePVZVdXAkozuy7PVtU0Gl+6wSDJ8/XV0qJLdWP7ANqJeSVTAbFuaLi85V
ToDBJ5vR7x9jiUbmT1mgkxqWEunenqHo4u8Mdp/JyjAWc/Sa+kHZNUksvqcEnPJi
+Z2IwujMovknrF8ezdOqNHgXXAVys4wV5VOhqZOnHbQR+yurxsTgcrKtgfj2dIoZ
uAr5m7JWKoGXIStl+KDNCRmTGfbPwNSE7Svscpg3f7rsr7nH3LlP+I9Zg6A0wSZQ
wovnyXRg9f1VdRgkIWfu+kNT8Drv/APLOoyP9RdRjUtrXxoTU4SVtUCqeFXATuLT
AR1RhBsVPu6W5sGJ2U8MZFEqfA0rJK7QRIGlqXpCVxfIZ52dGpOVDSu6Y9x9Gx6r
xwoC4su2dYpTZdS/kYeU50mPjSkE9Pw50Uiw9chkmubmApNuy6eGlVF2fvleur6k
kuwVcdFQwNZBOZudK/OGay0E20zTmI5HhEtvQWUNb33TgcygROizeqK/9mxcwz5l
Mq7J4PfE+Tk1002wqU1CjR5CNEfPChBXRcW87W0T+rFZSK8EDiYZE7R4Br1iLFoS
Um/tsS5FR1s4jKAE6RimiJc1bAy1I6m362BkYmuaTNd5MBDX3yLCdftk/nuWnC5E
dX7i0l7dmJ56kKJIKg0fun1CDJw4F18SdR+ZNs3SJrbz7hJM9OxME13iKNjMen/R
RCw8112ybzxzkI8BTyR+60jGE1ePhZo68biOlnF2lNg42aVJCIpkKx/7DoPLSVev
2rq3ykodo+PQ5CzxwHq59WjShDjrQkDu6fGOSCFNfMxLrIJYIldLAXz8oKA4mOWR
ksIHnYDuRM64sU5xv9tYAiz/PXKgbQefKCKbVjm8l+zyEhehvBQSBdy6nJMv+xUh
jqEpPuSVMWmKInOemQuZ5VdAmJ9ZXlpFsFbhWAGd+d2x2zcCcObWpkm/SG8ihXwX
SRHKRtAO6vrCMBH9UXEcThG7ToCcUR5FfChECstLbJBI3piBfwf5gzT5Pu4e6VMo
PrFEPyfVHZ8YKeGykBVdJ/kT/o9jjilzRTXWBGF1Sj4P13KPI3P77i10plBG2lHI
AM1XWHAllCPSM8hW+Z2evjEWGThaNitZy37bRL5vw0/PSSrsl7H7m/k8iXhT/ULa
Z9daHy/AzVtjk5hbJz0FufCSdtuSHYjjlwwNgZeqwU9csOoMVtehtI4Eeg6gMl8f
D6cCsRBIyvDafmVJOhxMkKXbgRvu9jsyLWxSdCmcwxtCgwWWEnmM+/LGEyhLklJe
+wmSRt1wanuK85iGVKN6OZHyd65J7ahePkhvrpH/c7zew6XjixP05qZ1UxhIVvoE
3QQtGG5fjju8GgA1kxioMvheEiFRYAhU6BQVfixzVfUCMrE1EHQRBIhdTb0dz7eP
jtqSqEkpM+JkPtLG5golKnXhdJ4my0hawa4g6nYc04iivWhEkTdrMR+YVVdzUu3B
0oX6DuuElOs4+nrq72KpODIDY4muPbcdTm5rC1EqcnjZG50RVlBgP4pYJso79VH0
g1r1uypu7cCtWv4IozRl2uUU1YW1Zayw0WELmlT3MoHGqAGqGv0x/xBYvR452eIr
9E+nf84cmMFLsEiJzqFSyogc4kbJAhS7734osKA71qHhFBo1xYxnq6qBwLu7Nyio
42fq4lthRrOny+Am0Wu6M7zM+MeibYI3i+jTIrGdBoTW0M1IIDTHigTRfktxISkt
3E1rrxqaFBxBsVdfKtnqfRGoEkmGeAYFm48xPVZIMC6QqyyuXA4lalBm1zbLuw0a
E36PkR9KoFJ4ast8NWO/oQ84D3RaG74kS2T5NCQQJ2iXNwMAYkOArIgelA9qEspJ
4cATxJFUz7hA4Fg0JMVfReFKDaisYmA90yT70TKKs9mj3ykWGo6vAy9tmqcBlNRm
mz2DHrD2+PC2/OwLm2mt14/uPziDk11//nDeHIx80GKFWk1oHoAKqXfCLwuytpvh
kl/Qz5Xk2r8q6ShIYP/s7hZE5P+Txuv0lDFv19hK1deeZNpQ/0yHR//GpX3tAnBl
lBzVm2BbhPqHT3HujitF95xd5Hk7ZjjMdeKOanDyv+7YVAfJLZ66smX6NJCTZhyl
rbjx67Ppclw2QLOohMd/vcO/jA7lKq9Mg6/Bp53xyz4f9nRFU5eiOHw+RLpjkdtk
kQDkm+515LbYfyAY+nYghao04/VEh5myqk86PNttZJKQTSyj+J+tTLK8EvmON54R
QTdNIzv5LPu964Vk2yUA84728R0Hv5b+tKu1A8i7nwJ5rGhIL19UWlEUaW3ZZBeY
+s42jKQDYskAV+I0tO88+2x1O+0l3RtIHYptnVbyren76VRoEJ8b02AirsNU6JQS
tkqJetGd5sEB3CttKDPL/ltorgV/VmesQLLuvLDJ+jUlaR8lToWY87JP50zto1Vr
qAZ9Av32uXvS9D0ITEdTFOtheRqyVvmvSnmcWIM7C4pSZQXJACjtUVGilDb9O2jo
sVsbSknsLE30FekHuIwsw+5nnunx1cUp324OMd/3pGGT8b+X5ZIUUgeBlaZ4/Hr+
0aIMNgGSWRz0IMIng4wGdtiaUPOtHsq13KjcP5aRPajpXAYg0cOayIQQZAXykHEE
3F8zk2OWcW/AvXtr523DesbGGBiRnKvjOJvb60Xe68BDzqN5LPuVuINnXXOJP3iI
e7nroWuBvl6fEYmYKwj1zBx5l934V9brVuzV44XotPSuKolmsXO+IfL8pgQmMRtT
5qxhdFctWt+pHRPpj9528WxYSMgevmsCkn6gSDSMngjziS/g6uMPxEDgFQm5SXzj
7NhuJoUagBd9Wy4kXHnSKChG6yXNufws6tV9GtnZRTyzY4T5C1GmGerryRUBqNuJ
9wee5JMDbGU9qCd517pFF+n7WBW/C1Yh9o8eaIY7BhJfthWdcZRkNQHdzdEnyejs
6RuoGFBqUDnN43w35/jGr0e4Tgy9gttgguUmUIEzhIN0pHbJNkpm/DXsU20PcSpw
nS5IrflmPZHocWyY43cXoGXIXxUR+EKylb1/tAZNW/txfnK+pW6CcEFZuJokxjBV
bLTb5dIkVYhpP2sd53fsD3FmMp2mAuMvjCHuWNctPyJ04go+YFrdM4kkvL3pPPYR
IGPMNi1bfYQcjXWq9jYQumWG5UQCRuMtoc62jxX7hx+J5gtTv/dlO+7B/dg9QvUq
vKkiRv3jCQRVbtm0Hialw187w7izEts4PLOgeZSUQ4yCxy9eDtDHUWx/q596iivB
Tz4HfR387849yXghhHXGptQOILVX/AxfRcSDR8PcqurEIN8/4kutn9a/Mdqz6BxA
/MXdV9jJXj6P3kiZm6EIUGraTDOY5ZwdshOQUvUuLPEfX823nkf3GC/1f6nJCaIV
QGxWRT1nv7TTXW8MoWpfHGP7ROk9hI45GTC9friblB4Xfq8cZZS0nYbXCVEhXTbt
f4q/5fFTcm6OSa+zDM1kIZmpT0urq8JRhN1HR8q1ghkciU28ipP5VOV35KF3s9H2
T6AvAL7oF2y8+JbAGEKlX+i7YDMKzs+kthUwV3ijocuPOxPWP+574V6LRvT7+xxz
rqkBXonkajMGa31r9VZZQ0EnD3OijM7Alp9ehZ2DHTeB2nNSmzFrvpYI7qjmG1sx
tMIWRyLIK/37dcBSiVbn/ut7F2IQWLDn5uEBDyF14usUCioQzzSPoW24CZ5pO4Co
yt0hJYUQ0aS21UJdBJ7yYSYtOE66efkhQIeeaJssTXvOYgIfl+TfB1M+0WxJTW9o
SuNNZhN431S/MXJNUlkcuUB4HHkFQE74nb6wJPicwfgG5USsOVpC3D4BkblCswp+
0xNPvi+vv3nzeL+f71sdEG7VKnmEO8NmT7vSfGPOblK55tHreG1dlOK+GWOO5sy7
rbPhiD65pWcask4W2OM1ju0+negqDeoW1hNMDDe9reSeJl+49Ek5hJV2dCkV6kxr
aXtMQOFu0ZuZsDyzbPDTwSGzBNjmOIgJICvV06lzr1/4bTrwc4R0XUlsXV1UhF1w
zSsJfovSb9IxCfWCvk5QOpojN8ti0g/aY7UdPiCBBm/KItAnS/7A+KFCbERKVCp6
RPOUn3UQzfkUWiDd00lxM4feeJ3YCVqXX4m7t4JuZByaxEwxv7Mtq6MvAf9UB2+L
OQArJV5V3nimclcVQ8zEYMCKgMxfSB0Io4YMRbJU9f2JEuMXK8QBdmtvYhEa8vBj
3PR0rGa4qLjPC3t3y5+ISO+rjnFY2lo9mCSAF4dBU241EFgy4q8dSuA4wKo5zlyq
3KqQ8ZkTUm7c4uY/BUgKuAji8qKTJTU9CTIAAFuSicYEhdI89Q3BYml5RpO6ZlZm
0WWuCGcjAGgmaJ4/1uMFWu/UI7zXzBzq/Zw5rQk+JgYpmrTB82XU8KVRLn5C6Yo9
cttTKk4d9mIkVM2EdJJNwzEvShL9cuIfe7LzXbhkQs4TqOXmuzTAvlewAW1G8dYk
RJrNEwpE5Yqz9XBsf7X+diLY5SxkfTAT31zbqepHbtAbrBRKx8uASIKeJmdNhKqw
oLf7h7VKMrMj4y7CWmgMJOMRfMx8F5uULz7ytNhaulyEsXqXnMdAidp5wW74QZE6
+Z9XU2Zstr0hk+eMAPxpAgY1XRZP6qUJ4FpDD4aU4AOPRGhF45poSyAfWVuJlJPs
G2qAFdAep78CIxWh15JtQzfuawfTYLmFBJXzp2kpuDwuh6k3a3XQFX3KuoX0TJaK
La3vJuRmLwp3WoOlpQnVj5ILdFVNymSE81fF8zjCMdYmSChCOKVKu5dLv+woW2UR
naVrtM6qEbhdN6R/QiX6Mtkt5c8RFtzSrEG29loC7Nccb4NsxdDB70SxW/OGHJ1E
cb6Gsi9oPstsc7pAaRVjBfzN+nvjNWPMA+ElChG7Tn+1QUFFrI2rZU0P0S94WwKR
bCJRQCi6+sKut60R3zjqhHBWJjIVVL4z1p6s1yGty0tTbJXFtQoCebq/q0VFV1PK
n+8tZ2GzMXUczBGXadCC9GGPzdASJqYfgy1N1bRaON4FAYkxlGLNsmKl9Y31iEo0
JkBe2+MNwrMFfJqnNHHUGYzT/tYgfgDrIO5bbdw1jplaSZBDp7kvVvjoEXJHgAse
fNysrF5jrV7gVtDcfo8mVoRqL7bJMRoXT5OIVnGQryyKL4wEPSm27wqP9fhcVCFo
mR9PBlDqNd7X3QvdhWWu1qP1JsKbc4iYDFqys6UMm5Ok6T6pVf+7tmoSR4buaOK5
/5HKQTFqqC4Pcp8r0CZuR8YL9+vArz5snku58+cRmoBkm9gUAszJIKNoGiBXvpbK
08wppkowAj4ws4pWJL8FI+f9yR2zIAtHMFBV9LrBBlo8aTNBFvg6CIPyjamC7fnl
DFVZVfgfSYRDm7Ds0qrADzFGxW5kXAOhyJ+KmAAoPi8RdRkCLAB0Z0Cc7yMSaN3c
HarcOWMUyyUeystjO+wkRavsHiCwHTNW1a7wODLeyTImI4hHajghmMdNC9C3N1wZ
H6c0pkoIY7WHqqEtGU3gPf5pHSEw2hVcD6+NxFQSYt5PARVrbWrz3WbpjYlxR347
wf4Otb4OElX7apGvZoVN1c0C9QyUFV1i+mObvWNwH2O+tgIVB6ce9zo6YpWoO42l
zKo8hvXc68zoX3fosUIzziHn4/mzNfvFFeQqTP+zUONm4etLeIOSzS5ZEdi+dOL8
88xUtzlPOKF++o1VQ5XqDzNS3UF1pc59lWAO0wg1uRd8t7scfUxtlU23vKVyQ2vj
8r5CAPUYSrPTfJ6NmVEGdTIFdebtz8w9O2h8+ia71MmFyiGNdpgz27sLRhlsX8gf
mSvmaryCAKEXWZIY6Mmcm9O7ephRKCKrwnJo55x1KTf/3c4LRzM0AJYP1VKbkEVf
+KS+xS/L1a8xzzOO4bcQCG0GWpKEKmVpMrgMNzRNPe0cTdgmpVmWbDzK70m88bxT
dHuDdL+K//MQmJmFiJrrrLv333QqD870OeJELxB1HO25mtSHVJz0xqroUm6sq/OJ
Vy03bCUmIrvNrLxMKg9P1j2LABhKDW0VKz7ZuESJ2nHyAAKWyAYGnAjG59hmqrpJ
VIyYI9W/sQcK8Dtsv2smkp3oiWhosIhldtFr+XRx9djnJPViz/hKw9oRy0h+bfm1
H/SwsMlDr4KY68rLeyWbUB1aJed5cNBHeO3WOxebeDPjazgCl7725wfwnStnyjg3
vgHXZi/t9WDGVNn9AOVKK5fTE85m6pYs3sWaK72MjbUkAHjvTDW4WNXe7l/zG3ae
+fMitTDKsWYVA3StCa6HpYyxbDnUIrV6EJCeocHE2in5k/R4bFz/L2sveFnbxner
PoV6UGBlTwQCAq2H/Qr51LwzD6VGK1t37Q4eNtLbGopJdmIK0t7hkJG7ONGOa704
9iJJ7VQGCq+xi5j+L2V1Z/WuQ/HmEVwAd4sd/o9htfcijzM8O2sLNqJ4VABPzlrg
XBdfLUA6zXgZKh+zkwhtwPfV3DfLSKi7lOU5siSZM0n8DbLa9jgS7SfhOToisfrI
uOo3cD9oUGdnSzo/j1Ved0SFgJYp7pdprdNjsZvXjHrzcVg1Qun8E6PDtls9MLCm
1Na6lq0d4OvmLNZKWPD0ZyB+AYWgYHrMmRYn+lzuiK8tESZtlHaz12JsNe450s32
GPi9sOSwXzWXrWWuCpLJFdZKyxa0fTrVWmLwPLZU0tnb82JceSQpQO4EvNrB17IB
dPmlDvVN2drsoM0Fm0fmzWY2dcH2RS+trLfKzxyAPPtQbSUhIpOb292lkJdZet2e
v8hQEs0bdWxG3TcE22xcSBRNOHM8Nyfw3h0kHze+uvzT+kfiiCzY16uyWfaSzyZO
J39txqx0Bh4WlkmVsrGm81I4QgeopzprKEii7g92AuN4Tb9EwgTRiKBssjw4GmJN
x0xpsoj0pi3YyvaXCN46nuartRqdb8qmi5v9HaZEFWzSCEUMgRVUPN5lrqr2inWR
mzKb/ivoPqgVyJGJv87UiC2nz2W+GTdEMVDpE165vwtQVhm7zfQ57kRDEyhXr65z
eOcnpz4XbyRTDO+Srf+EOU/ZTZki2zRGHtvNNFrHLspk/3asjMG5bMK9ZdZFroIQ
kRG5uwM7lMZbSeqkLQGPktz8+LhQ3VBrlJXgOfDad9CHmQejmUNeP0M+m427eCsS
m4atqpKAnM7y03LoxkyN7PJHVSe4Q3YKA35Lmve//2EvcAhtReEfCVZYdebVPSgt
CcOj/JhIMhRvoGbGe3qVWQussTsrBq4hxkDm32eu9CR6Xc5b5KXX38hANRbQvLt7
CYDR+TyLzUxZL700PfwSDHecqseYC6L/QY5/fCjGVodugcuZvOnu05qxYkll6tuc
4QrKl0U+P+WdfEV3Xt8kMJ+wouFnf9aij4afciYjTOyJFELgNwQKzWgAFS2SN1fA
2b1D8LPNaGltSJFs6P/XkhoOoONH/aXfFOLYE+bnHw9kwLmgPyPNeGQlrktuA/eu
4hZkBfDzmmfyHqoWDTkRat7g3C7NsVkuW2RrQZmfW86iwodSCQvXxqAaYLnbQTiM
u9HFNlw0u6YfDVq5EjkW3VV8Te4lBUowyOzPIDwj8aSHz37glFHXei8eZcQBD/sb
IuEsMs0m+NED9zt+NJHgZISSQah1SplETzXyN2KQXpE3FIbJhT0qcJLgDLVwFysX
7bz+glKBUPwzXibAkWXof7qB0OtEHQHZzCkVfEhDKPib+xvI5qbYDfiuTZZYCqrI
kml9zTcaHkj7UJH/YxIppbuaRNIhwTJVKaQfXHiuGNfVWMrMlArjnyU5XLhBC9mA
av+pEi/SJgeoT29UXD6kdf6bJpHsehDGITlcNDIT/QaNd2z3fqGYAMV15VP7/MfJ
+vdLL1MoYyl1AMhypZ7rep8tGXCEVaWUyfsfv+waAL/15w2I91d5fPQsfIEMYmtL
J/jGnwjSY8Jaj0GvJlIW9kvDvsM72HgIIDbuheaWD+WoHZof/h9PpAe0WFkJBUQ9
D+V/4hO9lCAX77SIhp3sDxyqL6sodi+g05J1S9GgOCxzJ3lwwau7D2uZjXrXcWo5
ftgm2FuyHu9w5t4aQwm/nWxQc3D2DzE9+EXW37r19wBUXGsk1Oaiy02t3wt4r5Ga
PlyLr5hH7xajaxDi45wHv/2dxX9RcRjAxwbX1MDfX3o94GI8Qc5E5PWlEKkrdbQW
OquSpqrzwGorX4EUgwOSr4hBeZwJRpgkIcuPetMKJ5oXkugNgswCb++q3QLHCMh6
fuTyAC8ylqg1fqNGdh8wX6PIKo582TeUBFTZX1rpNO11LRxsbktDOFbl1iU6LuQE
X2dXMD4A1OaUwb2zye4CaZ0zVIK42jMxSXfCMqvEk7ddHpF+fn1WDs23vQ12LMp3
vktCU86zNjPCDec2fL6cy+gDP9AcBt2lQQZoIxfwK8GLcymlWjselaCE9I+pu1h3
wkuSTYgwKwFRk4rmPZ5ZUDZr6V/OrkwLIGInkPc1qitD62DFc0uGROIcYct5thEC
eD4zeXvURSKkyEaAeoJqxywdgYRKeQGePNq/x+0FIuqIto4MLkYjCIcCHsWIWrzF
EIOitARB++/CCLe9GWvtOxq1RpL5umeVjClMH7GZsbmpucSeC3S572fVnTLDKsC8
4iJ0edc2tkRGY3VoNy2Vqf2fi/g+SeJ1U6Pemc9T+HaXjHH5TmbdzA78udfx8mQ9
sgV+jNa7woleKsyg+liRpggrm5nJB1DbeLbRhgEJ9gVUiR6F3O+0+vC/Gdq6ZzMT
FM9rtnp40JAN1cyIRh9QfQng6qIHbR+iUxhjdhQxzRGb/ASQ1joND8KKdq+ZoWIn
/SXFhgk/X5vhwLNrRuCstiD9S06WLdw3OP6EXBc1OSZuu42xc1HxILpLtaXxWp9L
08Ij9A9Df5Y9Uvv7gvUteaCZOcQ7OWsRZj/DEm6G3TPkRwvtvwOIivG1U9Y6trf6
Yi+slh0riDXwn7g3doaq1pDOCBp90OQPZyvtCfDwPcEWrPa/P9sDLezjfp2535jJ
UnJ0NRAKyk530Iw6vOu0T/xW00UGTvxvrwT8F196QZg49jMa85bgbNza4lV2jy7M
tHBi0hRK5wjVha6+BhZGbi2fkzkdkP3/F+V4neBdCB6CwJEpD7sIWReP5jK4RWRu
2CdcZNXuq7mziGOm+iJY229hXQpinzWcaHC8oWAy9odWdbLYp8dg/YzHend2fpQA
ZVPD8Uclnfr1SCY/7FD6sY2SbvzJe9LXL7x5QFBnpZ8KKSl3VTM2G8ry3qwY1xzf
MN8QXjHXMwQJ40Th9LzkDxGBB2UywYqi6dqEI/SQHOrGptHod/3KK7orJBlQrbws
gfuidwhTMh5fAEe2oM6NYiSJqhEiqeUe1qKU9qwYmRxSVQITyl/sAOAbP6ZNnuYG
YGYGBM+JzMw55rslEQ7sqedZxRh0Rqw5Ax4f290GMqchfXiylS8FvFQYfZKIoM8w
dbfQmCHZUMJW5u7kpX1Z6nvc+jAtJb8w1y3noQGvOL+Xtumnv+A4phA2Ulu/1Xji
5qYmFM6/quoJJHKkJ5IJP5yjYDRs7iMhNUaC/jE2UYGWr10VoLAU9DK53oiFL1Y9
9/iPcIl9+L9UYq1tnlRJM3k/98M2XTwTYMk85X+JqtCk3fUJktmKDXKCqKpQd/hg
sx/pw7F7i2mdcic78s0rrqPy+An0GQKidh3xRGEdoaf5/AwQdsgdZ953r0evhvQh
/+84Bz2n+4EADcxO2HZfDR8mO3jpyybUH/f0pjOaGMQnWG6+MnwXtX+SqaAfsE//
yDKVABopebnZFz2o7SaflTJc4zjZDO5X/2xdyDIqYdJBXEtSZzOdlAmOXQcDd+Cw
dAo/jzNcci7dSJkvSuddCo6zKi7JjCfKCVvGEQJK7Q3XE3bVYCU/iGy65BjtmMb+
57806/cp3kpfoYp7kxca27TKjuqXLH/wAGsvLTMpgEc5CFrjuQ9iMEzCqPj4x0/O
K7WFzeV3W2YcJNwIacJmGkQgnOJOj1IO+tsanMtxIHGwZRquxJxULFtEMROMjEex
9weclWMpQNRGnKWG4aYr3xOCFvFy5wK9hBa8Q1OyZvdntmtyQ2VZfEqb7Gr+gceY
1EUEi83W69/qSsKOd6A7i1zFtfyrf00h+vQ6aZCvVADh5onSIp4itbpWLwbIpvLE
2oGBHxIKU0SmNE2AeXrk2KD7gUl+sES316wp6P3YRp/3Gs2l134r6oIY+HpR0LIn
DhnTYRn9+AetjT9jBomrctVOsb7sBp1gprT/7S6loqaES/KSDkoaRdtrt4rRE6Sp
NFL3z+gceTI+kEnlBJEeRo3ymZFeMHQjCOIYJdOlAYQJcjF4ayuZcAH1jo6YRht3
5CRgUJ8c3C5t3ASw2loA0pksVl5lFXW9dVensCufFCrCPFNZsxSvzs2TtFhwgWfC
yocIDMbL+wbv/Yj9HUt9xMVLMDqx6j9Ka/VLcIBxyAR2gomQxqOfy5tLNAbXGHwK
UEyAoaXoCoJcyeJJhJ+5raREKPf2YkgllGAaNDL9d11MBzNV3gK2fgDPcGxA1hoZ
3Z6KgTqZi2Jx4BoWxKWrxu1C5CIb8aisBSjKgZX5UzO7eV4Ri8djmXri4SZDDIE/
QrIz8rLSzFHajQwBbSZL02NLUFxDQlVbDhaxsKWvx9yKque77GinnrYWsRgNfL6e
r5iq+or0TTnZnYMlat6AgTi4GIEQk6215dGHDXwvnl+bhRTwB+4l9U66F2Xnwjf1
4IwGfbu/Sl5grenu4O/sd8qHPrJpZ9Gab+kjJLzVjLir2UZWZ5c7RbmH4ubp0UDA
ng8RNi8SdmwQKop29u7ALsvGOMkpX5cEP61u9nMnhX6pKvVRl7Bk448oVEioSmDv
AtsmSB/47wYRB/HI/4VYIKLW1fOT465YaBUgUGKcY2TQeaI0htrprZNP90g2udtm
3WxgcZxRG5sFJF9SiahIuAWR34txGlzgxp0PRZxFFj8F8E3dFgx99U8vCdGn8iEH
JzD56OWu3CQmOu78cDuE6wB3OBmuqRrQSx3ptSm5/BiN64qDSeH3VCpEzbrnwbhs
kHegWsAZPO5pW+D5NTX2INVP9ez6IIYKv7mQa8RVFJpJj5HgVCriVj/KBBJZLx/A
xdWol/tQ+zO32K7CEYVDtokk5WgqXVErvEj4QqPrYX8TnXnYbXVAjCYPepdU6rPH
mJ+a6wwaD+Zm1URYoxOeA+adSPKX/4kDatFOd5b7UWVCnw4ZKrheR9OajIiUzf4e
nAvcmsfAtww6X7gCBAUt/E5iG8QYRhCwQiaB+NrajpomlPsNf0Z4l6/vKP2xGan4
IdLz0kDVQEPLvSwzqdshwpssFGjZXU2xUb1nQvjEGvcMDvWl0h/9rKImwWR+A+BD
h6sZbm81mrVfmfFPQep7lIDRxXYZzZaRFXG0eEkIfpeDF371LPp+ZUwXABcR0eD8
//qiLmHn3+aFcvfRX9gU3aFyXTXAStX1k5W6iBYbfSg35arw/IReFNzBFrTUGYUB
pGkZsOzm82QhdpeEmmqNHJAxgd9Q1Y4yuEM0rilfBa9pOrohA9WrEo9cZUor5E33
6oC32U57SOnoqQaaOukorTTVREmxCQrqSavw/mQUP/4kZV/E1jSXt8eMr/btHnzZ
86UJ+AKwQCQfHYtHlXloD3flL7PfYWHdEfZ6x/UBOCadR8xf/ioq4kQkoA5AqmUV
od6dZkWag4B3mGf0duDjyi77Zn15AtHLLnr2BsofdWYCPc48CEwNXLyimynJHlWj
JtfHYQ9fJG4Hx+2c8dstEyfSfiIbC1xI3/DLq40SQtRmsYHhv8U7CoFkkqjlZMpV
rN/9JACvR90NwtcuhcamsZVkUMjbVLYY3CGb4qHhNFDGZj0tKN8CsyqEv5zvug1d
gIjylrjCXTEj6qtpyd5J82vQGhcw8ZpZz9PoZf/yBHmPh6lgNNmUrkH0XmFGrB67
lI8k9Fcs7Hqjr9EbGra5UCFGT+c4VXkP5QeDHGGvASvIrGBONDHD1k/PgoW0LPHy
kI+fl0k3sEgnqb7Y0gSN4FNl1XjwZwsIZj37zEdwdi58jWyu8qyq7IPiBkvlxYv4
KscYSbCv1RsRDm8p+48LXX934rnpRPvUqGVhilzCi/mPR5k26jy0KTS1vbLkEZ5i
mkNz7MPVaWtjXf39DM6J6zgaauytduwUnfpnWNTIZ2OWoKsWlZVPeewc6p1JBEL+
QecyAbEasCvS2qKef5i2HOwqCeLY8VDxwTn+86uH2IdDPbe+HObPJ7572OPyGLeQ
mt3+ty6DA/pdhTESr5W8dbjXk9/XvJ/qnBxFgHTfbsU2dq2/VVpDAIRj6inb/AUW
R9JGqJ4PPrNgwDysupGr2JLlFqdzD21cuWJrEo1y3YRawQ4kCjHJnU+yKdua1O3C
24DRHKTJXKyTM/1mQj+n6KYkrpLlwm+3lv6Z+2WXr6gxsoCNYUYJG8j8fQALo5M5
sl5stMrGyN7u5hIJwE7xkx4s07AnievD20w4uZ2Z29idQwkS3juiG3/EJDnhsw6t
n41A9I8ZcVqV2eJrgiM4JWZl647Oaq7ZsZEj+WerkNd24hasXCYUhTvxo/kTdf+D
lS6IvFVhWTOf6+0Mg12vCBYm2DDRcjKzXk01ZtoqJtOmoJIr8lCGK7Goj6SFF4Ip
WDOIdr8kElVmjnirkuF4TuvAzeH7PIsEF0Fo/gm+k9yvlYclxha+4ekDyktmdQEO
Z3TiCW8NsGlM/ksfwJBlRmiOLVuG7ff5W0hZ5ggBkp+Q9DCP6tqKr2ItNoOfubyt
Rjy6K5b3eSoX1cBW6xYF3XHXsoL4kqdZbzn/DfdImlI6XCPFhoP0ZvA2QcpBofWu
e7BWSMYrHFIMfmjOmMaqb3gR1+9e+Pyo5NmGfoBY3TKmApiyI2MnDqegE+DxHhcQ
pWqaXg/kaWBoVjI6JeW6cBz4ckyDngmsPYNAGmP266rRXnsfFHbQHrROVhohjMWH
UpQ4xeQ9MaS7RBpmPnbVRumjKnfafUXbD2MUvRHLcAnPnC+0ntVoRDLUXxQp+wk9
OuvAYwgbKHWwfgGzt2jQVhVKiWMMEQv/u4qLHwUX0hz9xAnB93/J7pM183S676lF
AZtXmb7/+opNxx1Yl9hJjGMI662Dd3qcRzlrXV6D09e/MNGCQCdXXNuMvDRDx47Q
d9VA2CA16wqZOAI3vxwjj/h5WuBnbvHbDPPSqtsC+eVzK6blwatHQyDCsNZmwVtS
UkFsLd/akl68Yjtm4yg80nCe0DeqMwk27MHGbr9Hn57rV3EnL1f8k8SvTDq5N84d
Kf/o59EWrS+7/doMT9SWi1GLEUXdUioWke23sSGAqunQBrMztipK1yhySD2k1tDd
2ptVQLsvTsn3v0iyT/dA6dq1A/6xu3HqfQhhQhbAKBNfcxnFwY7bwkNvvtuUYUPe
im9PShGqzZJ+W81VFndz02KG0xqM2bN9TtE7PCdM4DHh64YSpdotH4URfJXLQJNz
Vlx50PFjxUc1k5SND2nJnjVFsd0flDOyR7KzwbHRxjsItf0nvp2gvPMvECnX6gPU
NOZwYFL746yWCVBd7Hl9dg9p7GvPfRcn4zJ5bom9bwp9AuCJnTDJ5hozuuCABc/v
7VQNIqT2/XJbaOTVAhCQ5y7Azb0AMzJ+oLEVGU1c4zGH3D13uLcNzt4KgYLh0xYj
rVUNUgrXCUJUldKPT3I+UFq+TFdA9OBvMdtKpOd0P/h5EUQ70IAAwotZqwJS+Lkz
IvcXe4WrTmjwsIJF2sA3InILWsVXGTdlHUSC6ZrF0xzb2cUGSmlaysiyzHN1SM+1
N0ar3ZY4TRU1AH1Pb+k0h2HH9HUM2YohAu0VOkek0EswNTUY6ZyF31rpislvyifF
0w+ULEixnJ+EstDlPGzeKuuFhGZgwKbcsdsikMU1wiV/VHLpEu4NI4I8RtlKPXtM
Skew1+/uRtdUE1IGjg+QXXGYEMrQZBSFQwdtvLB5FFCsrs+q8zAoHQ9N+2gHV3Hx
C6w23SCkT4QM8li9Xm8xbxc5jPi25iG9JCnpV/67JG2yO92AC295qP/T+VWYhT4e
QxwTkoh1EDEGc9iFgWCFeGXOmfGj6CnfuBbIk7hNi2X+8Uwp6DzEbJF+vTYCwBOv
exE91xfJnwmrBKWL7HTFxVq59NmZXBGZ8Xo6iVluhrwZDrdsoNHq3aLAF60EdzkT
l3USFv+njo8QR9pO0pbNwDgN96a8wAcpmfsd7aFNEM0+jK5WZQv7/H1DMZs9/FdJ
aVIyFnKifNSVYZlftmP0vFMxcXMo/HWJJzWr4dZ5g3YfBM7pC1OBIKrUUqp6kD/E
/LW8L47eDh3pvxNw0n+350JYJNnBTlY7Y/sdw5DIcD9C8yhw0YovfnrFZQ4ExcLm
9ydHrPUvWO/dXfrlJCbt3EJWqzknasCWSrWiawxyBpaFUJVZ4fEdFYTDN+GR3Avh
dECfwVruy9/rLF4s+M/4dIlhNvwLz3gzHuuf8rd/1nD/EeK/iSA5xxRVyYJ9D81n
LnTLzmcbj4b9VAhitW9e8U/q77/Q5CjXhdpJX5ZGPd5JQzHJNS67cnNO6X6MDITq
+XmJzQT7yGKJkWDYq8/JK+N//CazmxQq6dhBBcVyJ2ngM/njkBX9lkxR/9wm5aVR
E6nG4ekiKfWCrRy9On25VK7O2PRnSC7uSCggxG+atVqjXRHDnIBlR1z2l1xVfRge
GVmrNnGt9N+Hv12Fqd9mBHg9fXuRSvyknRmWlfiy75sV3wcm5r5hjS8KWhZ1IPV4
kX8MRBORKqAOcDYz50s581XClOFJXaoKsg+G7eD6s1mODFDs+D+wYOfKRjW/YDpp
OfL2pAdLqriSi+usHsZ317d+7/G8NRV/A/gu8yUtlr4fXFoA8sAsGJS46Uteu1Rb
X6i9e8kUNAsSq/LWAcuQLm0y5TZX1ySulSBgw+8ScXmZ7FaoAi3kth/SuuF6plOl
t3z8W0CSH+6zlegBiNlDKOg6n6Vo4lliknYF8Htcx4FTR1lzTyhA5jm2Knl80L0l
iE1B4z4/u5GrpKgHpGQx9B12VZPXyRc12wwxUKkoPxYcCLqh9aJiK9K2MrHq/rcd
gAXjGzsOIVjZwSYzGJ4WwKWTkk9ksDP3PvISC4u7ofv70cpWHBRVrjxbSha5Xtth
ceMlAYZs28rTqwJcOlwztb0u3KDgIdQg+TFoiIJH1B+bHsDSPBmus/7Xh2KIwnnL
qwyHwL6ap4InjYAAJbncfOkmMo14py3lm8rk+NFUk202CF47hYhDMlv6kma5DoVF
+XTzUhy5elA0AxFU69zuhg7VZjlwHLCIv75OGCkpBoJBJEc7OnUSsaiZFT82H6O7
TyzgOhShQ6mupDcHWu+kTgTCq8Sjn0CDL5Rejn9fQ+PXCu3JUp7dP4RsRZEnrC/s
Fzb0i5w6gCaCozb1YMLV7wq1YkYZJLVkK/+cd+eOReW7DxMQ3vuGZ6gAFzXBx4tf
Jl3+Rs3Qlf/JQvM/Ykk72+uqmCER7WSKhATqjdpFOdyatGh1Uk8g+x0QmgDKN+oT
YM9T8DYARHXaBF2E7lDQmWFR2NGv+r4eCQ6YjX+p1/r9EhLau7vRkZ+1F/286+x0
5d2liU2sS816wzlrBvVxvlHkN6WbCluq38RxjKefRswMiOw1H2bPW0q7uHI9e2cd
8EBovPGDmC3kK34+EiuSY5rBHV7Ad7Aj4U99OVEJqRWcLp1q4NRb5jqPiTZ+xURx
y7rU80+dc467Pgt2ZKDmKFSVvNFhzbQs7JyeK82j6MsaiZxT2Zknbh3C5f1elrYG
laD992EPowswkJ2NCsnRw5kg+GqvKm4+Hd4N6Enk+U16TSevnmGn8h+9GwZ3BFMI
eJWkdvcaNyUPzSEwFkDhbnCO4KfkUcQhnbZ8PG1FQXLaZhE8SnT3TDXEW/NqYNL7
FSCwC6tmWe9QiGZpR5rQo/aLRfwQj0+JyOQywwfNlUWoKvYejofUPdQ2DGexOwQJ
1s5l5ET9wJbgXTGYs4i5Unbh1EdOm3yMV4H1pp6gCM34kOOj3c6ClXCg4XAtANKA
8JA0pt4WEcHxjBpeT+TEP0bjrjPvi+wR+mpEpsphMuc9ZS3Rf7Iqfc9Kbsj4e9Ys
UQvfexj1rSfGFPit6qlw+yVqtOW11wdPH9/kFeNBtHMmjSdCKJyP0vn3OYg96dY2
vmculSiFCroMfD/doDgLqkjn6OSUqMOlf51NdePmDuOGK++u3eAuEl49Nyj6LdAP
BRV/mB+bByrMVqqECOSl7EoJj4TUK+5t4pJ4KRJ2tonShEkACjgWQXCnDwXATz/W
ZklXyvVA/P3op+niao4LsyVv5gT5ilkQzigj734N5AbLTkm+UGFx1tsttJDEK/Xv
Xlossi0XtjJJyOJc4bQO7QWQu7AZ3iFi488PN8cS2hd9sa7xukNAPNnJcnUy+17F
nnl496zoq5td8FppLWghGveSU6TzxFRhufMo/He6tM+ZSuVEAedv6gHP38LiSBuU
w6kJai78Vwks93gikbcqOWr38ocXW/BBq3g6QB7cPp8xRZe6+EICz7c5n79m0598
wLyN0ucWu+HSBxpAzpBLj3qdcwejTq+Nrbm9/qbGqUF+48zPQToCKwkc9csRkT75
h///PzZogvN9+0cPhuSx/p7l1lQuzmr3kQ8lkssFarJCc+5e/3kpyyU0DEQCP5JC
w+7XE2gFapQNSgYStZW6fc2OSw1mKinBPGFf1h3x6fV5FtbGNR2ZwEx0lkyaGNPf
PsKxeieRMKgWOGdBUGXkX3BRGQCnhusxg+B3ESe05XccoZNcBsh1/Cdn1WIbWpX7
GmT58YH+CVnaRo5ML40bc4OV5sevW0W97X4WBDDbJ00bR1IqnDDxXPyj4Em7mvSR
hfycBxm1GlOK/+1zLVhYqFPlsnZsjCVyhvUe3irmK3MMxRDRMWliUxjEwrVZb+S5
1iDSlEmobs1ACOfPzlRMnjAcrzXp/vZ6/NUaHeeedEYGknbBW8gp79a21ssTUJ7k
GnM+o+USbXKNbLJYXtwk9VZw8kBu758b/0Q/J/dME2YSiVBL7zdK6djQGwLDaSlU
enocKwJXy7tlTsgTNi8MA9MqMad+Z1IRRVIm3TN2gzojRSRx4eZRvvjwbLruQqsp
W3jMliz01VQr2SEbDoljZlMBmxBNymzw/IoExceG61IUfSzWyu9DnLBQG3LboBGX
eW0b/QmTkTLEYgGC8tjs15BJIo57YoGhc5Gg03pkZ8W27tWbslJyxcov8Z2G/1XT
yol9hXbwBSGcx1lVWLY/Nqf1GPbbJjBrymOMv14P3ELy43NJVAmccNL2wbIajLHk
U+CVFE0fl4hA0vVKjza1oXc7N5RaWOkTBCw8MreYiw78Ue6GWPXWLdMQ6zp3UDXY
R3ODMX4guBagqf8NroUfGDfTrtwFMJhIKAa1dbCVZvS4vIB4jN8P2nc5zVdmG6f+
RjjxbJldd9nwPipRUy6aVDp/vX4yJTltTRHGg0lHT9iRxNt8YkC2FSSTEBdRyC4H
ny7hSOQw4o1puJiRRO6trv9UUXMghiZZHmYvvDa/D/XH15jYEyuZMbW61E6PdBZN
V4XgWI+WOu6KPb5r9SM67Qc0HJndLiwJ9AKmKJv+LfzMgMBVw7VEfCIJ2/NLVtKQ
6HQbxVBHvwRIFw9ZULCzi80TrXRqaCLoi+5VfyOYkJ/Qw2LLQN0eNu3h0B6htTUm
rFuyzg8kr7FvJlWzxb6m7M49k0PLdE6eNDpHjpXd76qr+Yo3MMfHVB5KHMIYNyyg
LeuO/CzivhVGnFFUP+rYKTDhTraTi8uEzfN2b6z9gwQXWYz6cSD6pq9tg2Jlqs/t
OpsSZ7apcr1AG8PmZeB+rK6iuQA5jIv5O4APO1TYg19aqus4bO5X64XA8jTkoGe4
pDxYY4f3G5raPqpHTOGEbQgxRbyZgQ0PlDLIDYSFI2+FgUeCwRJVeBPlbpxEe/gk
Q+2GXL0KavjzXT8iZJpf4IqfGffDgIEEOspqlnJzMAahm7/YYuFrvhwymwFmFf6l
1KmXer2ZulBOzFeS2hiEEnQ/zvvvsDMvnozihqMIENGWyEzZOwRGZnN8xDhDwzHV
mLRWCrjRKazIR3j29MXRumZ2TqiVjpw6BElXBX5IFeqvB/QZLZWJ7Edo1R20+KTw
zn+9pjS0FKzaiB1nXyfF2Dr51pJg0kzxE3PRtyWYPs5owy0jT0QP9hCH+CdIp9Nr
5fjgEwWbZYnS7rcjK15Rbe2cUE8A7j7SFQBpaJMOk0Yem6cB8772NKrK4VCLwK5u
WtNEUZI/4OL72el9v2aRtnVWbzfZzvy7Z/1iL781BqeRFRkRc40EPByuxNKGTytl
+/OYSWSLoPgVhMmJClctesUCglK6h0WWL6IJxyaDcRMlqNNk3UWqZGaYcznLsSdi
wb9WTiJ7TOUofiwNqVtqksuIEi0hSYo1hsNwXA6EsnUyJ9kmvD2MPEecg3RZSFpb
cxMg4Ab0lC37sUVFW4umQPRCVl1rtkVZwL6AhxIIyBf0n3IAIiCNJ5YomxDBFwyG
37kBXEBJint2YcfzLPWB0UIIM0yqM0F+6HdoVD74kB0JD/pP/rc4QnfzEKsc/RTv
nQ/0fcosCn6STdtc2EUgggJdNKXgrRvlrafeXaUEovP+UzB2Jfh+Fw9kJdDLxPUR
Rj9GLlVGoqKfSPKAmWtfWROlUyDn7JBwENJcHAkua244ajaikWWRbCmwoRvVWMTW
qmOuekQkxBkEZlWrQYAc9zwlv0wopjcsFVQdHhXFbQu0oBCLwxX5RKP0XJJmngUN
yjYG/7Y+LsO2g5Y5UY8St0WRIyjCjQEGw7cf0bin8BqLOoWuXURJXdTAgWR6w02D
9bHRxPYhG5JKVElgPUHQ5NR7JRiw2MV/DmBwMrO/WjDdEGmAtJNEzwhybuYL9OKt
P1WlLqU8G8ouKtCWxTSE73o7ae8CAJB9FNTXN9SKTVZ58fLNeT7D+ewceisCAPOT
OyVEioThQD9la9UMesIzkTFkdMcpoW21fZZ8xV2BFlzuII4CnAIbdEBuXVG/xnA6
LiaOUgTopbNBvJ0iWfH8xB7JBLmFN077Xl2PHeAbkmgAe7bSIScChtTz2WRyCUv3
7DmNhwJoINghfrFvSg3tt1KBMuQdnGWRfd5ufoNGsAIrzFLoiiZnxFuPgN+UmNyD
ziGY/JfCkcpvlgL87ewC7kQHjIuQEA3vksj0Qlbzd9LCQMEE0ImwbZV+xnlN4LtH
hFrgQBKAzbig80UeoJ3mVJYKRSeZqpfrxfYEWJqFWOJY0PmJXK4LRAH4sdXwrX7C
WDAAt4iiAKyUKvO8aIFLxqZ/yZAsbFO26U69us7Thp+HdP+CmiHPE8bnPjUvqwP2
injKs9+kosT/q8VTdncjZBobwao3xGJw6OfeUvevr/2UIbKL/7PlMazd4dRUFAEn
HIJVmwG6zuI8n2cpw2BqPsCTAIyviYLajGhR+Hy/HSXrMnPJb3uV6Gr/FGuL1Nvz
XQv4lMET+Ouk++ytoIJvsigjRLBPq8xR5hR+I+Cqd30KZ03fqQWtBBCu+X9PnkI2
LtJEynMoH9YzM0X3IVfNM8iALRUFXBQbR02DUGC/P28ktCeXJkT1ReZ1CpTa6ii1
2Q4X8KDMskZDTNMOWlrHmhJkbpu+CSneCW9fY6iFaHlaKsBkMhjvXr11hZ58/9cM
g2Fvj61Y1pZeegljZ9vOtlN/panwkqXUlntb7XHPbapp5s0ybwqD33GxO/use3+n
v0de0o9L4JwdVPeOWqSgeESJX4V19LmIEpxgp7a7vzeWYEkCBvx+XKAi9eqtM+lg
zf2cCs/FCCD5gUDjwJTXLQhc0hpS9oBEon2VWZLHamqsKxgZHwUqPwLbOurvbM6Z
1CJUrPOGw4QUVor5Br+zFlqhI42OXVyX0RBIslEnJfpTLt79Mu+Neb/Zeet2ega1
qKft0uTxhBUEJZbieu3MOC8nSq1ch24ILGmlu/whtj+MX5q7FnWaQpmVP7EA1PC8
aLTDaZQPXRusSA0bOdf9z95ehqRnwcCwvhBVawzJjlA0ke5niUT4cU8fkVtNgq04
bY8PCCL/7viDEGEgaxber7dxY6Jk8OlUhQPGYZX3b9ThSowtdegnpj+Ir/qCcKC/
6z7pWT8fhd3VBfLnaO/nVaO6lvtuG6nSD13gYFyOKBezZMYTOznG6AGpJ6C8wrBM
8DCmAH+3s22hDj8rT9o2MLwGXxS1grgfTYEqPZ+D58RYkWsIIXmtat8bH8Y72J6m
ShPqOTOEIbuxpzqkQwCEaLB8zwC3Uu+xiV9Oz81U/z+PhPsklfdEL6xsOnNHip8d
uLKUX5OWVYl6g6EaFbmPV7kOlnfYRnL5MLl8X7BIEeacFbTi0nZsv6OQ2xbSeyHo
3jeuTaa4ysT2xkpIolVDSWqsL1PrSQo8AbVzURGTHoOSplxv0yZDPFIDOAVRqRKn
81mi4Caf99piwNPm7TtcT2otrfaqk5K1tpln1YgsZNJpfnEcPLEbfuajZBzGsIMx
cA5SUo15A8KeQQZSHQ7loHzb2g6DwbzD67/EekP7Eka8qI4QWCD6O7hy0Ber1I3u
+BOKlNbITB+D2aWy6OdFwOcNSuREKRW7mz78j/R0/YL99hlL3dtbbvjqCGKKiPm2
jZb3kiLA1WdMJmt0sht5w3lJjk54DnDnVmt4prxYUkv2oISfBxazhuiocPutWz4R
q4BeJtsfdzanioRZWNB4SQVcv/h4F0PfwNcj+SiMNsEYG4dPOnve7Fi/dN+6eG9h
oOKEFH88zDCPYxEfSUyi3TW1eJuzViihB91SvJfUFGhzRnI+xu5gLvLPUYv6feaH
vhO9Uc6O33zXhfcip72nNbyMd+X1F/5gD5/t0RMOJUEWPImcb5lnAshgLfHkxFte
5xAW8qxI64cK1MjvMJGKuLDJ6KOeQmtq229qdYMBpETBW5uDwuZVvlXVr2+RyZd/
H70iCPXl5jqpGH7XOGMf9InTTmcDtfqZvRj+hO6WokKE+z33GkCMHwb8VkrlYO5a
x5vY0VRtyaTD21T6TNUMld8cuquU8h1Qr+Awrdi161gMlMpbjou/uNMADQyve/VR
JV+XIPsMDmjiqNUtQu2K74Ft06t01xlehSBscsdvj4Ff8Tnkw1NpFJss+VX2E3YA
Z0LE0OLwCpRY55H/a264ne0zo2HU7nLuUwOvk46U4Qu3IcrVynRTd3b7O5zLs17v
PbKCTdUWIRqrS2/LJrp5AC3VQCtdej6Obj2PNG/C2r+3OgvT2qr/SJMRf73JIU6i
IdR9zvMh7gqkUZ8j87EbWcqYXcumuDDu9U5weqxGqaKEXnmRBDEjzWxZt0sHYgKB
RrN1ANE5RNTniEgS5VoPF6GTyaT6or0eed4weN/Etx0mRWhThtGTAMuzZCBFEByd
XdLcqL0YIUzCa4G9zugW9nDZIYBcprOSNPeVwRnJzztCcPrLz2Z/xcsSmvr04HTL
LiqfAair40dbvckc240ECX60AIX5vZnyBgEKlb0L6oP3X32GLgOcEWQisvFiODEM
mAHS7x+mTsCGecg1d1PnerJe6En/TYNgCsiMUOLA8jOyxRZKLgXKiLjsrgJONCm9
4G1eDlVtZ6oA5HOgWJIm0JzrEJJx6WpfDjnQouSOsqyu39eDePi9KQ0wxfj/JozB
a5gqlea5bdxb1GC8PfRpgkiTIh7VTw0NUJUvAfF+5UG7qY81yVOJ472/2wBZCeva
6Gh0u2VWe8EcxVlbE9zoEqDWPO7fcUhZ0GlEIDFIVbqtauXviBYkRSzCDGWVILkH
VfDvbtCI7wQVG+wAPB3yAq5Qj6fythW8E0NW52qQZtF0pv7zjs3XOwYq/k1EER3l
sqlwAoa1MqR2OHnbyMKBhV7aNp3jW4G8V7c2HJSREB4sVwRL6a5z0NyF6XKfRQGS
tTtmstmkW9xaAAT8z+D5zg==
`pragma protect end_protected
