// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HQ!3 \=I6P6\E_@7KFD\U]+7_-69/]80,PW 67 *'QG09)QZN('-WV0  
H]R,%*$77#=@3XU]^7L%.3[*E)KV$$+"RI*M@U7DW\8DYZ#(<U8U44P  
HG/6=+=B?$92Y4O\W95\L3%1F_>+R//KE8AY'N&:(0DXDM&C#:$>4H   
HR7[O.CHCK19L<DPY2M?[S;/QDO*9W4NTRX8DEP8@3^L[^ 75=&"?3P  
H844<C\96(T)*)*[I*T<C1+78T*77HOP=FJWC-9V/CQ+5C13Y?46NQ@  
`pragma protect encoding=(enctype="uuencode",bytes=6720        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@\>QNHVCC:D^V,(>.$';4)<14:(+R'"ZN7;U;:!T6EF, 
@ 1ZM=XL<R7CSBS10TPBY1AYJVH8ML=&DXXZ1YVNE08T 
@,6NM^"QI5$5>E55S@+*=^\A( 5_;EJ\RID#=B?/5^#H 
@N%6]+)#2W4P;CB2(#ZL9\-F''2&[(@NIKN("2(I!I+8 
@GJ'#F8>A+)6DX\=$,8]!JAZ[EM<KU]_^1=*5!G>FJT\ 
@/0H8-#3&Z+$\8R^1TK8^_5!6?D8D&Q::9]@-".!)C/  
@DAJ-&-YI%;P#%"][ON89(AV6/E&"*1JCH28I$(N+0M@ 
@A0\\HFE1Q2FX\[K183;HL,8WA7E"5/JZ%8 \L@Q01Z$ 
@;1 B$<Z7>]\=4US)OSV+VQ4CY8P_(5XV7\U'@U<9I-( 
@S^1_(YK.SL3\J/RGS5XQ#W?M8R! QMGQC$9(FA":B48 
@OW<O ,3LXG7D'I<-OX,.Q?UWN8 G*/'!D;?Y)KGC8*, 
@L5[S$[1_R$'A-"JZ:AMQ3FF"D]H+]3&"25$.<]0]H@4 
@9JZ%?;8,[C2A'(V^_ +M^D<U;C6F*/Z[);)T"K!F*K@ 
@[0^)^^O&5/,OP/&%H;0VEWB67BQ]Q@W<C+0!KSN.2GP 
@5MG/LP-.KR:DQ690+ORCK7W>N[K;'[48921$:D6%4BH 
@H,S=G'-]_.A!J4J7#Z]]C/0]I$$:J&IFO/E('$%KF\\ 
@.&NS%H/5!/VI$&VU\M6GSRC;',( X-KLE;'N R9F8,  
@3;2,^U758Z]!7B)L!+^HH.:=5HEEY.(2?ZLE>=8+L<@ 
@6^5L: $OW9XH65M)Q6&7=$:J1GR,G/+(DTHXRMPJ",8 
@D.2D+P^.^^Y=_&;\J/9)R 8$C!&$0EY)=-L&G*M;71( 
@H[#=C')SAYQ@I*Q5:FM2REY5=G0H%QZ*%M@I[7'*ET  
@51E,,9MQ9N9K%7KXABM?*G%_K 8D7X$V8[A#%>35\#L 
@"0H."0QZIN2CP$B>A&M/MKQ_7]\R8^+7]*/''N>ZIB  
@S2#\(<SX+;B>N*U+M5VHZ<:;9X6B+@ HR>=MD=C3:QT 
@5JOL^% 5 SO$.Y5J?/K,ILQK?.B%",_B RUJE'$&-N( 
@@88/Y$G5,8B=A!:*$=)!*W[<ZSKS"\\0X%JX4<O$EM8 
@:9Q7)M6+HD7"[M_'FS 1C2E:X%@Q$?AK(A9']&<#B*L 
@>NY50<957M*$<# "XX]^>+3>,#4+C55O"!*+^['!,*L 
@3++ 2#CL\UJ]UW[::X2MX*<#KLPB %]%POL/#KGRXK4 
@G;5LNIT=KG->I.D7"1H)(?Y=7TXK89Y<<Q^'JR",#8P 
@"[4\8YCNK)GP0>%YQ-H;"!'?2YC^@L%O:T[#2995,W  
@HKM7<OYR=6J AQRO60'EL.02,8)KM'O7 C[."9)AG>T 
@7] P(K\N)?'@!^)L]]GR\EUO8 'GPX0R\I$KDWQHKG( 
@[-9WX#H-:TDA1F6RV]Z]7(Y5V?$+I/*("!4%Z?-K-9, 
@9W8U@9(OJ#%@)0!!<C W39DCU F,]XV[_ZHJ49MF^AT 
@L ]DN<QL>'2&R\S2B'9/8:+A>B4.D P)XDD.TE>NRYL 
@+_X(Q)2VGV;1%_UMG@Q=Y#4.;&9CP<55H&<?S&3$R&\ 
@C>HAZ7=NL0NO>=K6D; VO6*)@1OQR9\F4HHCZ<^DYJ\ 
@= CH<.YDMKU"*/EVY#>0P596?(8RC4^9D-I#9-,^%$T 
@IQU>VW?-=V%\)S2U^6'RN&RA C?>MFVXM_(RH<Z&.PX 
@Q)84(6:=EN"R7]L4:"!2Z1E&J1^A^0H>ZTOKW+P0U6T 
@$<[]ILID#"_O1@MD1&(8.,35HAY()PY !C_.6Y(M^)( 
@H?V!TZ>8NS0_FDYA7+XTT;CL8U4T9YY9+KH[7AY!JZX 
@HNJ<ZZ+"+P@#IRMER W'R:D&V4_MW>L9& ['C_$<C=$ 
@3YG,R?YG#XF_K:4)[J;WRC"NQ;5S<]_KSG%A7'Z0#0P 
@1JZC#K.*#0QS-6\'F'OQU<OLF@E/AZ]\RRSVT5,#L-L 
@'Q8)_W'"ES\(*@*[)J4<;8/(EX@BGI).D"OZ-/7^+;, 
@X!TXI@(ES2EME7W.Q]W4_S [PP8VQN7N4_(YE.4X5TT 
@".,N<=.U^:N(-NXE285D;S?L( .HP:?@W1L4P-L#+8< 
@_]^@:_8VG$C$=^:*^-!N1OZ% /W<B2'"00NTW:?=TO0 
@DSX% R2Z,.IM7?MY@G'II\9C28RM,A;,6W[YD+X%E_T 
@:/J[H=(6SSK^QDK)]4Y[*Z8A[A$/E_15[?ZV.GGHWN@ 
@_NZ0NC;ATQMHJ;\2@8ANNP2_@@2><V4I:)N6!"LEO$8 
@_(KWX7D3XFL(*>R(,YR@G_J"%T$H2JNYOHW@C\\_I2  
@4/3)@6+68"P$;FAM>1CX<[KW6B>1?+AE-8;([VT'I2X 
@;/.<@MS LS(MN>0^!)4_A:A'C] -_<^<_BS.!JG7VP8 
@"%P>S)U65%G+/CZLM$BN#K^7N73%[^ID,^#6MB\V&DD 
@S(1Y^<KYG@9D<) K_F.JSSB"UOS)[;P?6)#_:U>-@L0 
@VB<18951)7 P\>MS'BGU=/J&'T+ YFJQ(HW92? X)7X 
@GEPG!D>=</!V*@6:TEL1N_\$2.9\[N5>&,L@84!GX_8 
@2^$&?10+W%HR]P(C8<*(W,^X#?+S$2N\4JQJEN@EX_X 
@Y]=/L#%!D8)M7FXK9Y[D3 6D>[; J QFO'!&1BX@J'X 
@,8H2;_ND3ZE (<,N/]88#+YJ5,TXK:36%,2A,CKC/*@ 
@38$G+8YF@AV)I;2(0V(9FUXZ0K9.@QIWD#"GCS9WO@H 
@30( I#X&3@M9 1OKBDC1]'<8[&Z56I89]V/E-"Y5> D 
@5Q?OI7,5;,]PI;1<1+E0!_L%$Z<;"6@O0:8 A/)&4?\ 
@60O""2A%!5N'@YG!4C.^&IVF?\P?Y)(PFL X13(4*>8 
@.(IWLH4L_Z$YPS%I0(8/+S;]:7*HE5)T:+NP^_VT)GX 
@KH#]U9Q'W' ME;+J3G]9K _XG(2%,7Q?*&L0;K0W=\  
@<80DP 0-1S=*%A*>0.RIA1BG>_1R$^TA_=@+/*4D2-, 
@0D>J4]VTM?M!' )(:FGI6 "5LQ#9IBV"P28;_8%W)JT 
@+.O<_><^M,#P?Q0BULB/H<ZA(Y$3*](S)"X?/+I+A/8 
@M1XX.Y%*?BDPA3"D7*&ZM&B;(GM9$YZB7[@V4?UWG[  
@+=JP4$W>0<#VS: "J0E.D#5(88,JN0W0:([6]VE@>9H 
@X'<53^&D5'H[92NY2U'4V!NE=H -,HY6;WGP]("(G4, 
@OFLEX7<;[3RPSIT*!TQY@%U<ES6[UR?'TB<Q2S :LOH 
@PMT,[10E4R<>A9DB6J5+.3#22T<1G\W^27.Y2(0()_8 
@Q%U)F!B%P4DC,>"804^L*'!C""3\FX"(3,UON4I+7/H 
@V;A#@^\DAYI=4O58M=-L/T53(SA'0N(I>0-IX0N_3[T 
@,E),92=SF.B4$@AZBDN5147F/VO^2BTPT5;5,X[PP#@ 
@TR62MJ3B02RF&0%)TTF.3\(!3<4KT_:CJ8Q250 J%=4 
@/K^MM!.*/SKU<O@I\%6X.5CP!#C>7-$7IUT/N)XD=M@ 
@GN"%E(Y=,^EDH3*X)UU>,&=+9G0&!)MS@#*5[@4CAE  
@&Q5LD*V7L3UV+>^Y'_M8S0\(")L5-HS2G!5JI6I%84T 
@BS*PRZ*#N6S7M\J+,R&77#^V;3M(<1+9L"FL!='0QQ, 
@0X.%O-GGF0NNW<C>OT^G+0[$,X,O^799*#,772 D[<8 
@DOSWZIUE-&+,_!M@7\^=CFI.^-W2W "\;#=2I>D"^%P 
@"$W9EO7^#'7 ^2J#9F=LW,GJGF1BHB>W62:22V%:]+\ 
@O2W&N891,9D/+,X)P:#U8J*S6D89"5\\,]4%<)B-7G\ 
@87QJJ3QJW]>4[WU&Z]G-:^,DKD1U\B&@YU:'%8=W,TH 
@1=0MD SJ51%0",6$UQIC0;(.9DW=$>P4Z:E=Q%LOO8< 
@'+WX@"P2+?[*[HRIK6P&[:A9RW?0$U5BB"I[IRL>N!  
@U-R[EC-.:G\WY"> G9#7):;_8!L8K\_\EAKK7E.\K*L 
@Z+NVM\<YJ[KCLE=6BB_.+%U0>U-EXN"3G9F)0=RA4R, 
@_8'.D*P6[B!G^EV+7"ZO"8F@@0JI@7WVA!&!4C0UW7X 
@_:N]0)3P(B,@._/_(DK/M'EFE'K/L!0(?[X<N @$%D\ 
@2VSOH*T(K[P% K?DW+T&<"W].]<O%@:0/[0>'_<:()X 
@M"@0>\_6%L9_O#4L!X^J]K*"A&/D3GZQ3?B[XCH5COX 
@M^/V:H41L:?>&ES48QQ=M+[PHZ+MQ/G1"KM,IJ7;E10 
@H_E.,W:Y1U_DN0#S$KRT( #-W4)ZGNED7BTN6S&R008 
@0/?/8ES<IH. D3-@6*5.D-6XWLQXA">@@2#%NM$N89T 
@?]%U"DA_\\$@H;T9HXIR2"7P'XJAE$O\V UB/A3&648 
@"P  [Y%D.]WP2BT4NE^1:8L1/AE3OY?-;!IIY13+[X0 
@YE58(C8\N,W?'#O"?5Z_@1YVG&.\QIKJ\$ARD17\)!D 
@P;J;J_/(@31"J07T*D9ZSK.Q\X!355":6<>%"CV4FP$ 
@T&')CQ9SE,!>,+C.4@>ON^,?SRE,K&&U:&W\F6A0*6< 
@2&?'.$31HZSS<E;3>*U9&;X0]V&Z%#*:%"/0Q7T%N)P 
@OD$7#VZU/%+(J-/D;1*L)RMD)(VLW],"V?XNMGI!54  
@8@9#ZM]^3X(FD[2Y_Q07SMC?QKEUE]YOL_CJPGD7=)8 
@]"CRE4ADL#!6=8S5['AAZT"E$WAZR/>L)S 9OJ"[ T4 
@T;+M:CR21=\[LT'#N8\J.49@=R)TH?;!RFJ' L0V?$\ 
@K>!! 5!50\4(ZE?DC$Q]@!A]-CR#0L\F0Q\ #0?^2,@ 
@(W]0HF@%%[H]U/#/Y3=AM4GNR"P"/Q/*GI:6U7#MH L 
@'#+#GOZ[;[H:9'_8G0WB<A-VJ\9>'H  GU\AK9&AC7X 
@1-2/I([&NOZ-Q1WW9OS"]#%K/D)2DFH0LA]']JIE]8T 
@<7/P@H(;JM-PD@T/>XPJ'N1?0D4A(DBL=MXLD_7=/Y4 
@)<+Q O&JV0V-#:MM /NFK=1->"Z)B!#T?DOZQFL58LL 
@%F92W$F-]U1R<?O$_KX9!YJ&E#^]S@Y8%-:]^Z/O3^4 
@0,L#[IO=9]/ GKEX=[/U<U:O[JOABW39<S)F[FZ#+MD 
@&^T2,+;I^2'P@U S;AE;CR84/]DQ2\: ;#\-32KC^.0 
@K)M0&W%[W )?&\?K+I"R%.GPN@9[^%BP*.IM.LN%8I< 
@#%>NL<H3<RLSWN#T;ZS-LM[Q[O?$4C1:OXKAG*4@4/\ 
@)HD@8:>K9KJ9#_RWC_U+A"7X@^WSC]&J\U7H]1@5S=D 
@9/_6,A]3\\K;;UOW(;@[S3#!Z^6[7VU*&N_1KB7\K?0 
@O)K+6'785R@N/O5>!WZG(PPV!3-W&E!0+%P>'[GJ[*X 
@\Z\R"SWFWO",^*Y>%GL_V-:*WRD1ZNE1UJ!W.I,6*#L 
@W*4EK9\PG,!1?]E%U)OS?YM05OS3F07E=4+M<"C$X!H 
@)?SN]#F(%2&^,Y=88I,1Q4=NS+C@HO-TB+L<-2&T!T, 
@C:B+\[6>)!4[7@2M\]%ON=(.<B;DFTVMD)9^#4RD=W8 
@=G;I)WR1#VN@],[*:-:OQ%D#6_OK3$)9L*93\KG^_D8 
@VK0?KJ R^R0,7-J%FLD W-E4M*%K777SPF33 ^J<GZH 
@[HJ^=B.GBU4Y?HEL4;RZJ5#SK0'5 *)0] D<+6&#83< 
@D?9NF21B"7BFA$&RL9O?@KN(IWHRC4;:ARAF0E\^V5@ 
@<:A'-!O*\7WW,G%W"!P,TK*S$U$-<(:(PFI'7 $?>=8 
@6 !W7<!?X(3\HA3#R U,34%@^+?03]GQ]8T@.2&16;\ 
@-UN!,Y5Q4.0Y4*$.$U1^^ JC<)<P>Q)/#E3(F<._!S( 
@A3GA3V[6"#A^^10(6JI_FISL7<PX@MD-;W78G%!Q00  
@(OADT)\^?$5E)QD\=AP\H).]3MW8& =M\(E1]@27-7T 
@O^D<@-O4.)_SL^K6 MO@3?@H+2[[*8X.K[EG= 8^D7$ 
@NG8ZA1;A)A_?)9&\=P9)Y3S#AE(K=K$"F:*(<+7N4_< 
@3[R"WLG5)<!P>UTB9N(-Y= =88>_#V: ?'J%Z;8.RC, 
@:1E1SXI'U]R>R_>K+Z-3^@7B!^=S8HS9U!OV3.6W6NX 
@(GND!<,E!S;ZK#\.+CJ6Q]H>!-JK;:9&;,ED&.(CO,4 
@QJ4BHJ:!PHQ+)14K1(9^X)_,:0_BYFKIG11%)4L0VYT 
@@FFK^0_I]*C)(-JJ?)KP\ -;KT<1\9Q9)9DYFF'M2XX 
@$2WQEX+<42/07)3$O.>)@UK6#[S?;('[E"6 CNDU1!( 
@=L0A_*K@?Y-AT_5PZ5(1#($#+&&D54J)ZHOEQJ!<U"@ 
@\LYPI%+X!1C9?7;"@0LO:1S! )F&ZU&KQ[+U>!?2\!0 
@\[^2N\V]=G!,<=M(<XOU3:.@Y(30+R$G=QHP$_0#9[0 
@9-%@E;@OD.,[9ZMJ,]31?C(1!GV"'6)9"\/(&19$OV8 
@Y.H&8>"6&==B8) (=X.6C_I_'^X8E5(6]H>=@>'Z#KL 
@7K87-.JS( 3G\/\WK:JQ'L4YM)L2F9 !U&G+@]TU&TX 
@0A]P0XV^HY6='Q+-U'89%G\5"K %JH1!-[P@F)\/^+  
@ZX'!K@[2TY(AM/Z*5MU<2K8'7:$$J"[=_Y'D?E+ VR  
@_J\NH\[HM5UCQS%XT1BQ?0*'C1$CG^DE>+;+]'C>&^  
@,&4$Y?OGTL:QNX\!5P3;Q7I_$AUPR1+GRX:M[=>UC>0 
@._%YZ'[M>(HBR/243MJ[AT3_[J=?BW6H?7?R\T+]EW, 
@C<79D?Q1PH(IR!,#0E?9@,?'HO_7FMH.V/&S%N-QJ!X 
@9(TPBF6\<(2H":?RBM!P9K16@6B;SX@7D/!(E%[&K>4 
@12^9[1*B=UQ,O^"\=]F_4PC8/-BCZ>%(48&GRTSB^&X 
@]8([;1F7KIU AZ7:)ELV#/%]D+4M-CY)Z'\A)FCL*C, 
@KU8AFUDOH_HL[4$1)+)QA#V=0.<=96X=AAD,PO@1;)H 
@W0Q?@'U9.A$PGL56JTAXG.C)=['[.@1:7O$M^W9S'W\ 
@UY-U-YO5(48-CHC8@XP:S=*W/ +$VZ@E4GR38R8-@2, 
@?")MP+3GNOE+H35I7(U5CK6W+:B;+)HR/3Q .LBY*8H 
@B@)20=$"2*<^D"4 1H_%:. /EYH]V\MN7!7'R)E;>9D 
@"XB_\NBOI-M1[?(-Z 6 WU+.?)_(!=9ENOO.TLTI2G8 
@BY7(Z #1P5;P<<;QFY!(#KGBE'&ZU^7V/";_]SSCSV$ 
@OY,@+7T9]-:8)L0!C40US@JA@@=T&>F=AO4#,5 P7L8 
@-1$)V@6:===KA J5?LTJZXJ_O!#-( 1(D-("_^_L*0  
@8[P?.K?+V<UA73)>Y::,#YI611'BCO6AIQ3/:-IU//4 
@#0S>8@5XL"WPJ(QVW)O+2L5O%J22F;5K9?!3VZ*J:K( 
@H"?NCB(D%X3GTA0/8W,5Q]O<#>ZEE%OEO\](+5#5;1@ 
@R_=;EL!?V&\Y^?LQU6T'#G"V$L,S\B!PG;"DZJIOH+4 
@!MY77TC7S/-)<XAYYQLAC,ZRV0USNXI@!FN_E,-VA%0 
@:28HH2P3"N#\ N?2&">)0"<2NFWY?_[F3OV6(7_N[?H 
@3@36FEF1W3]=HI.J'C@SG/&\X[A<)D.#MR-(<GC$,0X 
@,TA05",9[&V ZT0TO$A'ZC1EXP[G4GKV]_$9^FI[%7$ 
@> 7:4X$(QI[/<431>+OR/^ZIFH1D<D?S/7P^+GYJI9  
@NX0S2?6K,",?Q8HZX8X%H,,/XWB/",/7RQ/\/)$<VWX 
@4M,JT@T?#JJ619I%VU-O-A;,#!-;Q=F'W;+C,8&]ZK\ 
@1G9OBNYL:277@AZPC#=*=6&V?HOI[)4-(QVRYJ8(C $ 
@LW,.Q^)X%GS*68VS,EN<&6'ZS* _XIL>Z/2\QV3;%40 
@ET?"B _9Q0\()05@,8U;$2A53UXEESZ=P8M)X]=F/0L 
@QGTLE+ G^N?RK#\VT1GT+,\8FGTX\:#2OK\R0\J<O!4 
@I9:;^6=56_;R"#%?OIGH16UWEBC;P?>\C+'56-OS;7  
@#G 7MRK\C?:.2CFC;T5UDQ4"]4( 1CT67GWP5:,F6T4 
@)2?IV5:!\-I-M?3)'[C1W'E+7]"W0G7.KP?6%G7<2;$ 
@?1YL<0Y!K/06AEKPRFP>8"J:C-9]!E%G/R#:J/:!!7P 
@^\5<)VCGPJ;8\WZ<5\;#9LDCQ0I;M7Z[ 9"#HL^X!#T 
@Y?N()+_)^NE.KVD4#C'IA7X$]:C!"DJJ$9W;=(A'8.D 
@U(?M)=53%=,[,;7W;+K2Z*(AZRU^PW+WDXRJHYGJ7+8 
@)G)/YARZW*U#J'01YS"S*"3-TA_,<I=VRFG#V5VBN=$ 
@-?G+TE;45%/STMR?O EK5!5;_VVL0Z&W.1Y,4>.^+$P 
@:O+;OIK?YQK-UKAU;H7K3J7&/&:=P5>5= *=UHOM[L  
@AC:]=RD/>EUI=N&3="/3 A1V01RX_6$X435>^OVZT+( 
@B?Q&#GDPN: :D"SJH46)C(VGJ))#^>KJ. [29&E )K@ 
@CGXF>X8:<KBQSW.X,H!:-=)-;U:3L*;';5Q0G2:0&;8 
@YCV16WW9NFF3(..GT-3CK].-AYB>'.,P.5POZFQ2$(L 
@ *0E=0F4T:GO% Y:?P81.X+\E/&NKRW:X_B@[SL,3D8 
@(-]O=D0+38L;-T?/%%OFUIE.T0@5AG2H_0 >4@'9<>L 
@>(^0T3U;IN.H=V6YBC;M_#*.YB'MOZ^@XEZHC8[:0\@ 
@94F/S1GLH:4%R<Q#8&4YK.!7T5VX>"J4;:.T:$>-%'@ 
@4,CCZ(JVK29>G7;Z6^6[B'<;VIHL,E/0PMGEXL>U&W4 
@LX0!.^MNQISO$O9CO%>3,M'.!/L<+H;Y_( +-IF)5;, 
@]T=:^J1V7?06B"" 6:8TEXILTY I-;ZY%HT%NZF;U%$ 
@OR>C*4&+8&^RWP\*2@=/K[)*1+-_BU%&I#*R!9SQ$<H 
@D3=:NWCUA-A5KF'!-1>]W=%I;0_NF_]E9E<)0:VT-%  
@8WV$HW83 M[)O&;L(,\'7X'P>'F!)] 5X@M$?<;E13X 
0("IAW]1@Z\L+VXG5N%/Q"0  
0(;L[VEZG5%L& !F6HY!BK0  
`pragma protect end_protected
