// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:45:22 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fos20SFuHHKwaiioaQZ8hGcq5GoPBtxQ9Sf1mV3jFqpesGYHCLqOA6MLap232Mqd
RjDzJhlVmp/hjQC2Ej3WHNky7fl0TkiG+K5+H4QHN8TmMwKbzDsRcQJ0ZGsiYt9N
9mpNqkTJ/morUeJBx/2fxQw6JL3PYx7iuGCGAzH3+l0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
F4FD0c79tcZcEjTxlSjmxu2F016kDahABsEtNIgbRuGuLzShQHcLKYxbYQGIkbG1
jjaSPfiGPFmkcWHMMaZZthBWNTXJyos8J6ItazhFCJ3HDpVyh1oqZpP1f646LwUE
A7AQTqP+G0FOnsvdku3XtiwmA+7I67xhYxC2HY068JfPzy4bKz9Aasx0z/30a4Jf
ydtY54GZacfZBVWdWCi9yY9lgj/RhwaJNgMVFf4NPMe4OjfID/q8pRFxGrBFL6Ly
ZR1XE1RBY8AbbWtaxaYAWYx2KEGZn+scB47ESlnxWt4NxM9WcKBBpsIdrIQ6oAvR
wJ3BbgiYhrUpY2j21YTfZgJheSuruT+qZZCD9i01nC8tbfx3V0f/fZOxWQGe4f07
m3jqkTF3KxQ+NA0/2Ps16zpS3b0tPQGqxO8HALVi0Xeh3irRMivG797XqyifDrca
EVLhQIJr5bU33MvvHtH6dtTJfL/Is/Mor50LV7WSpIgcgG52tMrZY3LLTSjaZMbm
rd9Xk8faPFs74sXTTspLSi3p6gShxr6mJvuwVyp/4Fhr8OZ/gOJx49qEtwbZKbSF
ziwO7osy9FdTV6/JDBH0NNiCpoZAaFwX1DKvcE71SttGwsxpFNr8MEYlpyYm3txD
CpM6Gn6WGqdcwgxMMzN+leCNG7jigKzCwIrer/mq+hYqX3mM9If9uVT2OqkO/y5R
fPUpafEGnRPGHnewNxbFscTtmOka8fcags0q8eVtr1PZMYvEXvEomLzYmO4VH81R
8nnwCFhFdqPf/fSK840DWF01GiaM9XAcPSZ5m1oy9ueXFNnKRCj6GS337UHp3yas
QX4R0gDZrOArES9Q1Mms6+aav7QAd4QFdZeC4RgvIARFdC+TPaQh8m1EDKLZo98p
gPvJXhgVkB338TrTvjyiXEcFnpc5z5fbUNYRIkD0w56+F1pqwpNP3hLwTRPvUecR
l0/iB5ozST7B17oqoStriQUGIT3A43zYXpFjppn1lfWAhinuQuOZjv/d/qxHW6e2
+eDYwEfW3tMqF39RjsubD+IXKvJ1mM4Llf8vBj3jH/q1P5LjV1WOf4qhzgnj3SAs
d2slRUuIZERMd/N9vDXyp4lI3SdKEQJp3rvFcgIQLTXqu8QDS5UVLCvUPLiRSqcC
wEDc9rZwv1JPF+OghM/3/EM0P3ShRHXrnj12ZGUEIi9VVFmYfB2NTo36FiFrC4OR
G3ipl9SK4WggBNdej0pPZVB+mU+BjQHbYwveNLj7IjP3xftHwwzrftCQGcHwgAWI
rNzIbfzNIybaaRxQjgqKXQsFPbAD8PlbsPG92zdkPafMOeIl9ZWc0yyp/sCk1M/c
+Ixg1XoYdQNWzS+tJwohWKqVbYtgVnSeUNwiGorwY+NrWD/xy4x5v1Fv7KSLZH4z
4P48tooW25lzo4fh3ViM4ZD8rvn2B4fsw3ia8bf1jw9CG+bX6n+C+rPexyx4D5M8
w+28QqX3Q+FW4tdReCgnUSOG0pWKvMFMIwZkmXZn5GJuuSThuojfhQz9l7DcPEQX
1NuiJffg9bAnkAf0JWM4memnGU9lHn5tkUo7KdavttJs1EOQSbOOff/kB7fN9+yb
gOUfZJMTr7o9bTjhaeG1HCPKZ+2872H+waSdXyp68BDTaH69iC8VxFsC9m77FLsg
RNLWue4DtbCJ2awYjWuer7DcqarxaFXXaZ7KJ3hK5QMEpPnGeH+9CfpIQiStPEuC
LDOty8BdwX9+vyJVg9ELDx8cMjgXv6iGwwg+r+JgipguHecRScRXvXPmfr9keBc5
tVunmFK0XACx8xz0mEObXMWp0DGZHcKD2anrYTz9Uv2BdbwmzPcZdsar6GFlfh5I
MMOktLZYsAph/Pw5OS66oiEHQZDSe0HYb3xDEExZ6JWL0A8uLfq+tYv3TiEmIRZz
fCpPIqt4QI5ylDC1Pysup0ZGIc2dSOzAAbfcdnN9g8BMCNXvfq45Fjn+icmKeClZ
R3uAY3aBEH/naBQWjyqxhIJmwqIhCf1EAb6lyHvTc6xBnd/StwPkxh75/PTlrTBy
USpnpgX0IpvyCHpl83QX8z6n4fbL9227TUhFF+9cSxDCrhnUSb62ulb0tNq2oYrV
Gr6lGnWy3NgJ9Ki1lFBkm/jzLlnol0LZ1AzcknRcccPt7PW/L1tXOxlItH084T5R
majjb+C2JtM0IcBLD+BQSpmV4VhWkMvgkb/GsYuzE74VrptuocFMrwWviAc526Wi
JXyXCoyZ2E9J3XnvEpDr0X97fnMOeUCtZxfARRSMiZopSgf6GcRN8SjXXP+ASJB8
iBa1TYzChRzxFSFfcjij3YiikoUpQ3l5IUJZl9NEgG82GXlgooSo0rJWL9qtamXL
oTggnmSg+V+ECBy3sBXtFClkIUAMixL3T9tVudfAenCP7BEy30CY+7eegMwGgupt
O8eqj1szHGj280K8ggPaSg25NQeI8upon9SPvRXtF7RKUhelwMufQO7tiK2ORggp
Kmw9OS9Xwtv1MqUc7WPXbbO7kyKHiUCtLC3mkH3G8WVfu2z6vVISLpkmFCMuaw4r
alJz4wJXfyck2B/7qCzoqRHIuuzk5TaBMHPJ37Qp02Q6o8JxM3kDyLUq6ppw3SMl
G/54xM1CVeJB1CGN6OgdNEpyrso8iW7ffWCtzp9PG1MpkLpkYM5FLjSc63CGXNpY
t1p7HTWJN/tn4O4xifKXUW36rohjckTFZ2nn+L3n+R6XREUSnU0WKC0ap3SUKkIU
M/m95Jpt0YmeR0WIlcyxaYdAajqNpKEC+LAwdTda54JkO6hhxrWLkcYnQYgO81m5
FlPMT836fWuDaW7/tDB7Gfgenrqi2X2H+YoL6MXOQB+4LyMPVejVG75t3tB6O8lm
2NT4NJ6mKxZMIvL/Su9vZH+eReysiZZXMzVVIwgMJ8CwMyVt9OIVoEpTv/A+lzwf
UbUKB7+ZmuR7cKpGL5lQnWmtDkD3ZUqofs0ZL/d+oOmvva+BhmApLM67ilnoIW7O
2EtgKDFdnLM3EoFxspq+uq5qiKjRDWOVfMmNT9SWEO0OZPVpPnNnAi4uHI0bqGaz
vrtYqjNzYaOydWgWAao0kC9fwI5a4AzpSZRYY/TWOJP9rFNyzTpsSgW1Pq5dbvmt
sBa0VjXrn7T7tNK4/uhNgyOccMUyeCTuoSYrZew5nkSazuYR35ozA0A1bdyN6Ul/
AD0+gDEeBjxfC5w/x/q3FOo9kpTlF7X7nFVLpq9XwG5Bxh6bV1O1TONMXhLwjMBF
J4S0ON2KO7ezOLGz4t/CIF5djtEoTGH6TpcvvcmtZiBkyr3JxSKoi7GmQyvr389w
Sh0NukKHRjBBndjPPw0GYO19e7nT9RoQ4s+kgMknuWse8jjOxhFRLfq5zZucYyJb
msZ6gccBbOZQgDVw+NB+X3vMf+nbac21Qh9m+h2TDaWSNAWxlg+kWgwInoes+6FO
h0hq7nPd31FioofVh6WCRzGuQs0ITM8ZQ6EAuZxVsRg3PDgA+4Vse1F8ppsT7Dn+
CIKDNZYIpvJvpQyMtLCMqb/goEBrBmR9X9aSgkoKHGt9VLiuHju0Ceelb+Kzftae
Xj+uY5Ib3qUYLYovvvvJQMCWDx7BVCyJPAVhPsdeAjK/Cr0R+wZN34roa7lHNSdw
ISMjQHBm3W519dbPsh4FtWBmg9Whv1bnoraZZVgrbId2KhCcH3yD8UtgYc9b1j34
M6MR2/pzHcrUGUqw1W9FVr1sPkY0yYDiFc4fDjPqHNPtj6ld1qTYxhdRhXYhGJIp
gdQ/XTinFmiVuQu+A7cV4/q51H4f660N2+BOUX33kTG3H/c6QJyhL1rvFEKrscSc
zjKafhGkDItRxKyqcCyO2349zkUq+bN71bPhmD5zhtYZFX0Ru9uDGQKzikXGXuWW
PACx2tTUX91ETLMyLucQhtnf6Sjvk3nPbe50mG+ewbU2UfP2otw9W3S8N8u4RkiQ
hThNyqfTFtAbyYx5ZGwnpJCeT4Hppl7cXlYmyCxpaXAC6ErXYqG3BiL1pnDfdZKS
qA8a4zZpfotCtnjyw1pAD5xI6cTvMDYCnaSlCCJRKXa38xZ97qQ3E+xf4beTZzUH
ZWAf7Q2WkaEX9RPRvI3CYHOi0TTgsdiSJVLwpkgVH1QZhbCVMShh0LGA0OZElgNs
R1szck1t7JMgOLgRLiFggSPyW9CXOO00q69B9tCnqqB9PZPHv9FVh1/8xfsTj/Dn
sup3cQd9/dNQ/IkxTXW3GDl/qsK/kBHVE7Tnrm84Wy0VmyRiJiXP3RXXZBpAVaz1
BVJ2lA7xISSLQ/r5p5leUAGBroyrBJPB6Gvar8bX5RT/hWuktFLkY9Jn0rNUm3ly
5hew2lAV9pFPY1rhB2eQPjBeX1f9W+reylD+F2EOhK2faxfKC7GnUS3QhXNQHzeo
fxfS8oMgooeUo9NobTqYElF3digxbaIKkwUjTUyOS4Yi8kOYvYY1pbZ+wY8HYEv4
FfASzWyJu03Crd1gslv1iq2glFhbq9RfcgAWVjK6bLxr/d0xYXpV9dCZ/R8Pl1Cj
AYjkGf4JA2PRqIWN0oczYNajg3I18SSmPoiHdyfGdUvp9raYf25lQithAul44+VM
2uPY1m73SWiGUgjR18yhyo0nqzoLbXzMO9EwkQs5fTfDT2MNyR6fHr6DHAJXM4Gd
YuevEQQs6PxIeYhSygU5dwGTmu3OqFk2mcgfk9IYRW0hVi/ulBFWRAjqOVb0qnuZ
FUMC+X12d0Zpy1Y/N6p4ye9+NKQZfVk1ehT2I/FUqf8enSIs4PCPvUKntw1JH/nt
4HgGL1DrrYYWyv9b1Us9o3Op8aVjlyzt1Wkz4FIn10v5bYAUoaejZSMC9TzXsb99
bSf4/aA8DFpmJlNPisbztZKMvANRP3lPk21bcQN1xtzfeWuXMy248ywmwbUisxdn
GKo6IfHiULFUl7B9fgjTcteid4DgRSTo6X3CinH/12l52huLvoBGykf3UqQPi85/
HXTt1gmjY1P7Mq2fMupOeX9SjixZNLdTdxJEMrjF53kTx+KryjLprB5kaeHMAkhz
qjh9Ly7nXSqHytmVrIiJjFz/46Vpj1a2jnwllQhHyQpztcUid+ZXW3184TPSE3bW
Hc0OTfsJbIZ+i4L69uPcaKLa/qVIYBqvxBpVsOAs2wDXe6SFKXhTN8wmzukU9mIb
8DiNLt2vkayvOBpVV5HkGUgNiQaiaVaXCytQRvysdvpatJ74l4zVIQHvr38TGHs7
iSLBwZ91LI6n0SWHUL5pUb32utctHFj93PtcPqxsOLBPacbIbLFiDwA10bgFfobG
OzGJ9YucYYr+7qN7GC+XKC0WMyuugqjoVPQfAtN28Xj6gNkmRj9hinytrP63lo59
x+8/GBy8xp4O1QQSKrz1qciRrK11lvFPUrEBKfMevIWqaxty/xv2xYe5isF0Ni2h
rXHCZg85lAvjV2xOndZ014IdHDH67NcsoFQy6MLe1dOBw0p4TN+ci3HtiyFgNztJ
B8lbquYDFt0xENJVpj1quN7FfgTQG4Q534LQy0FiTB1Rg4rjGdT6L0g9LDQnxBdE
sFU1KrCOLSBWtBaY/7GIzD3kbTLVpooOTqHBqobOuxLmN7B0PqKAvVLHexD+luw2
P3Krz59GKq4VFWydI8cegR/X5DmCeCd+rJHY/YARDzNLzduUgEdRtUXB9ay+daHD
bM7An2UbxAOSahXoXtKtoe+b/rot9IggLxQTLDj8g/G6FOo/C/sUiDM470PIv4rN
zXBwZFt32SRsKPkKz+5Rz/8/+1CfKRT+QQTh+WYxxShC4g/dBfRfu9mSakVUWLpF
/xt1PxFzF68YeeNvNnKy7uoxAbyGAonSN1uPV5lMHObs52FsRNt93ZH1l5Iw3g0V
l/QFlVqC2L6G0lNeioPgPwPbnnpblT7Oqo2eyEdbmgR1LfkPcOyjBk83BZ0Ovvfx
G0isSgjM/gGqLYsnaeAyoienAEpOp7yAN5xTXPMkvP4DI14kSt82jKRyoJr1Mci1
RyJ/jqywWljR0lfpClKonhP8flRe8OKl3A6B69p3lgkDHhU3nXFJ/mvIgbS0hTuy
xoXyQljF78pmMDVR+Fy/x+rC4GL14MXKGO2AUgwrjubEBQXsJ1JClZJZah6GQsAS
qFNfnaZ+US4E7katX1qVMndoZnGyuieDoGn3+4yeIZ7EJwiqE9UNNhBrxs/f1hjQ
lIkMwQtccYb8Q1Ew69262v1RHpgq8lfBuBTTbVXQQPmw/8JnIJVsnE3PjqxFSlXF
Ci5hwN6sW+NMXLU47VCx6EODUTeuwl7au+rHv80qVsaWhzkI+BVewxZ3Q+sgMDwL
ytRX4SBLpumCdTR9c4GGPcV76F/9wS0SBnojaQEKlrj8M9DfVhpvinyo6vDSePU3
EqEtPRYf8naw9exkDVqwBVek0YKVpzgvxeekE1fNAMiANVjwYN7bJ4oL692tZNzo
sTU5RsC+zAoRB6jV2smp2fd61tHciY+/Yv695ROOlJCqZep+bq8bP9GD0t6nTqKX
3T77SN6ZqR8HXUoGC/82rJIPuBAz3nPhS9+1Lsp2Kljw+9g2v9fXwkVHpXp4O6+G
5sNQj8lw/06jI6HLOEFAJhvBvgIU2ZavToiAD/7RFbI8733RVWEu45DoJdrAsfW2
tbG4JGW9rBfNrsZ0C0jzuB5/KeGIfhHgj0ulQBIabuaoKqGOuYKLyHJ3EpwCPdFt
h674y98WcAQKpI8jTEDo2SjOH5CguCPlqn8zH8+PsG2valGtkII+vDvCqdTm9pF3
XgFora3ImWFnJFAZj/NJMb6DtYtZU1UJWzu7G3c7XOifvCtK1sl4oCT/KfBch5Ct
kPCxmMRTXjCyUSKdykI9pXaKVnu2E7zgw5JnrDm34V6Lzy+cV975BLAKJC0KvU8E
QhGZk5g1iFZ604GlCmveatH+vHSFdIOWu9G2MiGa3KdLHHjCuJedy8lKUL/tJhQX
+neUAgR6fvfuVxjNENJpbDRvGslLDZP03qfEy7MwYv6LSbvZJlAC+C6i5e/oAgOG
rg62nadcks5PUxUkbH/JSVQVp3IR9nUs2Y4ppDB2PguoHG9SmZsvSP6QGAYAzAPk
jwm5MVIaVaGQmS9JrXmYavTxm0EYX9N+okNXhlTbEwp8h1kEHVURbQPMmeyFX/F0
sEWapOaC48oenxaq1Da2EuVIDn3+DhlStmTyzD0+xsAogEAMSz4xcTkOqkfrS5Qk
l6tEJslMOM4/f+nTNbEZDvgSWzELdiBnlwcE43J68Nqj7Vy6X01imGnUNcPz+ViC
+Wn3argS/7N2SPjrKekDC4mQLihgg1Y76BtGvX0FcjUSbY+mQId3tF8ynomDkXNI
Hi9R7NvyrmWh+Op/d6xNg0KF2gtQ7BBjYIDWCj6XxQHHVMZIwzyUqBTxVPNsuNhP
tIsEax2wdv+Y7HpCXMvSOftGYJGI4iQqiwhnUwjVFZiBL9vtGvny1XLi1Y5jjUOV
RtHaFdZ+iwHqZ+L8Cphvg52wgodGFQ2bZmepsJt+ARAQ7hhTt6+A1/o40sVK+g5n
82QWfhfdLJLrRsAnRrGKQeojLVTTUCeh8cKbZHTdGBodDzLc6b1vkh5l3/AnJzcM
bgGrusguOlQBiEge3RfVq9uY7ddU2+DDcgCK8Z21goJ/uAB3eZyQO/dYYRUFsfa8
O8+a01rItbO6BzcX0tVEXB9MF3VA7rp5404dU1wSklaFMK+XXozYSWDoQHKkFBT8
d6+1Jl06j/yu8mXZb+3lqEVJ7ILGTGQ8lRP3r+jDxjskZDzPVpX4eMhXg+obwnZk
MySI+l9kZedtR5luTbntorZoNCosjA2yzx7RFgRSNLKSR37mhULgbVPcW6oSIdOC
NEpNL2htX14w6GdxAPiCjsk7HWkB38I30bIB3sA0dFEJvSgvU0CIm+wi7ZTDZc/Y
wFnDSw9BcAHc8YjkOR1XjjebGvL52HAzJ2w6d/AOtBfnZID+HY4yGZ0rsDI74FFR
yUVwppMWw52oeto1fgyLik2PDVCQzM6GcOX24ztlLJj5+XJbMKi1isniZZYzfMFt
fgashBrh3RYvXq3OI8a+KcAwYUHpj0HfBUi/wfMIUUaSX4Hs5kE9ERjQsgifwAGl
1nSyvEBtdv7bPonexK7HcJHFeMVzFMRZm7PvvXWgaOeQ8QoTToLrmPzPNGDUCgYd
F6nZA+TsDxUI08AmJbI3LZwHbmt3Q8XooRdH6tkCzo89WJllMnDG1yy3kqVY9Qj/
hQdq7G8yP/G81FZa5TXLGWDPhtlxD288BEKo2Om7EemaKJhKuVvUBg8ymAQ4zctr
FjLo9+QHRBgwQfX3u54V1CBFtA/PUbYveSRN8298V33d54hUuXA2wimOuVhG5lZC
LkvmPAmdOzxIinW8cbtOABlopZ9i7tWFmiPl5Z5MrNiBvkVAZtW3vMPfegFDNZVX
NeFNPd4hjvlOOdTFTb55qJtkv+87L6hxtnsmCCcvN0vVeP9BT5c8uKQedJ+2FBU/
nGS7X9CYpDRTbmNryYKCrBYyAMCl/EDzd4JKVIaN02V5LDvZXpX177VGZ5AscnSz
UbiLOBZDYX9IvmDuGtXmxFLEKtkxZZ8cOW2pHRUIV9r87b4SWKfZe9ViSUA0NgYs
5UzZaaosCYvHICtq9XRcC6pMqjVbT0JX57VERBUVgyU/r8D8YCtx5JxK6aeVhH+s
f5Dnm7rD4oZHVfFnEeSGkcVvHfUqmYNH1j0bq8Tte7AoHmsznXzL1cufzbMedKTG
oChY4JIQP5Rn3W3LS3CIGTI6PvYVKNADXVOnIUXXxrja5XNR/qTDtsrbhODSDejD
T4e6uUvudO5lgsHpcq4bmiQCgUpHwVnE/qHO3MB3cDFo65KbD/oj0KSsfn0AZahj
xNjgdAmY7ua2WzTVc5nEtHTkmARSDZqll1PL4Rykd2wVltzWiNFACyh5k7EqgYWr
h5eC7zd6Oha8QuymtSlmwDqvEuE/PXERfsEBW/pzY+1o5w1rQdmnGNxWF85vmk4y
6X7Z8MQO1vNA+Zh5V6EyaYlkIJBXq0bslAAb1XaicXxlZv6pGFoNJjh8o4BOUvMS
wKX/Ax+alDq4hnZGoIHAkWDuZxpQT3SzmYJf5QAazwU6A3uKWXo7GZ9muw0sNn5A
JXD1fW9hlMve/xoF6vOk3KbkNmsdwdJnmL9YUr9zfBL6EG0TeAXdTnHFcQcOqtiW
Vx8W8LDm4jxGoBzn0cQzVgi51rp3z3/1bcmuOD1AnTfb4LeKXW0L6AAtweOKpoL9
zR/1KN/6HQVn6+UtvK47Acswb62EjVdH762fxVWpiK8m9wJbT5OkDpLPkLGKR/qW
cld+snA33WnEs0iAnPqw9yPASvjdM3DhiByyw1qIk0k5VfxyzuWKMBccK9LFWVjY
Dc1OlTpW8Gt1ijtbTK+nfNpRlym8oNNdsmzoDjHt3u/dHcaUJwhFpww3GQgewN3z
B52iVkjDYZTx5lajQsAnKsseUtt9S7DjexAi2QD2KmTzj9uEiqG2XB+VIzmosTf3
/xASnhlt4zf8Q1jjMNZybZNCUAScL1gof/kXyNC2HV02pxL+iOUpt1GCByoW9Z6v
MzpyJy0xelOBQhaPVVpN/oCSN12c+yY3D6diqfQED7xhDQ3q4VOQMSXLv2zqoNBs
P83hqDFcfZXkj9ecQzFxhE31b29AqwiqbGl0cO9MOnQkp8M/LZUw3JNCsLBobQkY
heX40LwZZfsVHV/CSQQZmXDDPto0dJzW2obrJelRLyBRuLZduEPyUx6yEHwTSg2g
iuIvCIkZHxe9WrF5UR6tvckeiPSvcTawcNiCUdzW4iB2IeQ0KDF6/BPhQh/TJ+lO
NslkCDn7eT4mA5CHGrMR6HFu4OxbhX11SE0uVfqLay5Ck0OTrXfui2X9OGt+plNM
UQXAOfL01+TAQilU1+XpL3CA0rJ+x3gsIV7V+HYThLP4yTo++RPnmA1mYDjybAxk
f+cVVIPZR6860LOasB+CWOiNyuw+NTzdMrid1JQiNVRsUA58KRKhDouIrVqtnZWt
8mvhrId28kBjUNkwoFUoHu3Y982xvywb3AiKEg0LeN3Fj6eOczIgt7uHa3PsRRNJ
5QAPytFY6G1sY1fKaoF9QZwImT5TjZal+pQfprpFTlYSugS4BB63xXdWHjwaoQyg
8IivissGzbDSgpvsLl4UkGE5aaRKnidX+ls+z9K6q6AclYjL3fsIgOTXclkPWmoD
Lhlc/eVGZvZD8yS0v6DUwvuK+r7m3qPSlaZ1S6BGeRPEGl1VdD4Zr41Rl/5O16zh
SwFJ4dgg3AlcvwgCozpqEGtfVjAoU1yMD7+kq0Bm11iKQH5wbRxuYah4w24vYh20
q0wIRCVGzPEX0BLWPDZoevm2NoRIjJSM5TfsMIBbJFbgAdOE1IDvGMLC73qxdCXz
EcIn1SwFzKkTP5+IMSfq+Bwvgn4QvBewuWenBwBr3gFUByNYHCNzzJ9eORVbKjEO
Q9Ztfnp0CmCWMl1APS/fGuhkbLwSp2BwT2Zc/nYOH5DAqjFzmYgIgK3pWMRfojcn
N3cjyvnSAEsh5VjDPfUIj50VXADhT0Fv3NINx3NY/8G0Fw/vrnJdq1GMZIvoL0iS
+V5Vs+ifGI0WcjE3jxRM3RQmAHK9um2SDHTFHKHkgXVDZcpHUCXN18p5jwz1DXw9
ENaWGCn2jy+x1vPO+O8uo6UF9wozLhATX9PuvV5/zwalFbFuhSpZSKN7JIR6B4Jw
ptYLrrPJy7U4yPjI4a2BYxYcuiLAFRSGnNR37+kMXwCfpaqlE0svKlCNUXEV5EDa
UF4c4SrveGrqV9ik+fEQnp4lVUapM6vp1ICuEjqDhtcf//1VxlMlP2zR3eHYhAzN
CS1/UwmrrpHkTSZvZphX0VovP4Q8BnvPA9v9kr6GVrWCpBmFqMLqPrHALDqQdwwk
XKzgqZtQ00ilWPaBazrPWrLjCOxY8ykBVTxyz3dpejozUPYcoCVcSpMExbo7+1vg
7XYyxmFP4YfvwF1kLw7zzZXAj84y2DlzdAtA9xFYzc8Cnvcb6s4UDAk/n9cBO7e4
UN+HMjIB8BkVXAB0Wokbf32ojmupUoXvEJffXYiqjK/CcEv3vodv9nEZByv/Cm67
CgG3dBKVNZJq6QKk/LgWeaXmaH7akWjF5gR1xqvrrAnLWUDAk/Hq5J5WfVCxlQYz
SqDCT2Wwp5E+v/c5JNDZOrqPWma6AQeRZjM9Ta+Be6vXkXB6I/+xTEqpyyZtXV2p
NySv3DF65uehx4OK7BAtErVu2/mXMZiUdKlj92Ds09sXWBkpda6iCcR/BDDq5C6n
upFxvZ0V4yGSwExNq9J47LYl5zQuJekz3pMdgRMewVHhx6EIN3zADW2dY/PNopWU
ERx3yVyOqq3S2UMFewPQQbMi+SUUkgm8hwZv2Ycjm6P4C3r2kDPz618FJ0kGFAbT
cGTG6MmZOgw0sA9SX0a/24Z82Eh3vV9KVaYE4kaBIxrYqn8HEFv1qSxNnOGIIPqe
vbyk7L+7Hd05inrP66/t4VpWpaYOlj//pAP0QVr9+iP2/mRHGuD4On3nLWi/OSa6
40kvYBChv4WS1EGevmke3XzWRvSxYL4DCSE1pjatk6haZkCy4+F6994eBVSqYB1U
Kn3pyeccH+NWji7KQYP/rcDHewidD9uaBKEUCJ05yMt4FbYLUDOJWvBjRZ4ERFDR
NAxbGqvVgR1SsCT1zpNigsxEWYwu+mrFeFEmWzgyiUyZa5tRM5X2ESesqNDvCDm6
Z6zH1ucFA/E2d/wJ3YzqEilId62QhZY/q/KNaIIj17DfL3+OL0BY8M4Zw3BwqMXI
YIrf4OTzwpxDAYdORXDCMpjgg6TliBLEGmqaJ8YNwM5efdrjbdXtoytatBFbLtrq
2xew6aE52n+4Dy/5uqvjyG3n6YTY3uMF1vn+lKQpHLJVSOP9waAT4lh2T+2kGztB
ukRAxSvhtlkwUC1qkX2ty/jufweIGloiZens6VoxX1fUGQyrKMIXMqOVYTcpzdBP
+Qx2xwRzXeyQDdHLDkeLVw8Scj9yQ3uRT5Jm3vJCoE26gIqFmVzEARD8RUOxUFeK
qhxGXC2i9AWdVmKvImOjgVlGrtRRTZ87/Ioba6rLcW3d37+hBatnw1+NekztIya4
9j0FoBi/GMw40BiTe6DmwOIdMp2xHWl4b6yHj0Qcps/N9OM3JT44PJHCmxMuYwgH
xKJcg7kK8AIvSH6RxbPmeJPf/W+O2++CSZOCMUDCIBePcaJZeUuJz/JcnF0YIZDc
aC8JJXcWO5/Q06sTxfBR24+0o+RvLq51MOaN4P14Ou7RE/oBz3qzKNakD2FSAwe2
VJIZB4dpnrIgyiQBnFoYH3UWNbiavubEMg6spvew/tibGDL9+OcyqJ3jzlX2M+Vn
Ze+cKI5t+0mzF4GTWkDrDlm3K6FjZ/gfG9IEbknCUWmkoIQultavtxklgy1z8D8+
5mHD+Qo+GpKIGjsu8YM5C89kF/2ggPlnYa05+9iIygdzuCngRGeC+80Y7rdlwOfr
WAbg4ALl4K6NiFtwIYv9PAp1IoXcjeAp0viMrX1DTb4U4BWFgMEhPV9ARW0GOq2/
6T7EdwDKdSJduam4aj7jnHJ7XyKZw2VTkcoI7rT/EU0+n4qnZ+gnAZ9JvxTWF6vD
jw2iGR98O3PQGswxA1kGY4l97n9zS2WHYd0jj1BvYa3yu8kBkwf7YuI10Wr/Q4m5
ECTOLm0ZiTpvvmDRcSv7xHefc0Cx7vXeelVsJTvYy5nwWQRURRTcXNZ3n3VE/tQb
V/ni+5OYljP2GJ2FB+1SxS27xf9tWri6ytMK06sNn0WomY2RU/lI2s7n2u2Xcdrv
dgZ3ozs7iVZyGjm0p+NpR8hze9psgg26BqgWRxiFltDVSAC4eY74uV8aV3Fjx6ja
xEMQX2HoDE0V3sd8xB55f9kpcC87LOMTuMGDWYLfNdB2n2iKF7VGplu/jOTuB7jx
yTmp+PwkF0DkR4EUpvbOQ1pGA7GovjWRGN7webIN2g5wItjF0nWh1AbXY5p58yuD
hRLzCMYtMEyh/k5tI8SEUjRIeuyuTTX95LzKxdBqkXgOPJqMEYVNBjk/W4C149l/
os7Zg7nJeZPe8YSEbwu3BTfwMUS/9nWV4brqmN6C/Dr2xU5hqUm3lITxa8Wg2vHD
jYLYvPGvy5biftTFxcXZo53cg66YExfj7hFo+5JRxvBz16Z8uJhZHr5VfqxR7PN/
JxtU+Upr3lQieXn+B/LyU93sJfO8hIdpeaO5MdlYvQydUsP0V1a0n59fed6Ra85l
TAfX6/5miEqVwB3gBT4mv05NZuLSkCfcsClIoKZPkckiWrfvPWxBM6YT86Sik9vR
BaVyzmarXewWwv13jkuR4pDvc2dGyZPPZS+hH7DbBzNMO2POmQpXnVeBmtxUM/qA
20uxPjtq1Ift7v7FjTDvB5lRNv/pIFSV6ZRLz+cCqotHC0vv0e7dD4l1UceotrYG
kDqjSL5MPPgxpQ2Rzy6WDFZ0+Jfpe6mYpGkGm6xVYOQRiEJaDXFsn1q1RJ0auvHH
H8w7Eb2jxcuoCnY+7GqT7olliS/7/bEejH65j3jSAYUA8hHGytq6pfPM6alXkyBE
pxCK3oMs5rrAlhP8yykZsWtOnL9VlKWtariVhSlf8YVJOubFRSQBjH43TQqM0+LU
AzzPNcIKUR0inthLPb77uo6HtByMFHg5EQf6kp9WvCVIO//gjBZn9rlkP+HlaDMD
uKlXeuF1aqpIxiS3f8GaP6ndg1jEwT3GKt4MEWGQzYRS6PcSmGrtvUvKGZLsfylD
dHHmqrF/UFskpqPM+vTdnJOGWp6XuKMyv9afJCt33yISx2RuDfO/30SLAHur0Rcq
BXw4QkAFnqEpEIn6bQvOCt8i5T5in9eQJ8RmWwqkEENHBmN6rbfK8Oy8h04X575V
othmGHtwXuFKrG4J44JdB49/p/19tVoz1iTixmX1AbXWtNlTOdrrjtjDMIP0egqY
dPp/BAsX9qCLbh5dtDUQHLCc3KkqhYnjnJjHNCiSapTi9HJY0gWCaoO6z0wM2spL
/e/shyt7bwtQR21iPmaAQ+Lk05YG5gc1Gwg1QtSVcepQCH0YHjKoxSPH6fdquE1w
E9lCaO9Ew8j2te47OArX9Uav3OCvSsXNt+pYC9BnRXzWl1uAY0LroOSVD2f8VdFP
8fiPTwmpNhdf61ExpxtdbvjFvAA3UT6BVgn0V1NuwagrYX+6c3AIMe7+KcUsIPQk
zRFc0M8ilE9ACcrVk2xsGDx7AfoRut+cig95IVIBC2u7c8tpv8pLgRyskmt+0pfc
fCHft4gnWom8SO44CR+Czw7x1ZgcJtZ12cqFZem5xDcpTX3Zl4ymTViqncfzZQ6q
akGKlcuuRKTkbbhrFXqxfElunI3cy9N/ESANETnl75b3ztvKjVaPVKSX/GUeBp7T
UpqzXw5P0FQMn9dE7lcX1Nyz6NTtLgIaxLEZnhra6KbdeTz4djFbPAZMMZWqFapS
6ArJ7UNKcxbpcRTL7WyT54vhT0Q8ht1/ViMllcUtRjEK3JsYknlZEhFFc6uHqOrQ
kDPYNwl+Xq9cMIGd0PsZvbMR3fVEAdySNCfV/aMnNLCYpFyvqPMOrLdnJ2nWQtSD
HyMn/0MbS+O/6NTxLplYXRXZg2F+kxwFihX75THPOrWugGU4uo3E52OnXOwuTHYj
zlULgtD8NMdR9IgmMqnd+uUcaJHZqkKFdSDlujiGYVn21BYbe2RFsSwhGaIZUe0F
ees6eOPq2zXarurnGB8S7etqksQuEM+VaCJTPFCw/Ytiv5+Xm6pfiKQlTXB3/q3h
wUGox6rTEh+2o8vZ03H3hLITvcHhzhgSTAtDt2q1AivU26qFDd/VY0iEwBLAcspt
/AVTZyRn2CcHDgdADEiTXKIQbS62QZc1sk2Sh8TV2XteEqrg52CDBP2sKld1xpPS
HVomiJCh05b0rF5n5vtynqCvY1qdToEiuHTWQ2CQ6zZRS0zwjWd6K/eDZ4n/Xa7j
gJGUejxxOELpqqk2jvpJz1D+W6yK/LbUqAZbdFCyx6298hP24l7imXQZRAuu0RMI
3jd/rYz6lltp53J+OO6xmGCJ03yHopJYVaX6M2qpRghzcnvq1xiZOytH+Bth/cTK
vt4DQCu+J/p9yKUGB4bth1G7d+BAPBsFLMiTWGYn0aKs1Qh2DtY7B0QCC+fcpQEk
F3eW2ognfGN54B9/UpRXLaTTggOgkZqZPNkoDgbaN6ux24sPpRuyCDSJ+KW4eVkA
yyCTO+mNOrtGGo3KqKLpK+LQ+RMsof3lpLm+BKefjRIIVNTS9Mbmppo/BF1P3ygA
oOhScffhD6YX4me1Rq2DkFq5j5AFoJGf7XpyBZwrVZFx9skYvEE5fiuF8Ogg2Txr
bKBLrkyBqGaaktV0JIbfPIywVMxi7owbHVS84s65GYH1DXeiw43Q3MuwOX7fpIF8
DywtAO3NyLyTJ7ZDB9x77A/K75tH8RTID1Axz0+6aOIox5+JxjU+lhEG6obbrcVF
Du79QgCyAXqefy4PzQVcGdsUU5gFWgBcpKD4bTih6gGRJwZ/T/+uoAhCsym/CUqm
tXYAi2UEzXfxwJbKXr/Q4pVt3uCvkfuuuTv/uRPRza/tsiqrsrnkyWqa71cJRiyL
OL2uBmRfB9q+1CItzzZRBbdjPLHOOiz8lmBUo50Yzxa3AW0zMYYxRJZ10ANqdTUA
2hSdi00SXvCf7+jrMtgvOCGEEVUF2oM8sD8r0e1R2CxbGqo+taihzw0L+vqIHS5q
V1druid2BzZTstjS3M2ZDUmu6CPwlcv6xere8E9IVfrgmJAytyvCPc9SuWwLa9IO
rg07hOW4BAi4O5e4+M0zx3E8YKp4AzpNzt3PipI7Eky4d74pGYAhoGHGSgqXM5R0
RevW00SFul06JVjQiYo5SBFh82v0+NbP9RV+Z/wWcQC9rbrQu+O2j2Q+sOmCOEi1
dmmqD6mWpBLCBffDmNysY64dsb8UTu6AV3+YhjSQ7gGzRNPjUYMn9WJChq9TiOo2
D/mm8FPD2I2MddwTbfZ1l6Z1AFPWqSwZ3CyQieSa+CkPOmkAK44mw6gvstlaetbf
XE7BlGQt6/OiTAjIytqPnbPScpLi/T9BwoOjBuLOiXocLuZ+5BH0VUF+P9SWg93f
Asz6wY9B3HWlViNFL41QyWfBaVk0lhnFzb2F+q+FHHTpQFljs47SXpcXBPN1INTS
c+br/0K5wiCJ8lzJ4fmgWOw2dO2sfdCqZOVdxUQcn/p+MElo4FxSUO02WPsSX5V5
IKrC8DTPTIlXZFFC0qM2oKrtCULduczP1eNPSR/gFi3unVzrsN8BQ9cjObtmkp+q
EJL2xvM0yw/uPQaOt3vMretB/oEfRjbBhq7fTBuyf+HWXV+xQ08HeyU9gASO+JqH
puvNPaFAvMQhGEssg/+ly3fxgTDuxErhrhPLP2tTR0QS2F11wMIVbw5rw8Ce9UE2
N/3+iHe5MP0YBWtT4Al3H56iMukPgx9xAK9d6MVEP54Wx1Kl0XzWogwV39h0mITp
N0JhwBRvR+gWHLSbbZiMysIKu4XjKEBgfX7xMdubwnl6o103KzHRkV1fTM14KLAs
E1idz0WAhN0lb7Wgnnuu4bajrkCQL5FjecXpdBsmkS3jEwBikvLVz4mSKSWxulAK
N/934McAObBnFNlCJMLeeZmEpvdVzr3BkrENiR+RLOBKQyo/4QLkgbP0VaffWKMB
QTyjlEe4nTRg79rv+keVjnifwE3K4otJYPDBgjLQNEpgr0jaPeO7Vhby0Dh4wtYk
iJm1VMTe45engUe6iLkJ+N9x1QDQ38+Due7VYu11dt98IH+sYweTlDkN8/XBm1J0
HbMmE1BJJxWR/EJi/++mY2ZTARSIspveSjIuKmW5UMFL0XCGiO/1Are5a7XbqMe8
dkko14gHXDmExJOeLway64P+RT+WB0MLPboIWhgnPDQ7yKi37ZSS80OmFtOY/oWC
+C1abDHG6ie0flB3nl3Poku0qLuINgo7AP3LhbW08RImCPcostRWaILKi1HweVMX
D1PbZzYfuG0K8m323+mcW8gEG3odcKaMtSqoqycG5L3/e9L+tR9WiOwL8dYoMIK+
gbYHiw3DElw2CewSffLLY/PVqUaEP3EpHDPEvWMX6UlLE7MFhP9guC62ukuz6tyO
W4Rg4tKqufRvZRv6g5dlVR4EXoFJNat4ghj8B0WEREk+Okeno165pxD4t6XJbZJw
gT78topSFgquF+UksSqJCDxqF4HYEfWsEaHUTyk3KZgE0IASdO75S/C7mZuvvZ6s
0kDdAXwNxt81m9VWoaB6EE0hzN99F3s0uUGMOQIyRp8BjmP2AurZMO0j4gXPHifQ
WqHBSJWqxt2sODDEMc8xYisca2Sow2EYLLc4w+YFBNL/y/ZIo07BFBaJjIRNQRIk
D/dA2xqA0g3UL9wdDY0p2pFo0jBCBFqHxxot+epO+MPMsaIpqCD64X0X3LgwjMFt
2H5O3iHlIbR0zUm53jsuFSk960C6grZLIT5N85nt9wqDa+uXllYmBZ0eY32I7eM/
QRm2vZAPEZ9WHBdR361xZYeyGxEJT374KbNuqe8UWBdfd6NgqihRvuxRpbwEY/Ov
97nSMjTL4OHm/2jys4zHj0vo2FcWGURb7/tbQsCNwQz3AmQnkBkgqGrNOItqtEmI
nIlNeVM9cQ4GV3BCZ8n8vp/veLt41uofod9/zm7NAOAiI3UNa3OnUvJE4nHyA5m0
zOsUJw6EkB7byLBC5utqWXLXPUvjVls5wUsEy4U8b2kE4Lq5qChdXWNbIPnB0+Rt
6LHOzWNUNbVaogi3rxo35wvht955OWNCojHdiksVidtn1+rPtWfA291VXWHgdvH0
IdEyCNowaJCs2M5mRfJVrbSF91tS/gL3ni3aC1VwHNOxmDnTNZFdNjojgJPpVN7D
q4IKmJL2g2s24pOiqZD8T/7G3f5/kRZ7972smE1c+iWJWIgkDwVWOTZaDgRCt32O
nPHJZHGFZd5Vnj2HFUdz5K6VodZ43hHMPnkmIdol6NXLL5dVKN5BPIOeWtXpanEp
VLDYzPnRy3d739mQGvg6UDghFbv+ICHayuAWRMM1IYIuIHxwwTzrfw4CoVJ6rOeA
0LOB3Z/aOsKIjMCMI+3naa0QZGepEZGQ80XaCDlW6iqgSLXNyB1lX2FqdBEl/lYr
iGpXnMOfDHeQKt2UL9wCSePO9lojjfVh/yzA6dVnOGQI4gkILRQChqUMkFemmIIZ
9T/9qAqEKJfWoGDE3WQHB/KgiK+ArwOU6Y4k8KSDKgGYjeFCcGzTDKvMQ+QaV9Y1
k0E0l5SW+wLb4oY1g3sqNpUblhd/3J+q0Jb9jmD9HZ6oSF+mmUxHODRpw5yeFyQF
u2GwEbEWY9/srLWDvJYq9m9kkpcLQdTi3yUyMfmdZLsYkQKiFsKzaYvyR2rbCIOU
i872WSS0d9F8hOUvzluJtzC5t1IvObItFI8OQffkNYiVw9OB67CCS3Hvs5nMxdCL
2yLRwEeW+mYOwwlKPO8+UWQdeRsIeY6jT2BEh4zAU3E3L0HnoIEReaGO1PK2SN6Q
FZdc5fk9nxyBuWZnuLRPbUPyZYqV1lOK4BhTKp6Cx74qVTBtUuiS//FQIK3f3knR
iwi042EtnMiaa5O/xDmVB6SVXdwjNlkCFJh9pwId/rx2UT7VY01Q9xu6rhrP/8XH
wSaltlz/9DE8KmG5PHQm8ZE8E9lSOWgQ8LKYjFIVjUEAWw2FkhLAdR2LOPm20UDK
Ou4LfT6suLON9e0gpKni3P6V3IX1MoX+pM5F6U1Oym2V5p7j091u5phGmadGQf+5
GSpQDBOnzU8G8SAZ6YNaBOgxz18xg/u58RMWGUqXYhawtusARD1GntM8qlJBQXFs
WCExU0dcYJieZYwk9Vz9W5R52pvHEZLb2EEzcKuCZysrCxTJIwrhImuhnP6qf4aO
hEtbBYyD74cGobmh/Ar6T493LJdd8iJPDAqxHfCfVaazz92B5BKHfw/dFq/I+8ON
nukmpPML+AvBXL5fxEGQ5Rt8e4qz5CwsGiNluLcmaS4NVROY/6V/QLkK4tj5rijw
N9LPk6gQ6NS1qiK02dDE0ATClOecUAU3TrspDc7JTo9wArN9SfThNFrw3eUqZbjm
/421Kw1HKDbdlcccK9fDJGRRs2bSA0ATo1xXmqJerPea2HUQHnjbo6zVtQbJWSYx
O/v+WqT1X6kEXrLUymRw36uqmS6ZRwbSyqA67CS+irGWagFaxmHbmHht5TaZOnWd
3zvsGFnY6iuiUYEOT8xx6Yqf6YhKg0nzhxcP/y+6rCRBBQJ6T3jlTVntUG5qA9u9
hl1t5fqxGq/uEYA8CUwoFsp4jrw3umcNYSbkomWi+J8KJhMDmM459n1AgBtpxXlf
Ph0jZ+DAITkaehCGFJnbuQzA73AOJ4VSEIsmNTyqXs/gOheWZfWaqH7wcvDqv+o2
hkLiog1WXau2wgVG/EdK7aiaXuXB2Ae4ipcXH29dLOY4Up4HE2vqoOdgaGMIAu3H
qMHLKvBNYQClIc3uDCEMkB0npy9FXKkKUkHl4AcyQqe6PuCV/VW093Dgd2EU48mI
4jx6ybiHT1RUrWUp/qs9SOrs4Ot2d5vwbNaKu7xaMf5MAwwrbU7gmX6C+jRCjWn6
rJL1bjv5GvPexutMrDALBCyHNYBHC5o6j8SLp6JcDFlwFc2s7afT28L50IM+JFJw
WT8YLNeM6FWrUa2QpnqPRBUheQGbyz0l7TcDJ3+ciOfjD+O7QNymLj54GPf/V/Gp
WEc75bWAkfA3dRnrZb43IyIZ4KgfKyZb0n0VikNcjtwgIWRSW/H/awEb5yugGTZD
nheg7thG/KVoULIOmNZM6l7kmiaMxDRJCn9H6emURqs7Yv8yijaEHsD2k2n+JKYn
IMG69ImRlStBYxOEHoNDEycUjqVsRge5SI1y3d3LMatsSAOS/FuZHaOm5sJJA+6Y
J0vSqZTR8XRxFIiond0VpV7qdpz3d2HjgOmxdY99llPj3HHtvpRkVYKBi2kg7DF5
RisbOa03KArQSQON8/aHJq73+ieaw4RL0XhKVfEk9V+qo/nD9ygrQGpjl+t0fxiH
RzPJmi9JeybTAdlhFlQWEVxgxttstAMJcBzjqQNqW1Hq8g5n12llopFtFAgEfUwg
luNnW1THaVxqb5hEFyNUQMxyhfuTizJjKn48q/tsQxeKwzOk4vXfdGJGHrH9Iknl
lYfxv3XAoslHBWWAqt5ktz9PD6lwWm8NBvwTa5ENK4l7b4QFu/NnPhSCHbXFVMQF
hY+ESiA24ysZtJcdB4v9zKKqbU9CGcjBnzzb1iugwj5hSRpCTze4FRSCZGbWKBqd
Hgpoju41CminWNKhEyMTGTqLoawytHj76wMWzDErvld4eknBISkEFwA/1Me9LuTl
EkriU5elkuiWHNNgLQK6hdV0CzFh4VXn3UuBb2KfmzqkcXeI1Q6PtWzt/BYDRZTH
+e7xm5XOvFHq05ygEQLiS5QVh2G1v2HdUl+1rmE0W8iI9jG42PCT1mysgwF5yden
svAe61Z5kRi9gHoRCOljZCfhxf0ZE/7kv9aKVdSOJRo4qjZ0h7DeNPvAR5W8MrOj
tJ5UPDaYl9ENT/YcJweEshasyG2jeDpCm1Zg3Ino577JTCtEhrxhJ/HLND4NxvgJ
vc84/GvmRwU0bcyL+cxQVJLvk5ZxyPNFnHa2lPrzoGiVi4DP1ozWXHFe07Hm0kKq
4AmV3DWdVUG4LGI48NmR5V80RpB3i3JCz/5o1R1YaD9yFZT+zfjf5p7QlC+gT5a4
BWIRs4hKISL/BI6tNBXLWX59FKgEdDrIlye9wb4RZGpWPW3X05UYD9e8TFZpM9O+
wdqXJrZLThqmWb+h4RS6YrRCX1E+OYLAfOjGKr8Edv8MxC+FMvawvRx99UBUPKMz
xO0COrFoGSiwFDwml2qiasefyFHtyIPnoj90PPSish3BRwq0D36RuhVn9bTRzWkX
R1KRmlG41L8EizpqhnunOt2oBogV3gZrMSdUE8Kzp5PT60HdDPQkdK66RCM52s7Y
lGzSK9JQjZx7qfHk+azuITIPZKS9pUTtmdqvlSDG5Or0HXW3TtfoxZAVliO1jK/4
/0N/UiE7k1Q4/rNBjEL1GrbfzzxeKMRayo++nwD/6xqwcbPtiSUiF71MePamCGtP
0RtNZseA8DNAvLNyJnUmzMrG6bFW9PeWw4SToJtzYpQwShjO6xCLDQYsVwww0L42
kuWPl+DdgHfN+g+QfwXxXodM+CZ4EXCPhW/PGR5Q1+4QYYiQhXZbNnu5KjdFr28q
UQbPvDQBDHVAhIFe9GVzLQxBSL+kVkZuQ1IF+vzRSNynplJdWroQfZraAv/nSf1x
ufmFn+6HgBgNO5ancdI7r5W1dmnkTYAFeqIv+bYwDr9pm4uKl/8Ea9Xd2aVDZTwy
0SY42hgEokc3j4HJ3p6px30njGrr8FqjtJ42A3lFe06ZCL2JDG+SKVW+DubNEuV0
uzWh5KZXQniIGEeUAl5qtRUlY740VFFvF6gj7snC/cz4Ewi1uJBA0GAdR0nHsLrD
oEIykGCzf1pp9OqK9MTWaL8MngLJvbWJraidFm9msDySVpWEXiFKC3grrweLedSa
1SYz2aH7oZ2JlOqqnN3fmR3XjJd8xAIXFDtCC6aO4+lMWpTvUarvneYBmQlG9Bqw
xySaYHhy2lDPLW9KBY/UE33JlixgS+2gzWgdZgF7NkGy3If3ZpARjeLGANxbSL2a
l7sh9Elkt5MY/gibfDge6ha3SEZ6BNglfKvxSDBV0DcMDlFjTrrbR9Zn0RtJtUxI
ya3jZutUsa7vudqPqFbDNHAFKPD2LCvt/YpgAFjIAIJTVh60qFnNXVBkdbxWbOLm
u6dK3jf97CR24TrUKPMeEnd6IYHg6vtydKDw2YCz6xS0G7Ae0KfMizqVlNaru88m
LLq7zLJ1bzKpbGOmNrv7uboA2Z34oFGr9+tXYBVFNcMePhbntillrFiRZ/cqmzte
8zeoatp6G7c1URLoWQtFPpS1t0JPinSdsT4tyBWZSZjbT67NMB0DWk3NGUk+r1ui
10qob2dvNDrSBxQgtgwZYX90sUHvxTz4XHT4iZ+CzEcL+q0UgXcMx/Raan1uUCnc
A4OdQPHYwnnv2DjAz5PoKXngmU8uuT31L2F6zhCCYGV5AHZA5QHLB42mr1OVfNbu
50rMttErF6ZL4c5m0AmSAH9CfqnoJDTcPh33odVnAKzeko06Iq+L1/ArPkuuA/0Z
4vah4fKkWvDxL997sYUm+YJpntQwpUWDR8FWSZHDUH5SghOnslYyNiaq39zIgI/G
yZRLjrhkcxrYwg4j7Zk1BAZIflzz6yYPFOh6yihFWn3tB6wWotIgT98UzZ6Hczhk
c3Z7/4U9Pb7YPsRMWiYpYyv64ON7Dx7Q+7NMxi0Q/l+Km5s4+Drr55g54SBkzciC
Dn1MDia0GAz9VMBhXE4YN3rEU//1gbQfVq5op/JjWlU7cFqo9NgIdewjXw6z/EL4
KNX/G4wWtFuy8Rt/bqAyzsVGzWj/bQ/Sa8QC2rjMZ6D74VyYdhj1GZsWPrZ+DcR9
cTrqHsxq+5FeYKxgOpUeJnFA3sVmzH3sFCUhQGpn4skEnS+UX8kWfi1Nv7etTAA0
Nt6da6H65OXFIzGMF7EE0Rm0tANNFVyTW9pTV5d0UjbLsPzu2G4kLIZ4rSXhZ4IU
Tk1BMU6ce5B4G9P3cRd90gtEidyXN4kqk5xqUrH5Tah3bI3BJQo179aFPXGejioo
UPfDjbnHcHVL1MXi+wgrh2M0gK9tUNDP7TCZS9MT/WRFaU17vSvnpfpOD3gmZ/Ao
vI66a83fpTqf4mgucYyxNcX6gEMvF4RCwlJNQ3ed6Jfr4c6PNdMirYTtSbdCi9zw
4ZiBC5/i0DIqfLc5kjAVkgzM8A7doiyV4pbnZ14xKz2rXePCqNwoc1dh35MQNO3E
Web4MZaBgBersaYNcjQPc+I5YpBoeNRC2B8uHFRaHORmNfmAa4ekg/3F7+khy+ju
oCa8WmD3YPZPbKj6WewrHiO/vqRd28haYmRW/SMo+fsEI8MhIUOD90moX0VmtVxg
qv89i+7owfRZ3+NpCJ08fKiNJIBT18ietYXBVMMT1ehXOLKvetM4TJI4FVvzOr54
hj9G8My0bmFG2mMBs0ly6dES0Hg1sJTXIvC9D6V0/WM=
`pragma protect end_protected
