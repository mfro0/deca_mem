// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:00 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PLgNm4cNCGzfkDRYaul3AoJadVp3huUQ8jvPgFtpDiFYA+mxtcmXoeBiwPwQ/xNS
7umbVfmW9wk53x2NF0/Ua0EwxAKFrsGKb67PWxBVcYP9qtyJzRQne+vnlcKRs8+8
6Y82YbW8BkGVx1h8Co2zBttvsJbCYorPRz241pzwHwU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 56688)
j3biROXhuDFYIaUN3WTgi//VIJjkaTsT1/cXXlFfI0YG+1qb1wJGlXjW6DLgZ3K4
juF9SB6C+LAsw81BNJj5IMdI9C//NZgAePuCuPRJEorjuwuQvJHuhg7wCiSnj+iJ
eCNN5Q0q0yYxWEIJwJ2U0Zj2FAy8hLdVxpUyYJVDK3VtMTg23UaKJsG6ghEPxOjj
rziELQuIydKdYqYhq/v3HAOLSe1xTE62kUoCDgjLNUHGhR0AuEjpEDQFoBNuo6/0
dM9M7aXt+1r/5b979Cge0d4q677zUMchukwsoh6qG9UjKVo6cjsL1cn7LMQrBMp+
neb+lfXNFjgF+nLqM4vc8ysKiuC+8lzTt8Tq5RAKzOk71OW4xMtY0MTLnJ6gvUiD
W+HFEStZnP1bknIbwaAZ4n4xlpFIDu9Gb8Nr/YT8IzAm6UbqaqaeRhg03RF9E5pO
/hnFaZIztFrI6VEugfNkcFM4/FZEq11GkdBEs8LNyj9tpq/eSDaUNr8aXqC76ec1
hVa4E5c3LLgmltUELVjO00TfLtiFPtHKQHatAmNGPYXFRgmK9S4uczAJMj2HpE4A
+3szerKCXWF7Y/ALtfQzmDeXFSxb2xNGsxjwJz/y4wGCmc2A+OxGt5Gq6+fzPPR/
UYARoYfzoxZapD5BA8/e5M63R6U7cZ50l4ayzppogAFYIz8fizCVKODMuOGkMEy8
nt1dFpivE5cz5ycXCrv9154sXvG0n5DW5wd7kmAmr7e659HSfAMi+DoE88cLcjEW
pVw2p1WoFzJ995EQhvp710iHNmbzCN4ux6sulSQksQCeQSKMTrFMMToCjVT9gN5T
xnlm1gjPtTaAX+hdy1UCcmjoYCTAa2jUS6FvnY4+Sv2efiqp/JQrU8E7vom3nMv5
gKhE1+q/pDejRpZZWMpgaNuJUaA0Y9cTWJRXcxNwihUUKrLJ2OcvL+xfHrFoD7qy
uKFp5gXSxLgU7wCrU6y1DJbtoFkObPtx9/wFnsGFFc2Sk5uLAAu1y8YULnLV2r6A
50HGuevtskINkY1pYWWnloU2wnZVPB+d08nd/wq+NVR8sURn9k6Pnft3rVqCgWd4
lysSVg2mxVotFgL/hUb6SZTWXN9n2d/lc3y0tG7OaZXFBs7rny/iPK+d6n04zW+v
OLE9+hMHLP1pDOEuLnSoWRzeS1+HSEhudcScChwVo2aK32J+/eg5iP5GjAn7YEfC
m1LEkREEo5UE+qRSgGPyIg/w+Lk7KKuXX3t+DehseuFenMT8iRT3Hu4IyrswKZQ8
P1sAtdU/UkL0YMjDj2f97pfVy5piwVYr/cAReV7PyaZJ29Lv3V9JrkeHOWnUUCzP
/falQqSD5sb5dD2ZJAnSFzH+8mX1N7zPChS2jB+bghZ99WKPzhrGJdD9xlVxmFFQ
ecWjkyhXYwgaYGurTsd3pbkpsd080e/ARow/ebEwx873kAi8pyHfhRVZ607up3di
V5RECpTZNzvYo0dA4TrStyR+kCFlC1qbl0BM8od/tM3tjRhKc1x83eRaHWhVuApc
H5kTwLhXnu1hAI5STFf/3ZGesmFtkiVk/ZYhPuRynhXRhGG/dDcYDpYbX9ck8xYs
4+ZQdjYkE7Xj59+R8Xn0LPOkzR5nXrgNCp6kfLr0+WHf350YwJtFm1b3f6UEGz0b
t3EIS24TgaKwENl8TnHasYyOUQaOeoR9/shwp05d+6ff18tUkN1s1TrxzWGR2xis
NpCPHybCEwV31EMMNh9N97wUpgDFk7XB3Ea5Xr/02vN+lYPjhRXeh1t5gTg/81Zx
sQpGLwxz9OVXH02M43uP3DB43Qzbxh/7rddJwviHiP2hh4pTonl6frxg2fEotOEG
7c4wBRQXSS+8+oedL62y1LLVE/yoNG2zlZp0UrIkSsGT7/PAt0NM1mHBjCCgM9bL
IgMxFwt55VC7ClrxMK1WmTCFOC+ZlwekGcPPl6cQ3qvhsDX5CBvpDtC0qzVx7Sc2
FFyqJ+givc+OVkHGa0WCkGaXC0nqPFBWpFhSHvQ3gQKn5I3LcI7VCNJK5Mw5Erb1
nBg9EBERqWponnHiNNsymhmFZR8k1bM8RwznKFZs9EFJuVbk7vMB2HiWg4foY1tI
jUnf+/DTF9sDX9Ql1VoeoyLA2NHWmF7hi+Je8X4L1G++IqA1k2qpCJsDtuaQlJ4f
W5iOlLM6sdX+JntqQak2gGsEI50k/rG4gtvQ4IR7VA/Yebqou5EjjEoNxXwh+unD
axskssVGvLqeXeFMGBCQjKH/u6gt182+bO1KLFD23/6nGudJWvR4UDnUBhfXBcyL
oHPbOWSRVAeFXZP4bXfAJowl7fcB/IehdcN3JJrO5EduZmd5CyZTk0rXbZW8TfoX
4ViJgIXOhyItZ6y1xro/rkeNERFTgtSYt+LU5aPiAoBT0MSWcsEA9aaEyGIaWdWc
tby5As2Zy02K0sSXeR44sZX5wIheIA3ewawqTp4T7yLv8USDQbg896odTsgdgYY7
O6GqfS1nR0yYNm1rZSm0NggYW81Jz5lbYtlAdmutMWUTJsdZrD+uW9RwYoVzIMNi
LRSHv2Nt+ScQM2PATJKVt5hvFEIfL/ui7pLB1NFRBVIErcw0Mj485/PwE4QT7G6e
N1rTFe73OajBLg3h8fcYC7Zv+KlDKkMlNJBL9j8m6E911LRIGa4gGRsIDbS2a0WW
DlcWoY3o2LwJafh9n4gJX3rKNmiWyTh7FeZ8UgKlRc7jbqbZzbV8cmTUUJN2ZiuE
AWFGGGLGv0l5RSnRM2zsAuJd+4j6UleW2MDfnE8ZR5pQOd9LfgCBYvAhaDMtXn7n
ZnmWD6c24ZQQsjDzvLRchJq9oKkJm5q7crgP8vYAPvk476/3paknh9cg0tDHn9Ln
6TSwDBVNclgbpAAu/q+3ocgLdaBPIZa/14J0C6lC5Gp/XEZg8wrLaE9t0kMrH687
M/wbci0HzyZmky+usGwh3EQEbQiBHjcz87RUEOvB5IrdlNCA6+TyP6qCtCTa6TKL
m1634moEj2rpamgif3pv0UOoo7ytABC1jzGFO9zStwnn3s9C6cDTSY04GWxvQ2Um
c1379s6MLoK/djzpEYWSgfPcTITYcMC2nXX2LNun8uNhyjazkpHPieiX4pQFufRy
fT3Et28FJfIEP6Tniy3JQeTf+CxBR+fhTLcd9NzV2BfB2iU8koSQ2lJchVndQpEN
vT0wD9714fBHC6L/faRJB/QhyxQMscJ15WNqYNLwcCT50RdbhIo2O6wMkf67usgz
2if6txesdaOTskbWgqCOpbHLz80D/qgSbQKoWrg/IR4lmlLVW3jJkmK6D3QsWTtt
R8K9nYmiIrEpk36zUIdtFhU/lzno1QYJg7A4DuspID9AYNKC5prpt40JBfUXMps8
NSO6ElISdTnKTWMFtLua4ey2/3TZ2Lefb1dPsszzjTbfPNIEXan0RllqnGqF1JVS
p1UznDDAI7jX48fxvss5dD2pZ066fJMpbNE4mca2x5bxvffd1AaxGNMytVDmyiMk
Vs4GP7OFRDPCF+j3oPiesAWUZZkNBYk84R+bDFZM8QRsiXg9sPKWRmRmDXGf9yvt
Ls4uPgMZGGUSPLNNaporawBGP0LI96qV1Al/Al+l+Rd37xRwy6PuCJ+U9pHRtMqW
XEkVAMSHW5gJqIB6qQdaTEpGkZOskk0OOC4p7iFPulLzORLX5kzgYMdEkqoWZLzK
f3DWo2wxyGW+EcHSirFv6ZHawrhr3h/Jy+gu13SmR9MpNoVzSvwCiSkOAf67lamX
2WocoZF5KF21/CYwQNuA0U81eStynA83D097f8RbzT0Iq5WFi4FwKqUIPMvhULDQ
LHeo6N7fZC33GcradafaQ6LKcj8i8h5LMForWZks1QbS5my2qIlBFehlkQrwgaAM
iafg8Xb0Z1Uu6llueAeX4YTX1lnW4NHVXrDYmtnwtsWvrPQJ1vUDTGpU9lP3eJnZ
cpnKgIjyYD4TerAGyqxFWSthRUprz1gtRjD4fjo49ICKrzY3hA3ysh1NaJB/Pnje
gyjrMnU/sVAgOuuHq3OmR/RzEO6ZnQD5YfEMrbZQCbQoLNnCTeS6rFvAG92vipAh
BBwKFP31jhzz7UIZbGwoRCAFYXUjKosTpV97Wnu2yVZxPsWVxTVaQ4aN3ExS/Vyd
GHzQmn3Y1sL0jm1ZamTX41KDD8gTWclQbEVDCr/PuWVN9b6ot5NwOCzuMjP4DNQQ
E9KHoajz4VJMgWYOx959qlGXEi2fAqK8mao4x8lec/aDUS4YhWfrDAdSaT9j6akJ
7QKIrn8thaTVvby2elBzG+JPxvKH7BUR86hPgI7Szhi+rbPadBoYPAgGvY9ztNQY
zMx8OV5yi7t8R1a50KKi/1PGDOtIKI59c73Y0tVDMxce55Z6Y4OD360VnmSlMLTT
3twihUrh187QM78Hwz7eLMUs0P1x4MbwqtMj4Ua3br8XjjEjvVblminiADh0Iyxu
Y3uVipEV5fgfo/JXpN9sARO7SnmwLdADmSEPI1PPLOFLU5uIevVsimJIc+hvdVvg
HSVxvHY5mGlwQx+uQxETkN+dI5PFVzdKEhkf06YgPvJUlGOvwxcV8BvNHNqqDucy
n+FVrPTXLwkgha0X7ei3NmoVthWQvCginr2K6P23YEmgEGAXeuYXY3Mb+Ab2Q3hm
d+TuqzeGjrRoXCLZCc+n3mFfQ0b/ohUlnvdsLzZ3Wt0AXcEfAj4JlNLTO95m5w+2
KEgaBNa6fmSCNHq0QAeqxsvi6mhm11xhO/r3fNm1YJXJC+AklZNjPyp9T+VL8YQq
t0trlFkVl39Og0w/PokWjMHh30qa9Hc/3AbLttqp7BREKpiFgPATveab7RiQpcdN
pJ9WOHLGO3UHNnQjfhH/oCuBDcmv1FF2LIWyonDpkM8txb9Ax8ZLYX20FQGfsiN8
YIhQKEhTHDxCTh160c1Dl2fK1wBjDGnW/bVnms8jEJA1id1pbN/msm86HHU49Ze8
d5/B/deFjhGbiDvP4ZaKbXqPLLK9jgaZsn5D5Xa4xr11GPCuUZgx1G/4wPV/ZSTd
dfoKQQ8hDoXMih/AIzKgyI5/Npk0KjmujEtxW7vKkDOYikqU/XACxu4p1+DqTMdc
fqOPEWlWVjm1nvGRoB7TdqUitmU2rvUIk8AWFIRh/rkIP90R013yiVbSk45ktk7M
M+41g60GyPx+qmTCdOPKi6whH9OOsUW3BHOyuO3BVpkVYhjiuvoH7hn3RTKrUEt8
d+hWsdzl0zydHLQwSH7a6SpwQFywgBBEzAulckboF53z4fG0zSKkrrz2eOPA85B1
yFWXzxI0RlM6oNtbQ9KRfflcV1mgFTk0VgA5LTy/IKArUPTXhSYGvzgvmygghVVO
LnN7zBiFcG6XTZTHHODnb1nf5dNucPr1OKawgqja92e6Wwk2JAdK5xQ1FwnQNZJW
xBCvU635frVfK9xqNlBk4HSvlDBBLApJxy0qzPwrFRsvtYqyEThQ8EGQae+NXvBC
9Jf3F0bR3AntX0y+eCq0HTM9pk3SvJRP/SWMOCKiRF6XGHMBl9ijwVdbuGebOi64
JwBgJMBFQUiSNl6mN3VygTskyDpA6Ip6C0fXUChX16/wHxYj359DvGCmlCXFtcY9
r0kDusVy4Gkc7eBYDDpNFCe467ftQsyfLBhhkW4hiWvllkUXugKKW1R5YfDCBRWi
7ikCXiSBObtWk37wcNsO1Bq3Jzloz3nsZJQUuGFMoGlTy0gJpoXGPT4rJFGMQZ7/
aaU7VtzVzVkoj2s0sJFax7K1JJq4Dr/cBm5qMjq9wsSuc6xdYzRctDuTJg6xzsEd
lU8FIpnCMjjItnp5+FBh/5YsF0TpqZnUdabb3LMIUqt2GLCSp0/Xx+K5+/iqGeeO
hd5uiCrKwk3g5K3FsPAhydPngDloU5FQBskXbg4Pt3LvBQZ0ghimLdeXF+BSpWjQ
3dgP1G64lucKt7ifMLJF+xYdMWhg/cq+/kZMDJ3VeBhUwBElgO8g7sLNySDC2imp
ZmkNlELgZToG15qdWkp7MmFFF0NuIQ4ybSKuiJ5cVdaFK0ERuRe/Y+eKHCyQF2JQ
9YCE72dFW6mrbN543WWWsIYulaL1ZFJ8uUB0o4F+nTfJsWK5AgTnRvLkyBkDLUjW
TMR4rESX7+64s/gL+a5RyXJDX9w4ZfYT+mVe/yB9+ZsVwLimUHx891g6YHf5buXB
JFQNrW5fvvpmZX392JZTga3Y2OXXryMTLENiypFNnWJgsjJHsc77eM8zzqP7mGCt
v/qsVhyyjpjdzBSH/L1Qf/znbMyFyZdAi9RRXCMaZbBeVcLXmlpa2q4fuumneUyK
pG8ctXWuT44Yf0U+xORJxw/GOJ2YFFm0UGXjE3Ko9m4sfp3lQ26V8B1OHAP5R2in
nXWNYcAD/zVPH8cD/IrCEcB/xfNcPnMXv2C8dW2xvcVR26Je4IScfNJhuBo3bLG9
2w2g1Drt37oe0e2rR55LHtsf65jTr4sOEEh1WkZX53qQWC8q4gov5+5hr01FWDcv
C1ye8juTx16ARmS+6rBtPdpvS0ewztTXzt0TsdQoczNkZtt11bTAEwoY4Fi/DGbM
kz+mPTR9UkM6f75qS+nmQEpEk373feVZX5e/DnD8SrQSZPoLoPFXTfufO5ByJQWA
dnwLodWpjrzQcrIvVJRdPje4iM3ZveL9udXdAKd4neHJbE/ccN8t8RW6aFUAIzEG
RxjHAAE7zwDMJOkQ8JUtW3o29o05gCdL2WCMNHPfQzrkgWyQ+3wGNlIUq1GcaSmu
qSissN8Lndpoovn7x/T4SJlaQK6xFdAevFaNDegWx+W/fFlAsfj6k6bpjskq5Kiy
3nklExlGwEYSfG0qd0abVWx0cSydbZrDxxhJ/JVFj4tIN179hWI6kKGnP5BSs5oe
duSXzSXOdGCtwUmTejuGdyusQ5sYDb55lMKiAO+/nGTWtjoyzosBxgwWqttEF1x3
q8AM0EgOZNNbwaxn6JYHH6iozm5pZghiF6+k6tc2f/cGHaE4vlS4Tpu9vC1dSi7A
+yQBxqZhGZM2VW03llkZ/sj2TdOItEsJmAch+u9aG/YdVTtri+DETCBGR40XXNS2
52a3YxIhyJQfUQ4VSfVZP/+EM1ghRkU/EWqW5eGJwIKlW3OFZPkO8rAhk7kASpwL
bU557JxJY9ad8aaNCmw8oQDoXgHO47VzXaIYpk0jMyCOE/gEhB4zKqE5ipNqUKTL
FvJs3eg1XYhH7Vqj0a1zb8S0CW35TbOM6hEd9AvOw+oWPKNl2oooksdSIvJESRnl
jsqE7CwUBXw3iZJCObaKazbklI3X9+b1dWVLJaVf+2Z7aaJ5HFfwJHxRHeD0uMxF
sH+q2DMaEcPctj/GBJY4PIPTY1HVKjQO3w4GFBo1YRfUciEivr8cNTtY69I0CUNV
S0OC9ABjpF3tEK1AeGKFWt6/YaaCcRrLlunQ9hNrYjdKQkjGNfFBLCUb8r8uV099
06KjbLxL+2ac6s8nOecTg7WOOZUfQjGqe03fzORyNgwFn1ItMJiBsokWvJ5LR+0O
tsn9908clFCCg9RxUaUm2TZhHqQrwp81RqX7qpmSNOnEQyKT02OwMh05UTdfVF4w
pDErHIqd2mIp3eGjOCM9+asb8lgy0a7qyyODR4MbLY1m7q12qhErSjDqKwh2VokD
uiykpoQIaVIWtDyJCHjpQhNmCVWDOA2juKTTKiCIAJUrVz8iKZ03eyJ7V2ZJXfqx
dUsn6YGQH6eWH2zeBY4m1m3t0mb79LVsdtw5hfh6uyIo8nBCVGjOmZTNLx7X2x4Y
bqM24ex52+UsTalTEKx/haawtf63zuhbdwi/Y/pMIe3xqXUFBg9mvGfN9NVsse+h
Lrby8u5GNLGgcD6J/e1C0ExWafMimpYgnUnMjqBowS2hYt8JLSAt9CdH9R1XF2jB
1yG+I/CcwBtit1pyHo7531i4MDaMBNjhbY6JY6AN0nd/x/VTbafDfXqTpcHtjEzc
S6e2G0/cHCoWDVeb+rHmOo25tzuuNumLaC1VXADeYin9VLb2bS1l84yPe8Ve9kjy
cfhl8HZMjmFes3qnJcrswCQAWhl6DLZWwZImeFFM2b3kWAgTNVF84YHsiAkj2XhY
qgSvNP+rS84UYiRlZzz/X0vvCKN3ylGytQBSTBQuhhyvJYiUB/X226rH3fFPAqg6
ivAiLEiIGlrUIe7JFsQIcEOeV6khqcACYAYBX6PrRMAWDPf55fey6iTzzMHizLMV
NntT7DcLUWHAj9niltvs3FqcoNXJPZ9aAw4PEer4oNhFJQnWXpGyrDAj0DmsQsF2
DugZgmKRJXWizf++H9HG9NELAhrS1rTxIwY2crrk93reJ3OG3v8paOVBEof8eHkB
1EcG8wfL59nxCdEy44RHArVm/Y6b32OY/W8GTgeh+s2NFSfJ5O7kATNFW0kJ7EE8
Eo2k+F/5w88JCgWz/IQJHVv5PO8Xtq1ucnorGmCaGEqzFuYthIOUuOjVmIBOT3T2
nCpYoyVb5cw47/DbIichlIQoJZeCnEgLCl/LXDk63yO1ja0znTluRBUpdH3ILrKy
K4c/+eLfTe+/YgUvjj4amr22LaPZZs+ETgQGcHjLkVHk3fXQP4EPZtrndqVfB8nL
ALliU6QscLq90Q3uwkE+asgF2Nji0Gx8kJqDbaGXuIDmR+y6LnHq+6FUXmVg3l7P
c7G6o0Hx/U3GAxSBrvkbCFH06BM7Ih7d/RZsf9Azs6i/vgpCIZDqd/tVL1swkrqM
5pMP4CLhnQX4yq4byurEEBPIElBsGbKeLeOqTgyB9k5ue7mH+slOnDcbVvJYXelz
7fxqGyR8cvNMBD0p78/I3chd4Ddi6+SMistLXxgSHa38iGiPJhEaOBB3AwVlV+Or
WYJ0xegbQwLvMJiK6SJwVqJ87AcderL7NUkyUIquDXD8W+rX06ABVL3EJK+rmIRq
wv89UY3T/0Qzoz9ZfM4ZnwCIEFzC23YWIenOMUv+AkbjHdfz1keg7v4yhWYmw8s8
YYGQeTGz5WtRV0qyz/YTAyIQYtFvLjhjd25uX0yg/0n4w+RCqML2bXos+m8mXXW+
4h6jRQJu4GWlQdFBc+4WoEs15WojdsgcUXrxDR3UZou73C31QDYtBlfOmp6ooJKs
s4uSTPKdjP0uUdhRgFe1gZ/gFiaHT92ksvLYubh8C/CsIdd3VAu1B2wBz9yBPQTu
0TANnEZWMhtBnjdF6HUhtWnbmIy1FdYK7u7fR9WFLTV8RmHwduqWu5U8MlCbLkkT
U1ONuRP5X44y2acIyiBpJUunKkxXP7hU51e+CdgsFB+8rgVHJ81UAMp/awkr3mLA
wd493Di/dE8m/bRUlzEs1ljiUhz5Bdc32CESKGuzrF+ZFA165os4TAPuaSpiGZvG
t/0MpC9pOsWQfElUb9+TxCnBScYHe5zlrNpWnZFDlrchvxJAhHmnvWbS4cTtvJqG
MD6b7X66jNm/XPQ7J11PILApMrKWKlT9taey+xSfUrD+PsiT5j31JVdPZi+55r6N
+m/ffIFMyK1Cj1VBo/q6eey1TFzXj1rX7WzXa2HI3Pozztx2avT5qpWGqJnhv2Rf
rdfyeuhgy6lW1J66abb+7qMEgcuAbGoJqLnEnp/GRHv/gjtVzlJZkXy/CbjxClE4
3IYBLuu429DAc89fm+GBoeKEgpWRxLXwdzmxWODUdrT/COLVYHrqdhVFZqs+/kTG
GV/jhhuwImu+L4uBqiRQwEvmvrSxSxsDA0ntnSNIHlrkaNoUhk1om73uKohqW9IW
5N76XFTDa/Scf2A4A7hr/EN6oAbkK3/TXfj8298G60dM0io95qkuziBq3orra1XX
/mrKXcmi9IvhFPI9icHvPi+Pd1CR6fpN3D+GGxLGYzLrj2uN9oEwKTnB8IwajqXW
V5tyB3z6F+v0ulfWE9hXtabJKqilCuzNbP9+1Yg+dNqVc3PcdBKnf6fWzCewJTSm
b7DO4RmsBLH+BP23rYhF0Hzo/kSO7T5rQkYDczPeT3NwMT4noFGB4+tfls2xuHfi
Q0pVzKdNjApene9qKvWu9pGKM5m9meEHimCbehIyNei06QhZDK/3ZjXkNMLnGD0L
5fqZ6LdjDbMuzuvmQdf2f74YLZnvOy2N2lxgqzlWu6OqFIVCDyCMOZGQAttzs+aF
wBtaYBeeZmEOU9Wrt4E+qQwD47frG0ZX6kxQBT65/HsZER57wwTBBAhq0+JtDh3o
hX6GxJaDfxGksvfTb1GQXrolL9UFKC50nrHwJVauVCtxObRWdbQaZ886YKllwzrW
DfihRvoxREW43xyvpQBAwxtREghGpqWP5leGn6I7IGvUJ5rY3ghO6MxGVZpIMiuo
uwFThavhEpIPEIeUsjGVvIm5n7OQTh4T7Nkkeqc4iWIErbSKMviTiE6SVKhzaJfZ
348ekRlp1lU3cbnpcV3uBtViuZPMd36MyzrPEQOFYfgA0/cBjN6lR86PJeo4yih/
XKDuS9RdxMgFKWimgYlcORVmI6hRTYTjuV+L0N7ENvMw6xSK9tjGxiOzaSWjNCBz
Lh8Lt8wR9oVyuG/jHVifUhfXbFEy7lvZ2NXo7X2OBKrMrCZmvFbzDp51jXKVVNhR
1TWW+Evy/LYno5x+QONE4oL9CRdA5aPsrtk1byEY0gRCqKfcpjKqTDmRoJBgohyU
R+iLK1vOZyvoKD4aD38/bDyDAiDlqkmDbuTWDN2V1nmzCYOaYf6tcYJkUWHZp/3b
JE9RUCU4eh9bCQsEqPxFlGCNpWGm7oQFcz0sZTPCaa2mqoS4bMergb3HSNq71Dzi
+3pxBojN7xjLVwc14g9ISGzfyL9/g20MVMKfSxT0qIX+sDrDUy5fTDBMlYZeu8b0
WDsl5q040+r3/THkAaLGzqCc7uSKCbiFPtRzCn7D5jvghDTZ6eXyvzn7eZPgCR7D
5uoAfslQ4PCMzZp3WeMejIvAFTqOOrnHPO6g/6q0hVW0q6PsUaCn+qb/z6U8KTTX
I3jiX6qQVUbmAMEQJSOXan9df60LRQ9QvBHTJujONypbyRt7Z41n3qIKwGve1QYY
1UiaaIIj4bqa4rnXAWSr1bhpdzDE7UKjzbcIZOVpz5dP49ff9W5JtbKqbR6SlFPS
eDLQP7ETWAAh9P+TNfPQenSHWNugmGhIPxNORbzndp3Anvqv0nBIt1VZ8I/yTRi1
PMu8DVP9VC43YzbORl1BoJZ/33acleiLLutFLWbaYJGS0LtctVfFYt7fyI68IOc9
iqiQWdkHDRAO26XA07mrOobqc51OE4Ot+Y1IAiQRwpvvPSGSfSPPC5L/O7R9RWPP
0WhfD5lWwe1WSSH965V9UTEpuXE7j7NVEqzPsO5BvNPmf+JPSaK0fvsGQ7L2/goG
W+hJxDrAA3AK2h15RmRHRZah7tuww66ug8slPcuD5b1VYMtkZeSZO7+mThd7Ug02
UdB9QelUasZXWPcxR0DySzTHox9BAeCJFsgben7pHtu6w55zuIYWgXPZwyUhTdOV
F/G/xKz00xuhQ8/GH8vv3Gqb4kLxVVJub9XIszeBjvsQ/JL1XhrI+NiVAdxCKfVp
yOwmum0FdUKk99Q5g8phQecCFcfKZKKbdG4vRfouPuIrM++2+j+/pb4BaywjPLbi
sRIMX0AwPNkVd3OyeYF6PjLPzpzb3f3tnU3lITJ21/M4AUyBWKyliOEzU3ESvbfp
KnoQP90AFqLPNXMWUBAovMdAYZ0q5aDqwrh4DH/ha/CWjGNSwD+M4ipFFdYRXJE2
9CiAzFcIXl2/O3tv4JzM6uF976fhMFgJjxMB0ijJEOTIf5JFaVou2Ii0XfjdyE1x
KM1Xsk1JdX2STTN67CEccK73Ue6r9ff74ickKjMqyXB42julndDIyHAHhfaPWjAG
3cgnr6Wx/NSddN3b13C9gZzoRck79t7GZ2EcHEQQypwBnChQapGuFnZACxXltkiL
LBkfjbE1YAEOwwxypfoa+8MA5HCf2++FK/E3VIAPW6l+bmOUeIYOcpxHNMf3GMBB
xCy6dlIcb8w+ctj+DudCesfPU/ZBaMQYJaEp7kwFkKQ41jWtuagSFk8DRCCz+bPt
XSuYeNFqeunn3N2dNIxbqeu+G3bdV78k/l7YoGrpsZoYWlXEr6EwlGGSU5cG0uaC
BugN4kQF65JEWllWV2BWx8dkLJR7+V5TvTCbieNpdxYvsyhc0EBPgN/1y1VrII79
GzzBL1c/vFMCcMLrgnBSlZKyOj4T52ACAdGV8sRnYYxMw74H+8BLNwDzCj7Qp6KU
kdNkj6zvKjse0HyABQFRMizSTd1ulViv8BZMpjV/ey90yWxDZzX6t6DqF+LE59nX
pROXxtDBx9h+/rarUf8N4easUWdNHL3NH1vheO+HUrwEqwYf2S38nrrcczBCBKui
TBRvPcYk31AfpJrP4dTAG7qFl6N5LdpIkLnPw4+75VZxXyQzIc7h9Er+04fv2WhC
dfNmVhiMOYE4/WIPWp4C3ef0afZvhj7OoCNb4F+didMxQ07eyxDeGedzZmJZu2mX
X7Q5NGtaPmcccu6NYtdKoHO+2af4sAQGFRzHhWJ9doj8VrKhE5LotreBhcnvjx6v
blljgeAfPP0KZPsy57jSMoZbnV0L1Sv9poJBxdIW0VohWyjS86imdFM5J7CnpEg6
DEyt5LVBIvDAYeXADzjAU+wdfTcTB54lbCuvGUbMnV3jwLJLp8QE7DrpO5Yiz+9/
R3ukHyGPT58K47xO17YL5svBub38XOeWef7LY3ozOkU1IeBtw9wq1VJj9pNi7jk/
VTlsfzBYS1+bjmvvl9gHpCjokGQgfJMjKWvopAdVFNJ3kvIUEeirDe9Br+RHhSmV
ypAL2LOPM1ItswjZqj3Jimsv9+euVdAArUVGTYPZSaOLQFRQM4t2HXOpiuXFSrJ4
69FakrdQXhE3wNvPtETs+/B7rcTsU/64dCrB1jV+TaMEX2TZXt/MAp2/ZfcFoXTA
jKE39CcauA+UWR/EYiJto08tovHgOs1S6hK6wBeSkfXXZlfuInz93aecXNO/zcKr
81OkNXohzRox0MegdhrNDK3MANJWCmW2xkzUfNPiRTFYxvKIubRcUKEd52dZTAyU
jsZ/Ntffg7S41jdAO8VgbbKlxfkd5kuteS3peDPCneZHbcpzU+9kH5/KxMYRLt6C
D3WvWmIW6+tSwMcuA09fb9JMIpB+3K34e7+aCTOCt51/3puZkJxvixXAR54SRI+Z
ULvl7lSrSxeF+i1VjrBm+KvXuEFgT/mTdoaXc5a1MCPtaznqtPvkE6L9lUiIW7h7
J9kluOc9C+07nzmmqWmI/XSMnzR4vuPIoI691ssERpfsGSP0UfuFE/qXpLnCpeWL
k2Xypm0lL+QCwAvMBJXMzdChyLKRNZTmkgKlJT9xFdgIROWrM8fon38XR2DUZfiM
BA6LeXHAibAvGEX6H/jaZhQ5DfQPU8Los0kpzBNR1zQJT+mlkU5u3Db8toOxw0Bn
jqddkT/Lw32IAIGENQkqS+RMHoDmRgZyoJG+liDDOE9L6RT5tWCVbqoKXv5VWLlU
T+C+XIApZBpkcltWJml04R2e59VyNJhRx6d3xegrz81T9h0x6DxawvPT4nMIoQeb
d2Rubl4vcLL7uqFqeUbofkda+NonOwO0Ld68qhFZEBdYerAHy8dehBIzUe0uapId
hjrvFB9fLmVFLe0WqgPYMiVXC15gwSBjMRlFolNU2+nJTcAPClPPCwGR0FldeDs0
UhLrJEmzxBk/p8k3riHzfidSarePnl3SkhtWqq7HRnJiw0eurOR3WKmlDmJuMTxk
kJkYNpgZ82isF5whSUyu3BcWd+SccKJgJet1po8ZbOPhqMDESLnrvs62+fRUFINm
87D70hbMRiGGBJ00d9rvPE16ohkBuN7vPk2w0SAvLEnT+Wx9Y3YbcRzoiM+hJaTF
61tb7kX6GI12UljKdFXEABbxqzYNYmVE63bI3wRewKE4QsfzUsx59vlre9bmKX6y
SQbpH6s1b02pulyMfsKEfeIY3RFBT8Miekz/FH+krC3wq8jL/NeeCe2AV7Xw0zFQ
gZ/XnjiiLWJuKUiVambLMXAt9TVNWgPCNE0/SMlV4dH2gtU86VUbyt2m0YoDCSNc
PLTrh/8uEnPoCraNOWeesa16lTTYpc6F/qo04H+iaonqVxAo0A313nUCJj1UZ2k/
uAggk0fifI/HpiUDPAHU6kIT6GQ5UjwumQdhPIqCkb1l91spRe5AQMxfH7lpvKUT
riQpJtyIr8KxEbcdNLDyYVQeLY5meTn/8CrhrxjpbvuzTcgeYpy6nQQxnCK5haMR
0tEt80pfEdu6YQObAly8AwobkZ2hnIRGyZONMJe3TNfKWcxsEf0WyIBKaKFAB9uW
S4H4fI1aI8BC5zHwl+fvs9+RxZRdHuzz9DLT3c2JEfep1OpwdcQUmITDCliRrAva
BAvYxXqVE2vWpx7iq2B4I1r2c4nJHgYqvIDs/Ou9OXiugCsxxphzV5zAjVcFmUE7
H4GWcrcKTv6NsU5CBc9wZYVKSmxSautR9T3Ex9rG8IEAlX2KdBbqIMqaByZE4Jpz
7rUAwwTWVTyggXIqLQUsavutM9p1Uv2g7G46XjIQIPMh4Yo3HZonwHUrziti03G1
jjFwHNrV/YAgxfqrZT6QhR/zkBTFWDQqvAdpoh576zUXcZTKOEISycvj6KVLTR/K
45zJHe4lwf7iOP78lmnegALaEsoMgnwl6qaWIOc3efRwybzOn3OWtw+ShSj6bzbV
CLH+vwKHijKttKbXSOXkU98jyswKkZC9ZW0+rf61fDdCZR2gcP997Kk73USzye1L
T8+A1nvD3/t7Bot5k4SULRkVq+w2rCdIS6ooI5XCcKKsQzZ8WfIrK9hMXw7w+TkK
38L7bUmpQOUH1V1a+9LVOgOGJ36bW1AK4Qfk2WfmoGNoOw69MRNPXipzikn7L+Oz
RFHKQOhGuvJF82XAaaeq2ITf1e9iX47SGrlC1o3hJoYgydn21P6X29REDbvTUayn
y0ijynIAZytbfB+GfM5LZS5EBtAExbIR2clCXYVt6sQMvv9e4r1Xc33yYJF13tiY
9awqgDjRtvsfBC7Xnkffg8OQvT3OVdqXBQiDwC43nVQwJVPPvWNTnmAacKbuSXZF
jen2riSpjeTlou7T3TurYGor7goC8AwVSEyj7jNCNIJp56MxnUm/QDFr3s/65FwD
O/2XfXi1gZblnVrn+IGuZ9OuD2AjL/vtzxfDoKKkkv0CLVsdA/6iSpC3+DYl/mlS
WHEn5UHp4jbVslNfJjNFvPwSqPXRAy7fx5qBH87dt2A/TSIiZT8/n0DOiJFr15y3
++l28tD0PFPQOeEWNvi9cs4HXtsRDQ0DeLo2Hjz/CoKnUvNSV7/QBDR3L7lDYgXb
Mmuf+dsRJsf9DK84umPNJuYtPYJypocHW3HgZX8nwGKZoc6hNXAKdRUJUrjma1vv
sbIwu18WOZYf3vMZ0hrK8JJzazR4hlNgfmSJnrdFcNt0l5RTEEi+5TeZZOYmXoSq
as1IaGuSaNaWu3GO3pVrTKQzlnXsoRIhifxM3FoTxeUn4pMuBMjLqSS/k+fJzM5F
PybTxoVNv8KpbbG3CHllKb3w6UozqDl/6z/5JXRc1ZswL2MED/LNZRJ2H+WtJSHe
dfHYEDh7dtXFcLy+sHIjRt7ZXvtCMTpiFOg5Oi90MamfAeCHrh9B1m4WFDEm7kyl
P/wpFM8V+Si+aKOU9uoanpcRR4lNxL5hjJxNr2RGt5t2iPN5WYYpzrrD8R0Cishd
H313AJSeSxsA+kUgWbsEU/5VkgImZ13mf9YS+/Yx+k0aLybymGxctyQo6qAWyPW8
mqrFL/r7Iq07NGkDuDER3cY8kgok4VXVjRfs9CSx45SV80i744NvV9RlB1VMhFas
HWqtnHMs+WNDURmbHmO3/Tf31/FzOxt2jfrR65WHiCTMxoCp/MCbBFqAxVq0d6bM
qC2nBUzNP/Fi25np95crFzV/DB6ztpFEZRhaVcGeC32fn21WDffFolzRetzKSh2F
GvNk9amJjY91LuclMOEyqLA7jfPZ1SO0pMnM3/Y9623RmZQBpBlyzmNdQbma8msU
TUEsuUA9JkUD86Lm+NlljmrI2xP1qQWwnL7d4SMK2z8HA9xZPsflZ8/gJcR4trFE
cG3CN/BcnlMLNbLL+VqkpFeir/I/3gncAQ0noKEhxNNwI3HWMAwJbmu9AzclEIM+
wsy08SnhY8sS/nyH5aWQ7ttWkuiNYXyfOqVMRTeAQnS2tkHH1fzQC4iKzfMGgyrD
DYlCZK6Sjmt4B6+Fy4A79eJr20s47K6um9RM+OV6krgFe5cvvBC+FwWNnet8lffV
SkSGz5kufzeA0IbCne7l1eRj5EbKcwzKqoSd/eGCpiPC0Cck8Vgj7UVFbEZpHa14
leW2xpLGkmTkC5eRNzd2uRrxHPJfCVb+K3p3jewb8w34u6iSq4+iGwubfQRYD8st
OuouH8AVwrQE1FrN2ghy9Nb+HSkqPLZmZAPFuz7dDJnTRJm1VosHkK8++7X3Mgv/
cuJJ+c+OrpE/xiAqzfY2ze2i/azHTgBXPTsNBLb4GtRAIZ6JLwJi3j9qIFLX9HkU
tTeDylS/EdsFIugJqd4KY76inbpBEtLj2DzLvQ6FOrggn843xednJWBOdry1aalC
bo4Z5d1PNzLOcxau3ULj5mnedkcLF853gVFtAml7EyaN9XsFSpO59T4SpoZkr5RW
tr2OXqbkCoXL6qZxhadIgCxViU7biKFXKx65XxZAxvxrOjSLbuUSAL/Y9h+TshFp
SiCdaj95AYQZBP8JL8z6qGHgvm5/8CdHQUolgVEPTD1yPgjYsYfwlDFwa8OjCv2a
uv1kx242PghRJeRvqvQuXX6f7e0/uuhL75b6yLOyjJF4aZf/lASHf6Ueh93Rs2+I
wYvRXznnDnL/AKw6L43B1mHF2w+ndjtmfaQ0ZVtk+uBg0AhfF0YsYWjE0c5XNpT5
wrSG65h7L1z0K1d23X2VGkpC4CgWKUCWhA/3iNd8E9ZtbF+vwwi8DwrEBTWXRXDo
f9Pxdc/hlyBjDmHy5WeL4JSgyYTJbV93Zs5+zC7qCetPKDdntVsDaL+oE/7+toVb
B/XJSR0ztahZhr7Pc1ksh73VhBi3jGPMtVUl3EsoEzwupMwts/ZtO+XQ/neGUUNY
T54eu94TPJGC2e2AiSuWGDED02XLb58hRxXuBK5S/GBVrFy8ryPCmOvhqPyMwVIZ
OJj9iBOfGgkwDld01KoNpoBfdIO0m3qWQg1/PPwrlYa2URwZ82uubH0spHeOZwC9
h6RL7Uk+Gz+eanIWEuXHrxoLepfljctwDV1MUvRJIpIiaqWd33Sh+Tgr1qDa7SZT
nnaspzq7oxUIF9tKyrs7YTgEnNp+waF5GKUJD/tdD6oOLXE38GVMGV3R3jSyg+JU
aTGr685edNmqrmj2pQOVZhVprZsfaMRTkSxUoG/MFNVF0YSn5qTK51a3XHAV5uxk
qzrZ8/9u2O9UwB9YjHLpkFNq5xiStzGnXBCG78yUSq8qtwIaCE4nm3JeXUEg5dnX
2kBL8ol2szAXWy0G9NSvt6m1qW53qfwE1PDVuJtJHOkjY7hqIfwGCqMsneQJWeeB
D3T+XTBnrF2ek/OErreqlLpXiA8dYzUNK4x80L8M/ayoEZYsvvm9Y8nHdMNQhfyn
MLOL8L3+rr6PBowzJlQc22eOtzgpuE8Rr7DpzoHnrgcIa6bSFBE5g0+IZiEpD5KI
4VMqZ9jRmLXB+q1xvc9mYl60Z9QHXJ4wRMiOc/wngTMqj+sWfRgmIBuRsjDVTTjK
nJsEJ1+1tgmZs3itpzjOqSDrUHV5muYYhZMNfmxVazb+yc5gSqvj1841ls8Avsyv
2RaZHXFet3nag17brrPsn5dvUko0xEvUziEpM1F6O/6CNmr9oq3iWPIcHs7bhuC/
bsiNKlPgvbbR9e+n/aXQHtX3IkaEjgUGOAd0rEy4CynGVVL6p50Q7M6Q/7cnAXN3
PCWztcH+9+Fd8SHAInhNYri1RpAuG3IihUrKWovlicm1bBxTlCsku+GminfqKC0B
h5qnJ+YFoCV/fve4CzaxKfS3jy2lIq2EiZmvk5zScKgwsfTbgBckeNSD0Cw799Wm
avaRbaYkJekvAfA+REsqLgOHNUi7aAK/1RYM/ViDT1AOAaSdI8zbxi7Rpi0BWNUM
nrkDCVy8TGq6m0B2Q0b0lC/0uzzf5i+dZAxaoLQveIyOW66gXQtc9QAXsCeKjA2G
cX2rFH9JFUzXXkutMNkuxhH32Avc6YY+I8hNPKc9NgS39+ltS0jzmsAB/wQ7KURu
we001z3k+hejf5iS2hHykXo6Vg1qSYNt4+sCy0xNxdN8PqejGUuk/d8T1NsOaeXR
cmOnL6KKnOQQ5OoqHhPGHyrmceeEIJtk5rgpcZRuWgnmaWtZG2R+VDKee0Uphsqu
JZJ0HXfo2x0P9T6X9hK2NTx7aFUY2VLijXX/oxhI726Iz+yBnOosWDDhShS6/w87
ABizr+Nd/Rhtkv2gWPeMgBetkPO6U6V8gIU41g+EfY8WLnzKVVU/zI8LtZ9zXS87
+4560coumkgPUFFyug5tLG7x7ZeMjL9Btc5dCUqVOfUT8TjCZefVs6zjrW93WcDY
aj6QsLFLCrEiHr+CItoyYuTf8nonnJjkIl6dKWEdXUQtVKpUsZLYXjAwF7mQU3JA
FgeBIxt6BVJJXbwmUbdoUBZcSSkkuBVI82wcxMPeKTcDMZt3Zq9myD3rlP7BvAby
TGUQBPXwaGG4t18Azmu+GAexdtJ0rP7S5ykEYS9v+szaFyW88dub00ilV0zoGMPx
xKgLMs2h6U7pAJBiw8HuuiBDmeIkbB/WpG0QCcB1zAVdp7iMHW1vVfmsVR6Hzqfb
p28dCHQMwvENombNZ8Eb/a2p5dol4DnVLD8fC04DZAtUCLPLK0FB0jSn8Z7CTNLa
uDOQZML3eZmTyap8oCzThCTIlPMu5uVQ0V7GbDLQzq/XJtELPYcly7AjIywxd6MI
I6Sklf/tMlm39ZqspEPXFVb9AXOkrLXZTGK8YOE2yu5k7ha1Tols00YITwWgrEPs
ZACfQgog7hbLfM2ZS244vxV8IN/q3lXMSvXJACEAkQYc7Q/6+Nd4bvrjNv8nXAqN
qoRcZ8DfjBlnRIXkgmzGnE6Loaw6F3cM/r9XteuJRJcQ0WOmP0If4UZCwHC4GEYp
92TwdTcWZTY63PXM+hT7pdAw1eXnv28Ld4NHLZ3ZAc/dafgbl7ciE+E5quXbZ/N2
Rve0Q6bHl+mbkzOhd7YdM5dqzbbm+7V+ERqUzVfkxGhhQ5XWl4UBTHuChBaxmi/O
t/XTN6AKfH+NhxxC2Zs9qJiVH8Q29N5hfC53+p4KFkqvpIcn8CLSHdISDRgFNQXo
AGmp49Tc9gO9bqUE2ztZAOkxTEPzPY0RizaZ4ZuUZU8n1mBTYC7WbkgND1QYNJFx
iv2RmsD/lyYkPzrDixfiG591crMCRnpyfRLbBxLFc0XJWVl9L06EpaGn13vDPnE6
sfatWrIz1G3fd6N7fP6sPxVxiSuub2XbkLYJM3pCzTrFvxSgOW9Z/KFumsK5KxS9
IpJ6na0SdMh3jPKhRX1hxDWc2Cq56Fmj1icM5kuFUZUyW4tzi6KbxABxVMVnsanR
cIl4UExJj7Q+C6T8CbCoEkMeMXKfaCUE/q5O3bcaZuIJ02eQKO5dy4O68nDkOQ2m
QtZxnlXraL9kX4sz5EJXk60XlJeWRWwGLSRZq7KrTXnBkV6N6ZwuOf93xYPZVu0B
Oez0OgAADFCDZIZCCU3GvrM+lPPs7a2/SpqS81H3oMi8YrzZ1xLpZcdt0nULpaNv
Jg8yQ/zkRcRMWzxNNpDIc0Fw1PO5EbvdQZUyMjMM0awi0Yw7on0IjO/2nItjLeM6
3e73nS3Vg+K6SK1v9e+uzUKfJ1MkgTOqtcbW989J7juu0JuoJQsbd3u33bxYtdve
ZsoQFl8oUJjKjFXSWiaFqtfMPhJlS2fpj67K5pSr0h+f/b+1mEYeCwFhcP62afkS
Qbh+YzBz3oiaQjFjB6uNmETHn9FTUKoh78TTeXavdAsUIiXwt8hbqyY8lWuiwSuh
rkntA/OpEaueRTBv0DmEUKqQiOpu68mS/SBlds3kpG+M0JkDGgqpnVMILuri5Bk+
GLU4T6OpAUj2wM+yFFhIA1wvxL5VCkox8CvQTTo7W26osslJR3/hUFQEx4dcgP7d
qWjrQ33lsupBxGFWxiNPDPVYY2/MAy9qJ4ty3KBMDOZ1kDkbZCFmPH2R7DucvD1w
DpwHuMD9QqFyszAjORfo0R9+DYWNnSCTO7vMK7KSojX9xkOkBJHO/nzcnxst5cLs
ZxyRmo6hVfAbdMT68hjlriLsNKPHQ4hACoVauRWlUikkFvUaSxWLBDB/7cJaXdP0
97nemSxdObt65syaiGXN1TXhfPhwDiT0TDp+5Szvai/gIye95zzC+r9rWOm9646J
GNPTVsZsVoR77qoi0Ecr/DcqwGCxs4IEDinpxmdxUwFNJExkzcSZgA2p0R2YwwYj
4TTxHan8OkrBSWpP04WzX2Sumf5CK637pXA6A6tMHAH3+IaEURE5WTD0q9XlYgYA
dIA3Um1CeTEqiWHw5n8mxvbNFv1bf0PweyXGKLt8byLDEfUapmvr2zwUOca1DxxO
8gJETX14j7PJbjDU3jd4mGCUY0L0tjSnHjqH/Btq97CCo+I0mUeNLEDNf3/OZMFM
DqrHejQWWUlVN3/Ly9YDQtNkr6vjjZ86vcL9V2hjjYf+9/RaeRmaKFlqHpMaNIDQ
xp5FwOgyCq8VjN3RadoK3r2Z8VceUhDbJAKJ/iN4nox/iBQZ3LxyBd2mRIN0mi4h
y8d/sE4sIlmNhsspWu1NTINyDCPM75bxZXbZ+LfL/IBWFXXgi3wTh36+lIVcyQml
szUDEzJnE7ncUqTrIwZ+yBJfs8TrIvfdwoDYvQ6nu7nmHyczSpCwqBzoKhdeBQBc
23M8rXw+1GVPVOzKaXg4UYpHOkoOXeuCxYLgOVUk2sGU4nvJCjkebPMEGcpT/jmq
+mARvYkw7pjo52ABlsxlaO4PJRCTFPpvo3qgufdg7peAu0+oyXD8UDlMRc0T0KmT
8ZYvW7TnqgjtIV4Sss1OJ1ht0ac0F1fPnGMqLG25zIlRMTTJLroDFouw7EMSeFFQ
Q+qUALCxaMvuWFberfkxsy4ElW6weAYBgFHggXqXCWJ7MSzsjfIz18gVoUO0bfqF
8TPyX1ChMwJC4mW/iFxURfFmboNS7qFF2KHALZ0GN1Du7BXYgYaHQ5/IOL7uz85Y
sHmeuTrl+tE9yW8kGaPEhlRjHnVR9MKr3+Afug9aVray3PxC0C449CTGmrUZF7lL
/wgYMUVCrFubva1m6K1tungsauuj0jWMMc4ErKzE06zNbtMWi7+siEzuamOuT35F
Y79xxP6dNjxla6np+erymMAZInanAaAK1OzIyHxGTTFZDaS8jR8tbsnU4rjrQKQM
YCa3geHhYtRY7i3GtJI1rFe7OXUUlPFMxb4NOsr07Ar4116xLtTYpoYocfjkO3bf
HLgJI8pXNipYgOg+g3dZ4F9Xus6XB//i3cjQpKEVUr3FIDQ/mTz/sdWEQJuV4kdP
CUVDQuGFr120yF5YqIPXw91uMpxGUzs7q3zLKZxclIyZmC/gHElwd7O7NVbYdDRU
I/8g7j4dVhikTe5O2r+ySG4KnQ27Kw/N0j/CxjAaf/3Lbx/Sm8LQfoaeg04TJqnp
o3hv676CSW6t5asQIByqBaX0QiFJ36CLV2nQnG1Gok45te0mumMrIeFy12lDCLyk
GyXIlGEdYgwH5xyuHQTC4QR0jzx7wkPYSAAOi5qHVhNQZcRuREmXeHSGxw05WHl9
Eg48ZUcS3F6eZI+1AW+lAyfO6vnA5pg0NnpT3E1xE2hXZKRg+OHDJhJuwclg+KC2
47ouvcP73V6o6kSOAWudroF6y3zLFR+QvcOx5wnnYrMzCCLGhBxECj1qPnlBQk8b
P6zud1wBQFLx9g35p3cNhrXklPGA1a5F8U6b8pb2YZl5R1s8Fd80fOF0vsFW2fQH
3PM927j+RCpiGNj5d4YrEmJVqcRUD5nPWHvhvav41BaJRWUUPVf+VT44LVk1rNi0
IgvRx+VVA1tH/pZERSl2gSj3XAawMTlCdxfzA59MElboSS2AmHDmOyxumvO0FG/M
26GWwWBa0nZ7c5KgVsY94K4bLeaoTMb/QLIFlpjrhas6Jr1VuKFFe/QQgN9mtANJ
dTVnzG7hdoLkvX1bwJyrRCKEHQwi5gLb0ow6ZkwU/hKKf6izGsPcalTWBIKnPneC
zgWyCKN9ZkTbUMpNUxpfY4OIPn7jniDAWU+bJS828VzUs3Vm5AAj9CrQs9/n48xC
DKyFf9SLyjBwy/DS/ZEVOP+5pkMMnB3m8EZShGerEmr+MqYEXmY+zrtMDXL6D9Bj
zPBnJ+ImgE3sCvhbxCN+CVph+Dg1cpo+zCnVRFtlOCGDdC16dJ/nLVjTM1G1CWmC
yqEdiVelvERXvig1p+OSTt8wIkRF0mWRyfPSUrrLLjBIXGo/Md1E8AHrtyMDSInv
TQKmCH8hE/Q4m34XfPam9KHRIx+7HmyUn2Ur4KAHkZdFP6U/3GqT3s1Z74JhcWGr
t2skURTl8mAGR1WQn7FotXIH/Ow2eHmqnvEHmnYR80m0xEzU3ZJk4sJhX3xfrQJr
hwBuYUvzdd0/Xa08ZkoRtvd1yeOyG8Faz+0uWW7o/uWn+RR1/ev5cS5cstRg+bM1
qdyhcWWyjNBuY13PT5PzXJoN1j7QPCh12wC4LdcsEnf5Z4tJ77VfwDCxJXWOtBIX
AbtmKmCauUM8LLYECfr5S1Qe5SP2DBfnR62y40tz5NdsrXjAzWg5NDu4lFUF4nAi
fBTLB6V5fjWqNUgeVWx2/vojh1oslC5qNUAnwMCPtccTLzXUpYe9AE7ml8mUsP9g
o1lYFn4wWF4VVa1Q4VMLk2tcAAuLmdzGjmN1T8aYEvixNSr257P8P3yzrEZFJ86P
hJtd+qItk30h2/MafnC+GHLYxWTgO+hrWUS7MfaGzkXmDr1LmcX09d7XAt8fGu/B
6SCU1HWiUpJ8Iyd4FXyZ5eqdahfq8F7u0f9sEmfO4SdVOZ70wJ402uZVadRMg6YV
upkROFzCINA9pxnisPD/LeIHvKtJUo6ZQM/aYNmTXdn2T+PQXo5UsHufPCt3wuPM
voObruYTgOtOUBEDi0QD2tvgErcu97Fb4F3kSmKPIPFIQceDV1O1qKKZ+DdAk+xb
xhcXu/IwE6fjetPXb+Qj0JXPx2oa5wbYBXeoShPgv5Tmeg4d4l2RQ9X1EITDdU4m
rKu6Q57UxTsidFTXUOd4tXkyromzOPAg3cfB9vTcMlnHmLvOw49Vg1g/nxbcsyyp
w3Hn61l3JM45bbWKTvCux6ZIBS4qjCV52INPZqxp0963EqUFaJWBVrEQsvLFsCSz
AFGVq72MJ2fZae/jdB/4lf3a7tJTRj71w+iNSYm8G3AbpftLJPPIGEk1vslUy+wy
qy94Nh0xnkv/w1ONcm0q6WjBY3C/BT9Bhj4owPPndp1IvwCrFZX9FIByBUKEeTe4
BA7PzX/AdiyZQYb6JrRYEf70Yr9fmfgWDxaBMknPAu3wv0osKWI7iWNQ0+JviRZZ
qGV6lsxd6JCQf3+OhIyQMrevShGnKnTG1SUHewS5+CIdNXvcHHLk7xpq3oX4aTO7
u7Ws3O6pQBDIrYQfz7sY31Qpdk8I1jVQWWz8w0fyn2g64zQFwIJ3dvVvhAL38SRX
DT93ZuJjShZWVT73UfbJqZMivMJK32pszEzVsEGYqpVlOv5vvgqb2SlXWP+sLlPV
rUgeWPR0my6BlXC15rQuXeU1EbSqlp6KXvJfucUU8DMFjZpQnIWPC78/tVxOhrQz
j4n4oxmeZfDna5fLCLdz7vxYhpiPmBGv5ftd6+yKNONOfglXPsdD7Vz3PgR2hxA0
qsGbtSUTGEWP7voI//yswcD4ttZ1gJvUt6uJNFx5i83F0pUnRjNbaTvSR/sbaBSS
DF2QI8s5JNXh3CznycPC4lcWVPOedJNJorSNmZsRrPbWm2If1arm/OrtEMx+DE7T
wGRijiCeJtUGOcz3BGy+zLWzUbIG4q0RT/ceTqL4yZMG00/+89TrPpFtV+BJ2aKO
plcmOSQvri2DDpOOqVNaHCFhUXaDgfEYQ2XOr7z06I2Ulhi6JquaXHDgy0Kuz/CA
c8LdTAWKQOpy/8r5RGJdIhDyZY3Urct2aI3CpBn8ognaupgGxwKvFCRkPdQc+5Rj
13JMx7eUS1cbNoTsM2kRxMcuydYXJWSBf10519q/jN4IVDnODLqzKs7oZRmSNhU1
f4wx8JkH8AVlMxmXW6zmMAIeQf/cgD7xtTY/bj4qkLtiF33Afq9Z3giUF3Nuc0df
LdWqxq+iCWiDjEUn0B0kAm9PCEeo/VTaygNLLaL7OxIO11DiLa/BzsdErbHpDjQ1
aBlDCehrFj/8152apk4UEVdnF0fZmsCABCBsaUK5DEDukYeRzQCLepBQnqcuMbRT
SeTzAA2xZxO3S/v2FWfIygsAEprrBFVP1Y3YYLxpUyuekJaIEKH3fBW69ql8fk1i
JeOhzoj7D/Q0LNMS8JJWLz9iVm6i2Qjp6lmAZzwUtayb17w9tAg0knza+nPOkzcN
Z9XGSHHpriy7NAviPcdoivIah8SPEKl1pb9n80AyBmtdTDXEchv5rJrjx2moJzQG
2+rzo2McUh17PYnNhbrxpuiVKBI8C87DApr7aoRIECpZOBROdrXtsrgD0ODbT9yr
xZocFWH3i5A538mMx5o/AX2dBav31gFi3fAZP9z0dA8ghGfcWHAIBbJA4mLeLm4Y
wjmiHIhsUwuYbDjDjFGYZJxlG24y2lLNC9mlmKwKcO8oYTzWrA3ZEUTy4fZp7Z2q
NCh56u3Zmchw1BuH/xZ25zV061SEx8Byi5X9qtLVJwa8A2jkfaxDrzjGCPe3dN1f
OdeMTtp126mIq8QTZ0rYTvzn05U7y9/cOgGN9J/4u4cGxqFPkUDMG1mlV5H97rG0
w30QuT/IiSeVgdfTx69yLJq/HbF4yYN1jX8YVw/zKu6j5l4dJgmSg/8NnUQhf4Wl
Bwd8wNFvurPlCHlxdyF254692rdIiz83PsHdw51itxVJv0YXtBga0nKyhMSpEdg4
mDDuNTVnu8m77QCxTNrkdT1jXovlTUqTHOKXszI4q7Vb6TL6Gom7upuo9uTlg6MK
7U5mgcNjEdwmlE4BGFf2z4Pc1n29B1Ravd5XhD915QkIaUCEXbr3HCMi82BpGIBX
5WT5BywkUBaKoHdfClXN6Arye8or6i/e/ZlMpTttL/fF71xA+EJs8jt90GISQLsd
Btoi6pCemwb6DgNQwbH0Otc/l4GcUCgjdlmbwbnAlgt7TEk6uXsQq8wqCfT1b/rp
YzmScl4cZN/Yx86P1osqCDk4ou/zgqJI/IY8H8OyH7rCMXES8m0cj0yTR2aFI+23
CeTGM+0FAkYdMToRoCw36PHREjaSydJGYzB8hZNVo1cWB5wEOzcdApNHi6ke/UFn
1eg+XbtKgUmQQV+Yza/1gtZor8bziadDnKnW0NBAzVyGzLRVGQgqUDq6jG+GaAmP
Uu3j5v4uNLG/AhXVKpUi9aZCw+34ZygU9Cz88sCy4c3246ko1PR9wr3v1Hs7w4yR
zfBLBLtIbErc6mC2wrtJTMDGYX56ckDr3OdQUn8Yu03K/VQfJ3jH8H3jg/Y5uQcH
bQ3cGJYFNbDeoeK7sQ1HcSt5YVkrW+usHM6RDfHF8LNjYcBZQYjZZdgZcbmusOkp
aD9/MKFVDI5MT/DJtOlgargRCHk9pVvSe5XHWKcYKenkn6mvTT5v3LpzuH/st/RW
ASvffaKr+87vGTBh333P7f/CzxPqI97wCuC07kkDGk42Pq59FkdORzao1NxuInp2
vwr267PvXNkqssTlNYKGVIXIKBDRrq4JeL3Um9m8X6GPgOSsb4Qm4wk43Jf8zEhf
SKmIYAOTwrgKtPfot0XSUpMXWwwCmPjXWawO4/V91hBbbZjwSJbimxWnOiEPZr1V
g++X2LrjW0ogfEKj8wiXLwoi3S9jFPKUtdVbv6EomV+5M6mHkW6sUgvnprGR8Qim
v/1N2Lx17NZvzX0sDLMTsptglw24nSMMXmAW89y04wSZVlIH28ZHvWUmEqK7yFO3
M+JjxdH0TuAogR+Omp1Xfi8pkBuuDJ27s+6dLSpby9zhwbAzAurIKSxYad2qcW++
6JdaLGjeon0pYsaNPn7TOskgh9Rd8JqwEkFtrsPaaql9cQsthxrgC9ROASH2jRTB
hTG/uacicqwQANWpsIsXQEr71yT9EdB4xWcNeEj/cHitxIru+1323n+NwUDFsrOO
sYpUgjRyJEJwtryRqARsNoi/GRSE8WrN0rlJgHFWrHYFQreyWjAXC5ltDPuSideq
u1ooB7ef+YTffi7OeHEKga75eBfydU+6s5Uda+Oly2ZXr6UyVdL+VmH8suKeTSeF
VUWHE0MvKSraQk5lGRPIjXmTeRafLSg3BCV1UQlhPLcW5SGkg1d/Fs/b6IsxAFMu
vUnZddLCTxla/y+MvqcMpjL52pkElt+wiO42rnaas022Lq3J+FMsXBQfCOhxmuOJ
dOl5531gYhARumNyJT84yIKJYUoELWZJIgYyES5dTon9z9owG5TdSIsh9IzxpoTw
pCi9E/ikxrbTGy02RlGd2M4ED0Qb9m686MyQ7m/ijhEEKgPylsSX9hEuqKh7jX+j
oAolIIW+7EA/XKQ5j58jiYHFUBG4QZFTrwYvBY0aNaP8yB5Z0p29bD8wG2MxEin0
JyE1geDJ2D4NNsjt4ovMuVdDMCrXKJoE/TLtc4NTzAF4cHMx9LRZ3IOlfqErASUH
JcQ2m9OXXHSOumTgy+nYYdhVmAd7XK1riHglPWB+C+gIAIoevYc8JXrBUQxZwNa1
Nkj78Y9Fx6NcDOyyOpY4oRduKyFCrrMZr1JtEQKZsA7d13aY8+w2DupdAHvG27WS
uMAC05WsyHwnMQXne7nd/kt1aorZ1CAIrni/Unf2Ivy4ZHpeMUODztxBgdEkhfHr
uyntTwUe3uEOOWv1xhD9Vi8EDuTlfOST60KsZ8FdHzZmqTRvXrAgYZks8WwG79S4
kyqlfa1ko9xzl+RjCn/ceC9CbtXhOkRuhweFG8QN1AOXN2A4Exe+9qJ9HGhK/kAn
Ei0nQmcgg3m5m9nSmd5XwqX9c2M4m8K38HUaxTtHzbtty4dmosim55Lg1kKn9mnu
JZT7W4g8s8iW4Y6rcwzJpg1Z3YwR2n1Oae0HEleQ5Hw0ZRlLRN9yuwowQOBH/kos
ST7Aa16bxBVEvc0UjgctNoC2uZ2H3M9qLHjK0IueeQy1l1jG1js/Eudyu53UI/Zb
6Ebfw1o+VXG+0DRg+iVmMG5VcLxC9VkznPX6wUPEVhAUstJh6UzekETO7auiropU
pJkFbTxQ3fItn29PXNSTWAuPYMysoyxClRuplYtpJI9LxnrVDXUOtnnIUkCaIToV
M5ZFPJQw3Fk7xHJKo9l3/OiW9zoDsArPQGhaqWQ0d1Q/vwYo45nr2PfxyMIbyfKl
bdACgYNyoM70LGaF+pWyHkDLMxTeP5Og+0EnIpwG92ZzHYfSwARZIeJPkE5CpYZ7
0ZUZc3OPQq3uOcnpP0M89ZX0MhoyMgaknE8wwiot17ne4j2CHxO2/ECcJaq6KUgN
aytYZIB5d/JuabvPPhEvi9J6fKuG80p5LgyNSgKaBIWI3+huB7nr9x3pNgSyYXla
61bd4mFBxnXlrblPV/mASSeoyFlf1SSqPotmlmNAPCtrShT33zS/bh2VFX/8IXGk
zU/j2w6FoZxsGW6QYbs4lDDv17aUn1F7fXYuN2w4F1/vTaSUvMDxIaF0T7p3NVeU
sRDGBBlFjqxKox+PCaCgfeglwluQ87yDYEmvnYrWT25bwdn7wnkGs3T+6CDqGdmZ
qKIDs2QlwzDK4gc7k2UiL5q8exiE3Pa2pAOTQMSgyPs4HfpmxepoiNUnXPzNh8Rc
EtdkOINNYllZgL+E52ByGmPKfkUv4kEuq5U2XW3ISTcbiVh9dbXfczQDiVRvrlsp
uVcsmR9mHFGJmx7d16yCDCfHSBlB/9lLPT01NQR2GlQEr0TLd/m5UrmuuRgspT75
307vqqZZcd3ylQaYqcWpB6UezPZ2UjNDp+nX4MY3NwDeO3/bKFnOJ6EV4z2Ifyo/
ZKnVfWSoFm7c6cQVHql9H43BpmPhQrReIwKf/MuiogjdaMl9WkyA2ZSJ+etH0Kuq
SGy17nrzCN0ovQFmaePlrqaD3/671Eq8PYYq1vnTu5t4MMqTTcBZ3Dke0oGSXEg3
CUCSHP+sj3Fo1058K1NTIkzD19V0dy20zhxTqOKObr1vNSeDLapWFURWshVJTXRt
9AC7TLLWVqm4RehV48uZhvUPbqqvhp2wSD1sLk2Fj6U55UCIrqfu35rQNp0YDAB5
XmMk/Q09DAUqq8JqqUyMplEyjPtCsR72+UdxAdb5t7kTj3YIV2RxraALula9dsUW
w1RBvsxRat2y8HUj2FvhyDScx8+4Bw/x+6q1M7IJq7/Cz2ovZLQR1nqZpPX/5PS8
3zl5rItofDWbEneVbGPRnkaJ24NmGctWsDmFc84TDJ74FeT7An61TQLSfL5VlmRp
SSaI3LFjKKG9oUfpGBlvcAY9zIyDqNt8xVNJt1DP1yNO3LtC7LNKTT/h3q0+exiT
1iumlEG2GTBj70EWAhGTCPdoLGQ/exlXegM1l0QAiNaC1LSP3M0E32gCJq+qKD4E
I+vQir6r4TUKE1a6bpTm3UzBPe73HZZyS/ExLv32biqzpAkTn8zJoKbt57luOBkJ
kqdZMXtdYqTiyphealwTfjOkPdyRm7E6cKk9poqa8Vf1Wgk+NGi5YTCEUZe9iKlf
3DTGDsAQjJ24E++0jKU1GVqnJAZHXo1j1xtTlr/cUmqyTBOEmoM9DnhP23v8+7ew
hH/NCgGuUFy4oHM8TluuZpc8uxLi4lEtl6LDuPQrZHfCthuPQeBFTme+mbgA50KB
aX43lILDRMBQhNBRqXA82IC7NyZrIFopGvwjdWMTBOQvTMNIsSif85MNvA/hgxds
Nm4qDxjLjlMQafdU63E3KWJRdSZylJRlCCkS9dEj/g4HE9TU0tB/dM5Z+Bdq3EBT
Alew/2RmMfTJd2Y5Kp4djqmjQNnYnREBN/JXJAKmZWSOYSEKX1tEk2wpUSUrNrMM
FiJIFO2ZZd4ng6oGhEZtWzKwMb6lDDlg6sglBhpeDYma57CVFAvYB/2V9hjba3AH
gJpVVU8pGkVHMRcwA404LekRyyjlQpUD2gP6t6GeZeEZySVVdGRAR+Lk4wP2iEeI
YYw8BL4kRJ+Od5azYV+ex3wqNohnDiLrdKnv5kEG/T/8z5eguCK1xaT9xASdYW3p
1paJiIAifypWS4pyHCXIuzxP14kkBNKmo9k4oRJyC5K4uklxPHZUlZwQQqifxYiJ
4Rkf52BPN98JdKKbgoBagWZnY3jIb1BbkzdFz/rKZZg3Yv5Zzxuo2ZauhBcjgafY
kE9dxZS3IvPBjqO5NF1pPo/MYtgx63cPiw6ShQhDZaFzkoO1xlKw8iECe7tliaIn
/47HG+wBpPpCmuhIxnq3Sg95pFBvDI5jGs8gdE0IyH92DX8TYHrhTP1rAnET/Zzb
z8tje/Av1II8DuKJH3FizFUOhvXhqRjcdtne02X6y8dTVCxHmJNFFGHnoyAgf8hg
ueCMAlyHCrfAvQaqukhiSYNoEfOZrsv4/3EsI7bd37Gphf782mFOvXxMXJ34FsO0
o1gkSwryPOqGU2PECOOKq9PlHQLCAMfd9xV7ztxGZ+28Msn1+USYslaSkDaD5OEe
0ogLI+djMS2HSBCDj3CD8Rx2g3QZDiknG63svrqIrVyCs4aDa8Zhna1pgev11hE1
Lrflq0D5A2p4fcg7Chi4zOuA4b+toSBJbWKwZI2OW9VpBvCxURd/9mXuoKayCOZo
JRMB/VCj1TTcT5mtSH+idtjsSJ3cMFzVRAcKvT376o/mx3ar172WbgwZSsxmy56L
b6APu4tK3iYmpVgJsSqRM+sYxpw9GR0AA0IkpfhUJ23EC4UKOtfcKf7Xy3yzvn7c
yCBclg7jXAaun2hByM0lIIHcFoRSNzuQtdFedHLEok+ECDpGX4z+wfxBFndRNQDp
WZz5tSFKKFNr3f+Yk+LVy0KOmVrmOYz8eG5F3NqBsGEfC+bsYpLQeLgGxKCseKyy
Pg96QdsihBbynSHFnRSCv82HxB6LiFbDXHGxja1AZ4z56QSOc5KkuXmUTEEJzx5N
Gt82M1XuP7/D11uWcPSB/s5tMNegvqoiD1gOEPTA83Mp0sF245jZ16oWxDzRGHzL
/Dust2IbmzTokHr6l5+dDG0v5R0qY5ju8sTiZosD9jDCYuLapgZFdQS2jhIGT5md
tuGC2Rutfe5l9y4YmB1b0SQx1sW2IldQ7k+cHEoKkSXdCpOUF1ahC68KA0kKW+Hq
WM24hv98/04whRjZaiGyWk7Mi0s6G7+TrR3aWoabn3+r5f+m9GtYURMD0ccQ/grC
VXbQWuj7CvKrznpkGvdl31slQKuVkFAndbP3hrMKlgdVvnJO7fZjqaBdxWO7fS3M
hEp9VOAkLEpuhTxrYc/2o2E3IfgKU4okpFOdWjJg5nvpQYzQclPMWvP1a3fOgju6
qxYuRP2X0bohi+o4tnMStl8vVzYjS5SxGPgGA+Un+pD5dQFH+3IHFW8Dfxp5h61R
rG4moem++AreytnCITIbruY21DAukZcVP69SmGXXKfWrDX9if/3JDDvQT2rjzTxN
/MWNjou4++eBuzz9IIHJdwc3m9Mss3On5oAmhFfATuCy1jE0/DJgy1EIkm8vETIT
bSR5VQpkEBpBCqwIB4Sfd5PKTyqcE69i8nVxa5gCsOJtT/e0tDqpD/Mq8xQVuyFE
8kN0t2XcPwpiKa1HjdiGAXij+jRTidARYfhQst21KwFx5ZinTLqYNBvqXcH4YAP9
QujddqIqhKXfn12dW+X17EZ06m6EA5xjntJuAVwfbp9BAy2yn9ppPxC+hmSRzPsI
4JxVm7sFxOC54B78uSw1DAmG5Xmo/3CFSyT3ziL+d47bTJDxhmzKx0oYbin+Xh3E
nFuRQSNzqRjAsec+IieAHdePBtBWxfGFUnuD/2HQ0qwi8te9yhNhJaJ6sTBOZEFq
HYeorsanDIU2a2v/oYZ7T3TyDv8QoCBmkobTIieXFKs0vCzaSBHqNz4FRf3DO5rp
UJjHL2iCIqK6BFmrYyaInUwzWFcW+aBudhe+8r2hy8a5vO+v4VS7DVX4XSLAcbPv
fSMa8uMolRvUz+1O9V3AVzP1K7fUk0J5LtDEHv0WsTKA9HXckQx6URq6Z3uFw8HM
4fmIXRxnmZAdmmSSb10WXrsLW5loafn6uPtEfmjrd/RWqlQmp+fbC6iQ+rGRDi9i
GyOTuo9sRYpVUz+qV3Ue1O2c4t7ivervElG7r07PY1FwtXbW8TaNxu3zz57eFoP9
AVMcJ3L9ZLuC4NAoSZrUumENiY87l0aw4h095fV3Mz8WMnjVQN7GAZKqKc89gctU
lApxRMpv/+OKGoTiaNpqBXwn8W2H0MsOTz9kVXKD5igGbOEtS4Mj6ffDZJ0Zqrjb
L7FHxccDEoMaCGYsinQpXDDbouBxJwg6uNSnSTVsx8189c7usJXkAYHsbD7S4ci+
OBCOcLyPEJJKTT/KZKM3eHWfRReeYxEZH7ykVWHUYUki+RxJIBzl3w/QtghNAPsX
clGsG3vtBWGv1DF8NmvmFfyzKGiDWG9qYh1vSUEh0WGYu2VecQDz6iAz6SV/khXB
68thdDvWql9vuay/yggoKN82J8kJMp0UbUwVgsoABuPveVldrJzm5664aqWOy4rC
aNg1uFR1cJARrvw1Gtl3S4VXXC+nknKj/0NCVUqldOed5UFMn7fPUFZKNjSpYAww
HFdBH+9HyD8vZEXJv0RA/mt92ADBeICq6VnEC2UxS+WWa7hRsT7W85v0Q44psJu3
xehHBXcOqIlbmeiCYLRXMbSmZgdHDSaufJZLIRTARGTdFwC0ldK7+R2thS3qRU5y
ujY2VslizN2N6RSA/so/S+BXyOnbuNHf3qeqGpMbeY8dsM1sXjL846MuzoF9X55k
TBY4t9J8Hx4x5Q0G5NMoiAbgVZQpTV8zTU9YXSDaAeEWU6u3dOq9l9RVxpdTdg46
d/nUsQe8pG6QLpgDfFOIEZZT1iZlrXjWAQkKIsD9YGu7vDmcmHbc22WU3KE2AELI
93BkBDDl6+7VWd5wj33D8xdxy/JDskQbVYE3ztTGDh7Ej6wzJ9/0RivCOePPFIfp
sxLXf6rUeWRaIiKoq52z6EGbqBXxlyguuTUjePyZMtj219WU0i7tyoa9LlymLpev
tLRk3+JT7ma6vK9yWBVOfWCytcX34ph97dB/6rfmdByPXJLUbrSVZhNtgJ8bKH1k
24XFaQlPNBkfMo+cOmN/PXObCPMsXOgmvqjdS8NX7/6nn3RDQtg3K0aMYafukDJm
QhJHBDepuhlEiy5/0+YuqCUgGCEvv3O1jBYJ14TtVyxvOD9l+OkZKaQzWXVgkoMB
Ik7lxwvqqka7FMNIANzWiH3ZvWVjyfqF3QOnTHK2Zbq3LepbwYvWReOgB8yDAUiM
4MsrPfjnG3BS6FmRFWyNwrcqW9YelUaBgHGVXOTvh/J0RSavQf7Cl/ufXVrP3AXJ
KS9h3PU3sd0nI6AwHzLK8gfgq30UqVXNzTeEw92wG1if7pmk/+DJLR/UyggNaDmw
2fVKFuMpZgwcY1DkX23RddLbTuNV5yFQ0S5vhcZ9Rb4XkMrS2Gu2a3G9e8lDohaV
psJh4ylcKL2Jvc0K+KNmfUGtRsloK0nlkW2KO95Smitg7ldra6CpG3TXl5/d3bjE
jaFxSmUgVvywqounEaRwsfVHUfb2szxdWQi3Y/uD4tWHQGffEQa63n2l+vdpr6DB
LZVQiq52F1hUjC8RMNf9ZJyI18cmO/zAMT6BNY8RrWoXI/Tjdc2L8Tv1OaGwryIh
mhmuDN5O3SykNc+0Jc9e0li1KCgLzSn9kC9xZ3+vV4UPOnHeyeu3Lkz4gFWZItOV
SP0ZR6Yc6sTDkXLLxB+yhY72eC1Mlwn/VdwPA4/zM2myxHk1dQ44rNC15C7d44ap
TeVjPc4M4CrEGjaVAzzMAsuzPx0I1mIWgQb44gUVlkoKq1HblCFYhA45OgmKFe7J
hH2WT3/Ky7khGWaiQkrGi+O9RnZbDBI6FCAf7WeA+Yy4K4mQlQZrZ/H6tJdGqBXE
KpO5bg7rNSGHyKn30dlAp5E4vx5YEa+/igqCxvSo6wwYt0hdBrkD6/oJHpBf2a9T
RjM4lyJbH6771er9ImVeDToG1J5Mryr/ULwRlXjJqQvIolOqP2o9+HHiggA31UtL
gJh1tgEssPs6/mAjTF273kC3Mg/iKXo0Iu+3UbQA/odRzXl2UUE7dt4xSL97Ixk/
7s1LJ94jexD3rCuF0fY3srZToAGI5KKBwKQyBIRInYPoO5X0i0F0sOCzwGnRoEHx
pVmBu6IQfyeGflNxSPZnvVvIZi0DuqN5B4dUD/jFztj4e0cdwB5gKOA8anhgMfn0
pAXOHZnwAfzLLmQRiqq9Dyh08ZXhlPVVsxGiZVlDx2FMfbkOAfI+GDKCaEZbkl2d
9RRd4bN/Pfzqh1xYVdqlqX4JEETqONYWxHlKnkKhQxeknjv+3K7lcj0doT0V0mS4
6bhSw10k38HDuufA3nWXfdFvQepbyLch0EGUWMVwF5mhT79RDvLgmT0P9oiUh1Cp
2edaZEwGXxkTqS2u1lO9kFq2J530KGNkx8gueww0CBshitw1r61EfFQs9ODE7py9
+SBGVQ33+ynzLcjToy7a4z/455vf5vn9y6d83MWAf3hARnK+xVgRaDHKD+GF0OzF
euKXzS9Pptlr/7XptnyAl/oNIlPiJcW/rtW3XoYo6KP8cKiTeEB9oHeVWhNzHvKO
howL0cpoKl5kMi1EwGeiGYS08Fm2ecFUxUX7rv/YPtNrm85NuTKA66I+0hHfybD3
tCFE2pg97ptVRU+6OyoOiU4BGfPpEPqb1/NYDPZFLZ5wonbqZ72gAGQYB8jmnL95
UwB9xKW+asygWAeMBZ1wDL9nnT/EI1czjjug0RqpwCRvqAve6QT93pePgO397+SW
c64Nl+bWmlLehv+pQ/HOsnr2d7AdBiUwhRqFgc43A/zEx/LLyatO5+6L99v1vdow
3lGLxCKbUQ9cZtvMi7TCAFe3keKhvGIHd0cn6USvEA2yBsAxCBHwqhSqZ/TLebHf
MtrWQawhytNrYOxGyhn/PeJmlRkijK0lDbPN5Sf4wVnpLrNxMXqtT4bHvsIm2R3J
LW1JYqvNku9UVyZKtci4pOwzrFVvvxAkX4xLb3JgKKadqZ3Q/6ziSxgqOv7KFWSo
n5uzE2Tcu76XAjXrxf7OTDfSmfUaRPRnFrL/kl/Esh1E1RKTgbYljOBrvLJDhcmb
7627IoePAX6zb0dm3oejyW+1qwtDOiVoj7Lm1ZxAmJjKjhtyFT7Jlg7Bgo3xaeSs
3sZRk0LFiZ9VrPf6pyFkpN4+rqP9BcDo8ei+hAyiuShlZw8vfoP/IK923la+1IUr
O04t2ZtDIwVY24LxLxDipOML4bXxD8H8G7XLUFJ7E/veTikW9VGbxQEOACIVscM+
EjHphriwKoHbbgTvREQq3ETOGKabBknwJT8+Utc9H5UsOI5ZOJIC/r7ksg5hT0eZ
dwTFpqLbrFoZyD72UiiBZm5peM2M9Gk6MXX+iNW31DLT4YHYgCkj8YK4Ah7NX1hU
0uXpvja0TM3FuM5wUkb1ELh/vEuEUs0hY7ROcw2YvOarpvdg6ej4CUey2H8C8/9C
vdlgRc3SAyWHfUVKRY/tz40QxY/g5Y+5CJRe7jyDAcSYrZGbZ44aqxx6iGiT5gLe
BPC9kOGw2hLvf8/uOctzQEogeQBkHoU7k9j0G3uzuJ0Ql67x6ELkwReCJfvg8gSK
bjdaA07JOXQYh2ytieB1Zv0miRjzA94sL2g+PQJ6kvJxs10N6vnkutr++YXmxPYR
gnxMRqryTukl1LwN/uoL0HrStlBJhVbVjfMuwajwSBSkOPqu3CjvutERSfi7TsgB
NxiD7wL30IJwAEW423wpVUZZDT5/nkIIBeqhOWuviFTVKzfXTG6A3JzJappymAwI
VJptjCAla+3h8W1xv/Q7ftKjurXtk2kDnemdvWwLLmAtw8fox9NQFtVLjxb71z7+
MeGR7rOqxiTW9zdcM0vNpEPT75DZ+hEG2Gl1pk/9Ix1Xct6EfypMeyYItm5+fgvI
dX+8zau2UY4e7HE0Kmzuxtii+CYW4huP9KTmCnb38GRgTEz6UA0iuM4QjqsUhiV+
5cZ87xn46Zy6b/dFc+QPQ/UWvvqKmm3Du1Dnw2u5iSyPS2lApH86jTySsPHqFc1G
9UXSfgRK8SmHnrLjEQhkRjMjHF7h2GtFve6J4q8qEsXxMcsdhEyr7FETyasUQHDg
70QqyIxFMrvQ3H760Oyp/sdDHVFIbf/sK2bC61kAthobj/ngcC+pGv5cdCXzY8HP
3/AIviWDEnLdWsragD5YR3KB/5IIC3e+ogJq+6kOZYk84camWWN34sH0Wl8kUXKp
E93lPQ4ZSOAoZc/p0Snbi69k17Rkg8PNXKdqi+LgsONInjGciJ08BOE5y2T9wu1g
J2rruoQFdBTguAQr0anfK1T2gM2XqmCwt+we5V3gev4PrVfwOCKifoYCHxEYBW3+
tbaDBJ7h18cgz4efe8VUPPcvWehmtjeyZCcJlByxA6b5SE97WmeZv9Ja4p/B5DHU
E13W90Zjpute/fHqezNDn7myeCIhvuml38NUMWJKC4bWh9EzalE3Fq2TCvMJ4N1L
Ij4cuyCOMEqlyRdeiOcqbB3TP+nCJEtOo99YDQhUuI22xE52iI32jleuz0ICv0hh
6sUbvKMMBD97KYVo2ngDlLPIbiAvubL3XMJiZoXob3ngPRWN9f2llHSlWe3a0qXo
TINSy1gbKn9k1LbKw9sLF/tgHrch7NBix+C1RTFg5KqWAgjRT3zoGGG3PehEQlXM
EuApB3C0to1g5srFR0qQkVHhpHNUdBwX+paqrWgHhf1o/uFvT7LBeoTGTDkSy0Y/
fb9rM8baEPYXxtp07zRPvXV5Cxn8nrYtG/5hLKrHS83ssk1sRKPfKVrO+AV/EJNe
PgZtp1nuxx05lxACAirmimE0evLIuqax0sK6d/wOOC+27+qGFofV5+77mJVGNA84
A/wdjZQuyCF35UeU8oloWOKQJAwzQMBo963UcmXlObyvbbkY5Gdv3t9edQbonND/
GF6OrIEsCnGHgAnqMiFwPUvRg1zPE+e6wmpKDAYLWISYFKFbTMDA3Bpwv0hS1SS0
1Eb1j7THErJfH7XwvI10UMgH9A/lw+X1X/uFjHf5UgnvN8nqYRMnt4m6wIngL+kw
0OF53l5qqx4NfTTU4L1cRBY23/GC+5wZIOn50iEeM2uJ5B7/NrvBKzp6GieVz+04
Vv8dU3KJS6MfR3OlKZ9Hqyfwdir73honIO7vEWy0o2ELbSOOYPX2lzoZOq98zDL4
1Zru3MkPg8KgiSB0nEFlqITW3F7GqorAiIG7190vEWuNcbOlSe9Za6RBAGZO7HrP
RR7bFsibbkWZNludnIIVFb5ZWZ1oYyMz3OJQ5Xptc2YVxgliLVCKWzBlp3NjOUPs
YWf7EgkJEqyow3V0QI5sCf28f1D6xzWBymQA2XxW2yJF0ql90V8LUpNWEDkLoGS/
+Sx9e8MmhKpKtKdOakZumOGlkMVECT0/Pljte4Os9d3Y0ESudBwPRwiHppS7OuUU
7CJmVJdxNKMbvXqBHPJHtoqvOHLQo93HoUxd6XAIeOFOySCPFFjZmR7BpNoUOIrs
GZvuxjrnzPoXpsDQZGpvc2OWh1npCBDOHq3ajAfgJsKl6tReDvwE7J2E0hsfdltC
BAZrLst6674XBDewh21R5bUY2G593Kq6EfKUjqUmT1+Z057FXqbr1PWFLquOy+uk
/7Joy4ogaaKx+EsBGOgjSaR88Hq7MDUhy3qnJ5cQNQ98sfLEnegDbt1x90Y+3y2Q
tDF+Ogq8KI6o2xyqvc5wwr67aetPF385LxG15WB4HjLTepi9Kn+fN1XYxtGMOdXp
UgkFMM+GvnA/pUUsnUDwgqeetXNtxuqT8gN1yQEmLECRZnARXSbIETHHs0Ak4KhP
8ImweGINZkuIa18R8bOZIcC6KRX90NwXkKYaBc/oCueKZS0hJtL2UtjwO+npyezc
NTqy0q3zKvLHmZtEV1R6eD31MabFxqg3lEf9yk9SNHCDMgE4d90MFOtG/BWx9ADN
CWL5Jqr/lMuV/4nXDprRo6hEDNxVnLNnGd9AwXQb89ADkdGfq0dTcLKMTXN8Lhei
djhHAr3pxHHvijaMVczRUgvKgIXRIV5m9Fyf/GVaSqvfVGNJFCM7Bek42IrhoLIf
zsgr/mJfF7mWMgSdJmM9gsOSiE0Wq8vToslV8zWiG9tdOj5Tu4yWclBD2UJEgP3j
vEiqR8BGnBIyO9EuiOMRLmeyNzUuO0CbbD9GVnQM6pFJRFxIbvR9/+LDhqKWlWbL
6rVR3db4ZYZ/MNo9pdMrwGkurUj7Krj9eOrbwg6TvgPjb4cUKRHmI59FcjwHMPRg
slgfkgSljd+UlFoj4wGXHdkd/dBEcHuX+fjJXQMmpxx+bMEtEy0g7aaWem5R72T2
1y1YTsm3cUDYJ49Y9giirW7SkQ/ELZ0JR4ryC5QhLtR0GPoZxYMXyU8fmhv7tZjS
toN1rbKYwj1KXTO0VDkkrJrtyAbZGIimp0llTTsqTby0T84ExlM+3jzAO1MQ8NtY
3ROQgZ91PCxf1G2U+zGwNeyku+KFcJcf4zO28lp5RB34zI3h4pQ5chBRNX8524zO
3vkNu4nTr6jpKOskwrNxni8LcVRQjqY8g4EJN36uMyYJaHAnSFg0mpBnzvcPjt3S
K6m9DrzlQC8m70iwmWFpQq2wY3g3OrTQyGWwl/BANrluF9huML7xu9GO/H+Vs4Xx
KSbi+B7//bY8H3270UnBqfey82JfwLZJ+WY39Awbu3LWQj8hLumrdq3TEzpfxo4o
nBaShDEB593Mm72spx2TgSfGZRs3cw/eOa0uzE/bthBsFe8hLPBoKczv2GyNWUrH
YxVDzgaVkMBaQCk0KHvSvdF5n9KfwqtrBkWBN6Fi1iL+SgNzXDb0itv7Ss+kWRjL
/Yjq5o5ExRcLURzciftpHGr4wbCZOWzZq2b6nKDBOyuJ+4GkKs40r3UnlJYJ97Bt
l/UkdytwqbNB56JCXuxJw3lflIuLIMKUjRLJf+afXCmv3T5ap915GtvLl/BxAvMI
+JdK0fBOSb2oCOjEuM5RjXik1GWdGJcSVptx9H6x4WQm+PC0N8V2RAXBi7O7Stdh
qoP+d9Y7PeSLlr+ClmOvf5RbGS3J1hkts4+3j7QoloKOkz6KDehhRMaFWEYsNd7y
DfgcP5Q54sKRfEPWZkKw2w1j5H18YV1Z/svmtefntwsio2/NgckPxFBxIvMluB5/
gxiPdaw031FXRB0941y327dl7Z7SoSEqlRNumQOD2kYvquIDG7u6lEaIHgpdmfBu
VVOooBxzmqvMG8SNeTO1bFdCCBkw0d/yGkmbRc/xTiLAcEhN9gN3DE5JAfxQhZyl
fVKD+h+IAsmNGEtwl2ZfaQM5v8SP0E244wrZRqGr7wTn0T7gj9CcxCeRn+ekipy4
mdR+2M0Ocpjo5C50mug29vmNk3FH9DNpbxHusJjzNaKUF1Q9y7PnHhHdbYZy0jS6
PhUq8z6ClAKjdmpWFBPdxHEZJNX8bjnV0l4MOK+lNN2LiPQ9s9Dn12EIhzMefB8J
PgZ0vG9BHo/63MGRX0dmbS9ukPTcIl88wZ7nm7nz9/NIc6Bzou7dQOBnIpnnFGct
5Syc5/IzZr1PsxzOoXHgr3mTlh60TQw969jVy9+4zPCfFrmJExCsdyeFDr3z9ZDX
YJgyzPlFJU5ei2aX4UFCqWd3w9ZrJu4bpTRiY6kCb0VL199R7Nrm4klL6XA/uwDn
A5vPdY/kyOguRxlbUGNzLShRGr4LQSNJq0rXwofOPkp6wMX5MldI/faK38WEW68Q
XCjsquzY1v3MG+5nSpYB5CUQgg15mrxzJwviYTs7wFOa41O2z8DHpHKHsKBzHSXO
b2qRvfTYjIhQNi131ZRgWhs6n4+aBh+K+VleGEuOr7VJ06ERP1Sd6I3BLzyIWA8N
dPcqBOMzCK19rlicNc2F0SQ85HpFKw6+wdKeZ1HH79Qa64tOfsnPIxYjNH+iXUEU
rvYLYoSLpc/ICdB1Z/SrVabRRIs8tu6h5NdmdmK8vDeHMYlgC2MiifDEJygfUFFY
NqHbVMTZ5POUbRl4gNHbO80DAPEhpV/pFwzokhzZyQWJ+LGAxOpcSCbhPaC8Fuk5
vkyTvP3oPAexcI+DhCZj3g777YkXUHEP29OA31/dvr0lAulbzlra3ablm0yp7+cE
KY8+u67fiAqCk4s0lMZYtnZva+NfCkv4wNtH5LAnnM22Q7EQV1QB9uMPxtqWc7jW
u7C9o/7wM/eDkPcB5IlrKhTpSERwsjsZwKx+pEOYk5BIwi9zqkccntJHGIDI9cMx
/QQ/8nsNebeyrJvlvI797au9dQEelCsMypGQeMjLTfDjYJMJ1SXIE4vb9J1qPKd6
ybGoaaR/YqIYo/0DgTuA3P4XhKwbvbi4sMejOEc1vmGpCxsSDN03LaH96Ew1t3Mm
t0TQ5oDZOaHza3BGF2Y60CK9jllyiRgSewf4pXtCo0K27nNarbOWbBnw4oxpGGNk
vV84Mr5V6GY9do4azOC0VFvicNr4a/VX7fat4RP94EwSLRcAZVG6/PwVlq9421HV
HdGs2orheUOyoXQQA9oRw9LVGsmlaP5QZ4LvNkpjnfWhiDH81qnXxJ+Xru7ipQkz
5SJx2UIBQ6UqvOXZ9qVRF/vnEP0Kj0IR7DejItHBp9guo1sD0i8GUVoV/mA1sYpW
doWwKYgRFS/WqZ/9nBdPPS79qqlxefAkf87A0Mizf0mL/ZeQ1+Kf6J4pfvYvleDA
qSprNDEpS7ilyO4wZvY1ZrLNjfIwm4afvh/jnLo2qZvJIuHcOeSO+nK8550yM2bY
OidLCe2f7+3ORelNrnixU7aIycA/7iqTspUUooFJ1dtbNlk9c5mQRw4FRCvbBdQh
/G41wGJXBf4/fRFJoASZsJTWWc8rJgVzfEJmuevddD1SzvW7s4APi2DxoGE6AQGg
pM9LsDYRwsu2yvpPKoh3+Hv2ecW4wy21dUa/fszhovtdhlj1Ckt1iTvpojl5NrS8
iSMfYYYXZ42CEArrOvg56iuwdGKnUuwZBMcDQ/VEjyrRSmJikIWMXMsxHt/QdPSP
GNyUI0x3ciVdPsntOq0dTuVWoGGEv1LmPoFdsV57ii9ECMc2VSS2hyajDitQmIxz
gcsSSy9QD00FO808te25C/8kdkSzBmyakHiBWFOGd2ct168ArSxVnenVo4aFoP20
4wNRQhwf1fq983w5V1BpMHRoSBQ/Zl6w2z+P+PQ0HqpLYUPlJpnMYhHMFk5vVutP
UJ9dZUKmXVjybn9zFwnQInT2wZ6e8nzXEu3elf1vFyVMrO+LwkqNYQMBnnIltzJ8
bI4v0U51Z8I9OMnDZlZ7mRfg+gyMAbvLzaS7qyGqvW6T+YX6tFxF+X68cm4M1X79
2T5CDLWYirgB5X+zUIhyPfvAMFuDbcXwe/IE+tluLLclg2aTxA75Y1EBcUxw6+NK
HR/nDUGFIBFu77D4AioluTN5eKtZv/pdNHYEKvp+6Iof2/VTRnrsAtdBz6y626iV
OsG8uNHutr5aZNAdEc3Eb77zhH3CS+VlzLR+Rf836E9srNY0IRHgARvrHp7e+jzf
OqBx2xDV0Eyi0SSTTi3c2DjSdbsPI2O33zGHXzUh/q4WAAW48nN1DNWUNlNeyFCk
3mNJOEpiDGe+i4ZUdMN8HadcZRqtFBbG6iGR6MTKvGR5DJWMGZmtDK4cjc6ttfvU
KMqlf/4eJ0XD/JBKWAw7Q+SBqZFPsvEsi83oRgFvxbobUWABP/eAJ0X+CQcr11zS
se7iGrNcvADrIta03QtbGC2E42CEOW29cDyL7yhf5WMKtBpoiBEnBmfcsgPgyUow
3b+pLKq8Ge/rv/MVqZ1xK2ixsSWavr9m6HyzIn2VHjtoA8i9hE9dfgcmumWCmDW9
oQWMvMMFAOu4U2w3tNf5h7qNIUOyp6gnUn5fPgnWkf4PciFRYbsE0xGrmk6iJ/aw
ucN8emsLZ1xv1wsyu3PMsQ8EMtpzTlstJjIVkLvD4OIs62YcVdbwofbeeMWg0wLY
PBVWfuENp2HAGM42I1YBbMPJKz+q9qvdlv2TqhbwUggudII7bPT1OJUufs0JOngS
+5/G/ZzFCMqGhPdcnaj1t5qSx88bWqxpXQ0Bsf5RmQ4s4OZfo8KKqYXYImG7W6mf
LZY3PeR0qkvYEYja3bcT38qCxgqSsGiixpbnHuvNf+mU5nLy73YQRX1AkFdTzktM
mb2fmbJb6810L/9Z7taIueMvTTbSkVIVlnxNBpeif/F6gq2pNQytwexeFOLTtr2X
cgAow1qCh7LeJQHjeFpEnKKDF/EUd7wmQ/R7cF4JS9BYHYy7IxyMMniLssJ5o9lq
sn8Dn8o1soHpZ1AyKvnlUEoxAl82yvFQL+FxGh9fboNIzIpbfUcofXEGtk2Ubx2J
JvxeGPuJVdtP77jzpBOWwkAJXkfqze8/VeYFAUXxj4u9KqQEg7tZqtiNEVGodRaH
ojs2M2HJRWZHwjlcQOIYnWhS+feij8UlDk9drxD+/RAK+5aQmXv0tp9wlOl/IAAC
BfEoGsupbkjZL8PXoo4hqb6Cgq+7VYpCX+Z3rDOVavJ+sVNL0BKLIcPMFAJ51uLp
cAvmAO9jEW6i7BPNRnlDyJRStjKVcrSpQBQR+B+5OORM8ei5TCHisorz4DEtSfN6
om8aV+dwSLWzdYiWnorV4JZg/tjkMSHOW+IItqdFbkCuUJ6C0fR3KjnLzgixPcXX
ndnrcfYrQ6IJU1BS+TYNTImmCqgFMMbVmEwMt9OJb078u69DdUFwxpRkNSM6y2dE
YyDcg2DW+U+HrHSkw2ruNysEi61KnT26v7x7E/NH3mta4BnOg97EWoCsZtgFLHOW
1p6Zv8F6HKVXoKhll0nikyxGQnsDz3E6Keazm2R++DW0aXjcAxVCq7L+KjuhFV11
rfb6TFKoa6GO9r7DxByKHVMLxZhsnykJzajMck7A35e1s4wDVnKzZXmCTK00U1hp
0ZcWSG7hW7McpveSk6a0e9R9VeZjBix3zfphnQ5rdhRRQMm/KluzZtZyMyE+ZHT2
2QdcBtCPJHGJXTwvjFtMUdB6ad7fDPfn1Ldk5A2vmouTzvc9lsDvTC89vUtN55FK
WVxEe7PDp7Iei4QTt+IXZH0QesUC3xVEVaPuJajV+KS2HU8Iac8bgmPYpzHpnhTQ
N9F8cb0JaEEYG0NnvksyL41Fsuux2KMbwVXTvClI71tjlAmtWhlN+MV+3MLjyClE
tGuaDUqCawqoaoU1nWmIuXo4HTdrEoDc6wfjIoocdrzOV8+HzgA6gEPQfwgMUfIh
DoSW+qYLaC0q1V7fLdXphuzVaWIou+bxl6Oqo3nm89/jpPdVHqlcJwokPFhFHfO9
YuYPmzmNiTFKjT8iC+tweCf6Oqr4hR59KSCXd4ad9fiCTNl05U00Jp4vfBRs46ii
aW/RFYcWuU0pB5hvU2WvMvIfmNwEPn/KSclnVljjJdjV/IUXX5qRN1lXE73uUZHo
EKJQXC5/tw+m1OljX1dlmFP28jbei5QLyCLtXHst33N1z4LSF+AGLiJr79optTl1
JhXw7dfoVWJbg77TwCPVNPpO/vYZEfRd0WM2JILSKQjKLdXpxvZX233YchHL3QRG
CS+1TBS9VambP6njBj9bjh69KNt0RaTjJ2zO0D6tTeJ+iR9jyBgMxi1IIuWAjUu7
fgmYaQrRcDdRj5bSfDfAQw/xcP5WmO+vPv6OqhVFWB10k9DH0AoJwWi/fZaG8oRl
k2rvz62Dk+Mz2HR/uSOLAZ456mEoou1p1Us417KRE5GUmzPP4WTpBG5rQOBE71wE
Tz5Ylqp70+kkirOMA9bgTz20AGHyyy1usDRkTDr4QE21wHioW0O34Kw8lqXNYhv3
eZUu1n6v/MEalXP8bi1zJE/IJeyabx4mj/fSTR/Zt/N10m7vwc9VktXuP20Gfygy
LjLbQsyRVaejPwj6FmHNqJ97XcW7sdnT7cAoIZmZOeiW9wxwXp9QH6xztLfB4mP4
ebzLJ+LzC/QHop1TjU+uiuUnSzvFzHkrOvpERhr6i4YlAK48GdxaCavUPTUW4e+7
35QJ4vlNxGCQi3YhQEngcxz0fQWNo8aM4f3SkRmu7Fn+hmNPrbDc5+zLqsdK8Oqu
9Wr9RdpaBZM/AkuP2pozzbdAJmKCK7tUA8HoDYjH1sXtDcSXex8Sz6omzWSB+B91
2OnsrToORanOWxGwTCa2iCJFVZs0ok4p7/68eRJDNDuF1fPWazv1iucubi8KoD/+
JyJr+ALMc/9JWLQKhb6TjgKs9qPJo9xAXLUxu3qaM8+NuVDtxhzoP7FgGbP+H6/E
c3LpyoE6pWXZkUZ7l8bf9quiCRNeq+wuLx5dC7sbHMYD1zgQX9i+XjzTeE39QeCM
FDqt8iTxMPrNVbxEnZpbowYGHeE7RzEShcVWMD/gGpFEqF4zHVj36mC47g7TS8Wh
sWZlib6t6PEJyGCUVZS9mOEHwmw9OickXUwwcF61j179g4igSfJA2/BYeHpC6Tdz
atYNLW2slV84mENgdf+rvcwIkN9LVtiIK0M8sgqhMH71XABk2dITuwzpmEY6CcEe
LwH4ZAd9f0HbKaAVRD2rkWkfkAhzFwm0W4E0Og7+fjTi1BzaalrDyjhzE2uRRVvc
3t5PlfhBq0JTxMFKHkiMWC1ZMo/YzXC8LuWZWz7ji/ZzNLSkMeJ4wITC0Ak6iWkO
nW2ITWCuRi8Kt6a07IcPhowG6b6v+bdOE8F5Huzic7zDC3d1c+pEOGtYwTBOiz0s
l2D4U/3eu/GG3qNS4R4h19lBj9lmhIabf+GgVevtxrcDR4x9+kKT7UTMw2DFPBM7
nMcxSS8QiLAWIArMI5p7JlLflbsq3VDTxRPiGvghCztmJsHke/DHheLj1/kiDISE
TEbG5Ep9nWd86IFZZ3ZXejNsY5W/jh1EAnDfEZIjbK6CNEbuu2mEoiypW3nt2sY2
fX/oShQiTQ4XnbU69ID4YrmzuQggGxGJzbTJh3qL8AbbjsmzMsn4fL00ISiU9gOD
jPK6M7Lm/G3GwzlJb7nWT6H6X194V2Tymj1BgTEKcJMNmNvPixAwdaPTgfCVeQiW
rT/WHSlW08dr2CEHxpwriC9BvModFUlmHtxsRnHg+RiCfGYGLNV+2IW62WMYQRJ7
6G7GRhxgOufFwwHfniBeOM9lWEv3qyjmuEFqrO+bwlnPv66ixTKOwSXsRM0C2pIw
nM6GTBSxQzwYBt5w0Y8n1PKXR2VKNv4AZmGKk9lOhPwE7HmwjtVknASQOqDlw4TO
daDWnv/yYK3uYPk6MNneBd31bjaVKm3fMePEu/slHbbTFqT92hsOV/l7gD3EUWps
YnUkQ/f9T2BQPnnfrPdJ5NvyUYqII+jy4K8+F3q2gUl3Lf4IPznimFJkFfjXsV/b
lXdN3/HDNJtxdtavwzX9Ys4gGFLuehI/BAOJtaGEFM0cdzvPMtOlkfzIuRIFzI1d
ZLM3mEh2ZYNkWvUwu8BkkVhfB/tmKv7DO/ut9RNXzLvB1vt5GWv5pkS49XdiaSbl
Y+OH3YyHjO/AdQJ/nDn19t3iaRWBQDEM6R36tTJbtzuFgDGEMuI5ctcxXwXRFoGc
/ZdsezirZOdHfyVi+fMp/swPA7Bmg4ColFp74K4hSeBym25a2FwRAS0gFhQJJcQQ
Sgte1ndHH4x8TxdzrNJA06pK/uh0YANq3Bl6mDrQ4N+pXpLENEYHtws+uTZPvx9A
hzfm3TIevcQAtxpWIK3+Sj0g/weZbzBNZ8/dRinooTvh7dsLZrlW5F1iyr7DpTd0
dc+ZcpcX0M3CwFJxdWJMuC5XgaXfemMvxh7xscPfGAgcfMbvEcgd7TaBq+0WO3Ik
m63Bns+Qw1ndklc/ByCxaTSKCy9RjVyl0mDgiP1tp9qYty0MXncrakzPFcwT1XHC
0JRwL9UGj02sQqmKe9plzeAn8cEo1cv1Fkfz4/EUTusbOkg5AkDU7Gsiy+r0Zbc9
/QBBtpgwUfqZB7J1glPcoHULfGdu4Y1XJx1ngX5T4wODOKO/gb99To95pURSGHjk
EIsw4u8dCaVafP3a20MdDGIruy/H4m7zseEAa83jZvykLwuzKkIBhjMnkjHuZzZP
OKcpP3wxvgZoabdZLVkQoTcZ8PI4lCagfRjmn6EbWnYY18Ba6CFMkVzIgi9u74Ho
+nN1Q6Vnblr7oLlJ+arHI5j+ei4S0gdf9Icllnr9qmWfIaO/W3zWPUbxcxGcZ/xp
SGX50SBZv4CGBEhsup9DgVx9g22f9s7IdRtkS7/as61O4UjStffk4yiAVR3QfJcm
n2q+ZgeFRbi8eS+KahvZALXQmRTcZD3NFuZncV4H0vadgkcIMpjdcVfcFkh+R54R
q2wlLxNAlu9CwLMgWgBThF++263HkLkTGAeQK60+TfIDBTzNMKT0vrvfaWvtjzJJ
t9mn+US2vzYRJ9KY40m5Sf8JZ3X1RfsVBanWV698pH+iCiA0Wjz/A/s0HWPKGJuP
yjwmZJdcsjUAMEZjaEjqUIk/77K/ZOkcPQk0kmqz5/Zf4aLmP7+jANFpMiyT1d6/
ZSNwSSNHkfBT+McKksaP7KibO7Hxzt5VClB8ywyarbLglvsjfnfW8lIq9stg94SO
6Ugj3v4kJU9snT94IJ/KcPf12fDJ4W+kbyKdFzk5slYd8/kboA6Fphx3A/VM87q6
aU328fDBcTIjj5LxAWO29CgtBg7CaoeTMzZN9MV6VPR63EktIsHt3x7yrpbgf8i7
cbZPiWnB9rDmg278lrmJg0+0xrQO951hzgXtzgv7iW4UmV/9Orzf5bjnTvXE1t9r
FQuzSVbvRxvhmPAVIAX7ZEjrsF9f9v7SqYIsi9ntt7O1Bt4aFjHvPcTOiJ0IiI5X
s1zjiQbXA8OWULrCq83cFhPrsoND/VgcghKrj7FP85IzooF16cdavSthF3Zwlz1m
TkVQoLHjnW8QQD7Ln8ChwUUCfoeqX6mAqo6VnuhU3xreAw/SlOa7Kdl2bpKaRhnb
iAK6YY71430LQBEqo6H65ER5qFAXz2FfV0auAfVSMNAam3pxe9Z/MLtSCV6t9fe9
VH2EvU7zBUZgrdmTxgOxJPRnI9xPh99EZ53lW18FlM4+SBTgl2fmgHp2Pbsju5gQ
xzzne2WFfgqX+ANViYdsExUzxdGAgXsSucqpjKvndmswVSqmTnZGVLxVZ8+upFsp
44gdj5si2YzGxRrEQg9Rno9iRmyDdE/4O8349d0RSwVw9w6t+ULFkPRKVzjQWbaz
M1oMza34rGPFNz+SaonVSvjpmiGkIUJoNJcsZhsgHPg7Yf8FdmKeWrvg4J7PSEmB
XtM3l+JS76w47dD3iHVnVaVeNdoiUWbK+KvQlMaYz12FNsmVq6p6gJ5WJO6s5LfL
Xhv8BJPXWsdGl50jFGgVpegmLlurHvQ1WOcDhVKVfCo+Y8eD41EHgh4yadcfN8+4
TYJO0r5Hxy+uslVdGVqb0YuFWneQ7/RrOxBn+2vgL4HuJQU+H4UjKLDC5y5EOdI1
89UfsZcXK/IkROcQmcZC2yKQeDCBZcU/yBefnPqvSYnYUBGC+TVAPIHvlaGXJSiM
IidIK+sJMujQlEHwz7jMT4/1NpiooP4TXd1F+1gKwDHSdAE+hhnHd6xMaBnL9cme
9Hhw6vTQbmnPZihrrj+dXRIUQ75czA92pa6mIgodAzSk8yNgA53TDcwfqEnDtjU0
fSBkx9VF+1r9n4oRUMtAEG5LY9fwnhzs5iKHEgG1tUVw+vZV26+9p89GLYUdh1xN
gkXTyyusGka6kccA0w7VaBJTOpC6dOIxuTpO3hqXNWxHAIWoveWJMz9WmlqPsmnC
1z8gQTrWrJgqDmYxJ7ACmb+nBfFcLinPbHoIxhWzRKjhGTDyjHkchJyFi7l2A9H+
dDAbPdVKpshYTBQih1nFdq1RHjHfmkaIuLKUHQQTJY06/TWL9uC+UWmekcEU8ly2
VRgw54ZBFkclrEbSivLAXxcFRnGdUl7hgQsT056605Jz0SDuz0jR82O0oGAmmqSi
Q5TN0kaE2YFXrTtYtocPRvXGCAocNVtlzlo6qcLq6Brbk4drKbV9zxBovSjV14bS
xJhWK8RPdhiOG/M/91ZyPNELFH4TUqI9fdDw6Qt+aqChAlmdkZCXHbv/IeGmkt7f
7gy+Z+Df6np93mXib2YSIDg3cIA2cq9E25HwJ0YPw/eaNfvXMxNYH53+7+EYKRiw
3cTmRWu7e4JtYezBbsJksKM/2LppdKw3q+X2RLie9dHIoKfd7Lp89jElyIyQ/Utn
56KzuIEG5ZZ8DIFd3OOzplmK7Totq1PkO8LrvNuCIJjk/FJJeZ37Ja/Xu/5bzDZT
zvUlebeYywTPLV2OUCEsYZb0aQ1ETL4AJ+UJC+AbGbpV7kGOZ93ySGTvh5Me0ZbO
he9AdG5OFwlf40YpZG1nQuJmH4pRoeKvom8vWgdgWuADIY8eDj3HVHDkLUWXzuEM
4uB01qyNibsBCi5vyDQmXBiUGXZCHLyGHC/bKBOwyj3MnW7EU4gZRN3VOorjH6j4
cOqXs3wHShoSQrV8nFiaGGbUDQCzxTnJE8lSsXL2y61EUNsfovKDQkOhBBmJZ4ip
9ci5YR+5aBHG7/V9Kh7zeenxxEYNQdzW5OmotIxfOzQvDOioanuZ3jxpFiA9mefh
0qUNoII51DNJB6dKh/R6TGnWQ2YZMSF96LEZOhmeg4VoVN5cFQuwJv9zEEWHDZRe
SQEWH/7/T/XU4KBS4qOMZQdn9pQMSrMKfmQh8xDVB3jjdDkNJbn6NsBj44yLufvx
TM7WExm0lLDZR7PunTqN63HL6Pgm0br96JWfpnrJbUCtq4YG+9jNmaqRwwk5NIPc
y4IzH0gQeq0hdzg+kW/mU9cOaXtNYoMdl7SRyfhaKF5g774IZ8KDZc6FVDK/zagc
+yUCywfrRyKvMalM/BS4KAu7isN5tFSRXpTTCWboFDOyOs2DgXoNWGryzomZVMuh
okqfSpBZOVbZDwmqz3WksAKKKJT0C+a0vSowsDU+yuBBw9tv/T6Ra8I82sPQ7Rkr
IKytz3VQ7CMHoL3a3KYPmGZUDhFLnBzwxdGvY41JtKfvGJNFrlKKNpYNows2inAJ
j6Z4oi9IGDWTpYDRDIjqnBvYaAXS4aSKVe7nPlJo+RFk34Kfa84qCAMJhDege5dP
v3y1pz814yGcPitpkXp9LTetyGqttcXIwdtmLanRAIrnyzMzYVSH1GcNNu4MyHMV
Tq6UiMA7CrjUfxUHoe+kzWMUqKtzbS4HW5MELG84DPJAE8LfvgtUM8TkAdeobkHU
uMCGDNEKeu53jorXqvZSaJDoklAPzLCYpn+6zkU83Hp+6mZd0Cft3H+ulLtHjlYG
boJfZsmLoUaEXfa7rIWnh4RDdrP8jCVyWwsXwSeetlAzgPhiQQ+Mdjhkj93zDCRB
A5LVZe9VD+nFKnm2EaXTUIRwwo5y3BQz4Z3CcN/k+MYKEHaWvpFp350/iw5yH4+v
s2Jpk6zHBIdNgmJQNjG/BDfF6lIdq7yBagWo80ravhGqrLdCgi9Dw2feTtD725sQ
VJHg/VZpwe0y62EC1TVK7jc1bqVXeUYQmBvGNdDioepQBcnTXc2E24Vc/Djw7RjA
ZuOcDBG686K67eBZH/baOkHDLzGnyDfR/wm3rtmSX4KPazHxAKsmJV4jMo/1sHJa
5hdjP4DbCoIOPjU+k0gcP2R+7bmRY1OfsAWtSNAki6rWaOLyxZizL4xkew93Hlgn
vpmbNQb6uUQaZM4eYTWY5XjSvJEy8WDjVt7TCwdOzUK/A4KSPmbpsAX1x0J95d1A
g2oYRS8zVHz1gXsn32zmKpvJEa+MHHpXiWLckQ/s7I5fI+EbgdxLMYieN+YBogTJ
6WcsVKht9OsbH+80VhB0aX4pVswWEkODp7SOAo5BUmkiV9BYPcBJ9HdmrL+h9JGV
reJC7ooAqE4h4CTIE8MMNNplJ+Pw+0GOwmfWvLtzx96svoyo3Gvj1lJiR0SPZ4oK
osrCA99u3P7K0HWZGucefHYuD+ZRFEnAIXi6KTvHQw28KbHoyJLMJDSDGcyzrf9j
vMWibLII58gNj3FpVlQpCgXcVyaYeV08BFcxb4Wby9YOUKOV2lFyoUvhZu12Su33
HcH1/YGbld5p3xRGzt50zXAiME3n9QOADDaTdGwNk7L/ReEa8nt918JgN6TarEa5
6CrfgZSwWED+5VJiSFITnAU16u/MB7rgb3rL2i1+WHWQ7Hrkefo6ZjFjrPtZiJkm
URHqduZyLUobN31QC18SRlqmFNrce+ZPa1d78dx4SX0D97T7qitPW7w1e6uzZLoW
sqdHs5Qtb0gerewBf7f2zCvFw+m3lml4ubARHu5dkTR/YbRHbu/Y6e3mJN5lpGQf
PfMXAMi809cgeEekiZOM465MFrNJEVwS0DLIbBAJqnVTwKiYkzfJW49Ue1Bz8d/5
h9fmtWFtpfTgW2dj14Nt7XARo5xVWsrhKDzQho6BFcV1bY4awYBSyguiL1ZW4bag
ay5idqg5AumbhlxaZmmhSlfcVjsK28+NUJBMCwWynA+9+C8OPJjon8ccoc7mq3Vu
tdiwahe9HkH4tgviCuai3v+yvMg9Tfpm/9OXzLqETaPzhLewLZpu4yUrjRlFcqmc
bhFD/w+X3xYNrLnCD2YGlhBlCshPoe7OxgnyyjmJwxgnf7OBuTheT4w2+lp4rV8T
Wb2/rQcQVj99Y06qjZ1gdDWAeR9BxC9VxHEDK4k9UIfdc15PR26GEsX2qxwLQtzA
EEqAkSCEnUSuKaHa+iENermoM6VpqivLhRpekWEdsA3Be2RhIDO1GlVfVlKaoGvv
2sq7xFNCeJgP5RI4HcvapuuC+R6A1qAT8s76GEM/Yato33kClv4xYlLGWRT/yiZE
FQ9KIjWQD01wDs15UpuKC2NvcYI35Svcsv+h73VWyNUj0ulkOyloK35FlXyQTGTb
7a7w+mFZ2aNHaNIJQ4bwl7MdMOhg6UoleObq81sV6qMRYvOmv14y2zbiTEADMcvA
cVtrj5fhaSY65XBxJhxtJ/ttzHM/c3LO4lN8mgsyoXCkLlmC9LyK8l9M2t2pNI+D
5a7ZSLEUBB/cOBJEukWJjvid1e7lU/hTG8oRZcBomdvpxfF2tdeW2BmRNmtoX/me
E6DpDWhXQGkeb4JLnB4bq3pyJ1+52VU1RWIx8yv4Wg0Bt0d3+y42zTZ6DdkQoWow
3sqOLQDBDrh+mD451aie/YPnuGduDi7VBzxA7hqdQCbHos84hIy1mgSkFkKe7Z66
XiFvuk5hvwXj7pZH4BCX5ZOP46wNEUkzldMUvuTJf3Sh3Hj5hj8PjqpWiD4wsQt0
2yVQmp/OaX3KhuLiYbUvn04mIVCf1ltXn/uhRTnveaDKw1UNT5U10zG35GBfVB/g
GxtIQfdxOFHjydq7YdZlXQOLMHnm8wG+GHXKqRWkBDt0cvUlLY83L/2LKQgi+C/R
jVX0W06AblzcrnHN4ORt3/s4JyeQlZyC/gWpm5h25KlEPAqdHN9N0S568sA4FDoB
2TUDnB+duqP0/bUi/phZPcc6eojUQGNd6KNGE61dewbJnWSsjCB3YVbV6VuBhWly
LZ30zbOhKE/JIHOlbCz7Xt7YHbcMHCJKDuciiGjzpkPddMoImEn0CrDp7fUyQxhb
py1GWzqKcN5VrAEWvXca3mbUBsI1wbyYIcNK/fgnoKY6mffJaEupScjQJdyACBSm
rAyrwOVw/Bc6wihxmlf4NVYudvwVtJ8dB7gnSCaG5Yp6BdjlGObvCAVESHxevE8J
qHU6Fu5g3OeErVtekBGvgYm8/JqntilAIYwvEiX8g6r7fSHACnD4GLr0DELnPNPO
/k8eaF2SnHFfIIydhiZEL5KQpQCcEiHGPjsWXeczmjjUGcTqyTISzDa/7bC4EE00
XqddzFYJ96pjWSNjBVrbfP2B/qyEfUclgMryI5x6Ffumj+llR4EnmZanzZCrw8Ie
5EvEVH94yjrIgyppThwLvmuDqc7caeGt0O7IqwkYIoIZlxkoXila0CgY/R4y/Oc0
Yw48hRFjW2hWq+0emoWttVVBUtcXwSULPg5QHO+CTmlUXN3sTd1CZHwUq3Q9mxh9
DsDlSMBrm6edkGBUfRCPaZqKgqjDB/U1BgdxTgTKrI4jK04S1SfESG9ctjc3o//6
PfQ78cwoqxsQMnevgBssdPrcGTxbrmvZjvuWLfc5zPDhwpxCe4wzzg0fVbRzHafF
An6v7YToBpU8vXXwN6N8V1yP49Wj+/XQzFQKrPwD+U5PuZdwv4+uV7OZReyD1BqV
5tKrFEFFeGSbcMPW6+kZN1e8bL7pfE9RlSsTCaG3dKBmtsUVZGedWwVhLOOJ+13B
Nrk3murdmgKO200OXGTea/2qHjkGDvO2VFT17rdahJrqMhKiNUsVJc7KM7Pw1bgd
o1JzHsnTYgKrjs5rFu+9rw1euk2EouHSAC3NaPzMPKDlDtIhlBHsAsyC1eiFe+xo
hTvHZTqnbcEK0HWXAJHMd2ilf4K1ycaFH4mnEvw5fmtY8EMEaiFOy2dxFEBXpjfW
1LCp8K11tQVkKjrDZfXbsQ2O0wgAoyNmv910p2G01rIg7CET6I58CsUR2Ry6Yh9u
CiRpLgN+GeCSMUozD+BHq8ffZCrqxFqRv3Dk3aX6d8LsicEzgH5bEVM91A5rjRFJ
S9Y6HdhzWT8lQMv0ExxXQLKcN6QPiQ3u6AC04DGSLN1S+peW/ML9JcWN7ll1KgAd
KTf2Qh6WiS9Y2VGmRnzZMl1AdI8eMw9Z+qR8DcHBdeQgfONwwcavhApFTV6i+kQR
UWnf4ae/zZKTf7PhKI5cds0pX3bDH6JMoOqY6jy7Q89qSBo5f8OOF8/Fs9ypaUSs
1/lS8S0oMgmqHlbgCeSgF8tP/9rXp3iwVwhUgcwCSM5TYE6FrXDRqlPV2i0COUQ7
R+iEBuf/iu/MIe2Aznnau9KaJpWB7R3eA6pdlDtvuh7UDldLMUcn1moM+AzUwmpI
9Koxr82CPYNcPd3JMXKPQ0JhhB9YF6wcIlFqJ77FLLMkSm9Q1uEy73a1IZywBNwl
sLZLx1rs3Wl40dv3f+pYK8PhF5z69xWVfDlqv4lZoFOJnJW1/EMu/xEaZLtS8ehZ
f2qVnnxaulKVc0iSwQuMsZYi4mQmjVHPXBIMgdOd3XNxMce4buged4S+M4e+l984
IMnTEqSIxLTjdSskP4dPed3u+ZSa0QJoEcqWtK3Rvy3nyobGN2J/9Qv09budWMR4
rfHIHPsmSNlrwjfOzGGneWddU9/k2LahkFougUNRK7soffk5gCDce9wZL9OrR2bG
eJZ2IoFALpH15j3Mh1G3vyXu7E6CnZn+XZrq/779d9lLGJ/IiE8O3D5jU6HmMYXX
zTjpKj3HsTuiU4exgyqBK6z8rySZn6tRTsygbUjlEYEw1/FVlr3mNVvL//srVn5O
DPJ6wfBN6nwOUIkL7Xm9fak6/p96HfoLL0jAwgR+2T/FE4D1TZtZDFziK4l7/1bi
QjUa7PJfwI27RH0MX26SwFtuXMHrJNo8K/90+/DCkgU6/WxGBQfsJsd/bYuwlzUC
1Wd4mX2yDTCtYMGZm2jN2FSRWRnlYQSFc3W5QnmsrYacHxy9R2i4RKteFayVyxV3
KUP/2cXK1fLfCeGhPOxig3N/V+L+mOGDlxXJRDeKbiUW/DX+Elm5Cvktqm+g5E6J
jdeScc+vJ2PwFtPEtJARZJdyngrfmY7w8OfNAD6ztFvIdOiQjNuVHvULBPiZeTj6
4SRO5zZwY9tPZz1TTDectiPIoJQZI7tbOj7Si9JiNq04D+tH6xrWJl7OnYPa1jCD
q1VEp5ogPk0IBkEPk/Ax9A3L5LdaDzc3PaMczzS+vH5Xc74JeFu2rwzWWkuptLRg
GTzK8syXNrafl+FFf3XXFGml3T3Rr/+mMo7HPqkxZSzlA8iIL8OxM8kWO30QWmGE
vCoPbehxkVI6fhDrxXYS6v8+ABUoPvQc+qVIZqzKTunZ3SsZMRVn0eF4sYUESc37
ORzUzDDg90GbfGnzMHd7aV2dJcxBBGnz+hpzGyL81fDrYnDCrvfaAR6dUhoAiewl
zOYUDodHEJsPivaa/3eD4wv14Rwpunhj2PvJ8NQVJjgNz9MFb9/G6EVakvg4oFHt
hu9RtHoN+QJ92l40AUkl8Y3psC2km4lY/+nUDHdLFmC8cpzS7xUrhxnEp006DYoU
/iBvE0SBFY5ojm3XAOarPKdzsaJw6w7H3PosOi0qhZet53rNJzkbZCqD5lT+CvLI
T0UUGSTPhzifWBH7ZdFsyunZgvkh7lvYVvyXDcO8ADfbR5XIkYcOpIZ6DB8yIWeO
15oovwof8NbQHy1fe6tvsU62VmvtSB+USz5X3qtG9CyFOgJPmzDmifCAed9Q9F9I
mjIYdDxzpfKxUYq3VsZ4Votmte/7/VIa8eQVSsN/Wic/+onNRjdYggoG5Hx2t7md
FG/c8S0FjwODhI62l1nO/X0r3z2tKwhaXcppm0DOAp3/ifbhtNG4z2R7BzU9v403
1GeE1i6LgYSNoq1AuDo+lxI8j/EG80CeqIGmBR/lclgSndn4Oy2m520V0FTtQ71p
m+s6NoyAHs6Oj90DiMgyNTeZmgtFFwnGMNrO7tTX3+t2PW2gVvWiYCflCjkVhePG
NfPkQgArPeJYc8/1N1Y/gUhLS+QGFazg9oQ0JBTgy2OOjVnTezYGsFkL4m7xrOaF
OWQza5Ktjj1a+8JCQ/9OAJRJpfC5CQbg3WfG7P0qb07Jl5LK/2gvGjQa746HNtGZ
NkFmCw5um45QPhhcfXQyV1cSTZH4Nm0/j2wCBtCE/EyXcqTwFr2hBMlIIelJlHF5
ArfSgVXbAvKhcARrtF1d+E0iie/Syjgt+502pYxNr8m7a1wcdlwsRrXDUe9Yr1MQ
9himTfM09oHOyUAHh2RaDKzu1IYnyfyFaSXqDBhSm63nl3k1Lk2uUykQIasn+I+O
UWTb6n+nIG4lDzAkE0SiqdErO3aaKPW4Bgmdb/SvSWvFh3PqxIIgt8n8bq3YmWaD
0K69CZz0P6YyZN/742LLb73U4J7+Oa/wHadookRezKm1T09JaZ88kLFiWXLkiYQB
cUZJAjkOQ0jGJJCzJdgkqcilqMgioIr4fS56RrGR8cXP5WenPdCzUJY23j5oZoQy
SDNNCMAz3bCjqsxTVi/vqyRgu7BaDAX8/gCNrN4wBAE/RtRVvwRZT+Mb5TmTRYYM
4p6e7eqdQCAnGEQ0Klv0Ntr5s9MAhv5mniPeRefvOj7g5HATqdxuyfS2w1gPGWDL
RU6maLzlQCa1L1+AvbcDndgrCjBne66eawMmgTYJbYJYycb2y8CLVzwQqkJEjdxm
hTGhPDvPq++VPw6XYqnW6/GTjIgi2g5hSJlam2fd2h+lBQ9BiNt4UJcKp9H29qFt
B5ancNmVZVURwQf4/toYGVTAit6Ie96t4EaH3Nyt1N9Sqx7QsyTSxx8mRX3R01WZ
lehNmnmZ2cVFB11HugTmQyTn7E+mtqfu5xv49FLaPxVXd+nxw2CYePrZC2v/6DZ7
ivQbXifiFNp8cpb+Bx2YZUiR4DrSlhz0sIYwp5jIuDNZT4dwRoLy59Z7dwhD9mXt
5ygQiwTe9+plNn1gEBLwtINtGuD/OXniCu9Y2BLQDXZ0Lkg3ib3AogB9hlZl0RNl
uUHyF2gRNBNJJpgxwwiHLR5WC8MEKcwmck1Inoa7ImXfCWzLGxA2vDspJrpEkSZb
nbdDjdrk3ep7mdE1xKhEYkrDGCQ8uhM8B/4GPM4FlW5MK3tdQiVViaTjXod6m3GP
imna2MClbsatkoRb4C5NiyyvfDplotlFpz6Btd0pxOQscJJqe0cbZvKiYBKZV3RM
xkCK6L0B9E5o7TOSBc+MiQlzF/0JOTuU+nI7C+NOXqh14lEROpdyCAvr9uwnTeuS
DdPfmhu8d8cT+jyKG+ptgSlwK3Y65wmRwJYavXoL7vxFESAD77nnv0EmcE0Lc/vf
XB1ZVuNNoWFhpzI8Tqy9o928oVAI2/M0P39cWrm1RS+TZhT5XYVruMrU6chlKvhQ
QHt4rQb2zjYoYCOw6VAHu9M4g45vjAk791U991GFAZIhqPn17NCKeuJv98VCvpFC
YboE40xXGQkYZj6m5vxb/+aaM9eRqlEijpa59m27Z96kJWHVatdbPYPtEFGFfG8T
Ia8/VkmD4eMrZH0GDmLdscgw+23EV2tcXZSIyu4hpPaSWbm5NLZ25A5z/gfakV5I
kkbzfP1XSt3vPeC+kzWkV2d2qUqXR7Qf/JR34WUxR9W9Z4YOg/dFnmxMEp+JR7yO
Wpl1Vq2VkyX+cjeB0Rlo/dK1BpElnP8HueJ+fMEEjNW6JyG9yppMOa1ANwFiL7Nc
ejELIZfj+SdjBQM/oxl58Du9BEaz4nBniuvfLkghibnoqO+JrNpbClAuD/ntjZzb
mzfGe3khRiEw/THbv+JPQjPOsYRlRr4PDHvFydSslVeui7iqVBZuBGBIRFepKg7X
kz095tESUYn13jrJmJ5L0rK0DG53JDo1bD0JtnlZWcgXGWs7jJWN5TFZ/bkf4Zjb
DqwgrBrFxXG0YkaZYlVbAvIi6vwrEoqrd68fULY+QQ/pwlN26eBNunF8tMBMO9Ch
Oktz/i7bf74mndWeTBCTYjNiB6eR54ZbW4+7AmRbHAgqat39txP9qo0cjP29Og27
8rgHzavOEDRn5O1Ku7/MVDiVJEqALUynPk1JxesxU7lMNM3tWpe6rTASfm/uikUQ
hzCSgim0JHsAXG3fUMbdY9m8JsnDNxD33KAZXK5rEOJVIPoiaOmrD3YR0KPqpaDr
jThXW4xSH9leiplNoJK9a8m09sD9vMhsfa75txYPeb1pZSUfgIU5H882FYwhxIBl
mQ3E6fGcu1w/XB7NkyAwAlROItCM9Q66L/z12UpKZKWVaWw4t/Cd7fwaahUBKb9c
mLCjw9Fq2cqSztC73+T5ZOEKlNx0/c+lsTDcXW4kmI68EhkvanclAJeD4ueXN429
cON0StYZDOOUxXZkDBVLGdMfJStJ1mOcbM9IuGhh6+jMsP1srynNB+ojHZDhDwqq
hyT70Me0xQH72qDgTmNjxFq+d97j0zxiuRUiNuNdl4lgPjgZ5W/V7/lCr/Ym28J5
riKtaq34a+Gp/onqGpEhXMQvIwtUcQgKMLnR6Yi+DNu9Bkno7dJVXUR0dlDHtLh5
W5e684JBfY/ALL1xFnHyKWBI6t6KyxuoEJuVOfFHTCGUxYBAGbpWofDPt5KUSlpk
ouH/lnPxw6cNAzPKANSKTSG5qiYf7PvdRSVO56pvDwDmnQEWruSKwwWA+i2KsIgv
X6iabxWZKu3SNA5aLRkl6UnwWNKEuJMmpwN2cwqxSYjY9+LpTCbEG19774Sje90w
7f7ZEI4ibItYKDbnrDCFoP6EPDYk3wnZQvblCekc6mt3+FOXU1XWfseB5fZJvyxh
tDkQqe6eL619RKNAI20rjBeMu9Zb4TSWchGmT1cNKF242+K557tX+x2Cx/u/3AOa
wkCv1pd7OGr4M7Wfz2oG9bsfS4DziOXRXb7iGB6TPvFr55/UB4fkDeRBH0j5nTGj
sn9xQcN5fbq1ne8cFWNXKQ22fVNqeynses6FnovAZS0Y20zN+HItNyA7mZtPiAHF
A9uHA6I//46wyyKTDjXYmqMbyrY20oLGT56XK7PmryYJnFLpOMENgbOm67vrBL+w
BmH2IUqt4w3RoRZqHdi/66y8uS7P/jAmyeB2ZY9O7t6X9oJtiS0OmNAbpXuFz1Hu
zkgb16Wtgwq244+dTtmKBVJ8cCBy9CahATsVB0yUq/hXHrVtnRFG1eWrNyAWPGac
WzaGtI4/qa1jy3A6v4c+8FUE0DLklWbD6sWtgw+EFkzPHFiIksOHfxWrKhF1Fa6a
S3G02UX5GPaQaxpCiEAKqAdIgzfv86b+Z3Io3tItY6SOQ+Z48HmCqF6taW0AWkg+
BD8Ie9B0EemBiG06CYklHY4LIk0xzNRXhwctPhzk/GFRbeeHvXaMs7Vwba1xo4Dh
d6QC6BebsR5+2MRl8MD+LyOieOvXaxu6aN5u7dk0r7t59VbkiOWdbnqxO03uSX38
YXgF+w5k1vJhqTjn88GOy4wMRmphbeFlDCV9LtKaP1Z+m4KFrGqy82R+lKwyLYdv
1FnjVL9dBIaweKOEEkk31u6DIBQsWku0tY81WX5GXQ4JAEH2f9mXzL6eHopP/jcF
2ZjyYnZ7XY+4jooKbK26bbaHeSlgTGnXy2mQW5DRNW6vl1QiuaGutS5jgczesG5f
KVlQOQ9xyx4iWer6fQrgHQuglALEV6TCcPe0/AwqrIw1Y1QpumX3AsccUZkbSYfw
xrYbxxT3AWkZIlpVrAZb4lqxUgLSfPlC0TRu7e8b+8zTTCQtxkWb+iDpkSSkoTmO
ZYBU6VV2tkkznas8KzeN2TnqnN279OWT0Jdqb5ha0uJ9nBkehjH5L68AwZqtiLLS
OzbNiECgyo/FK3JV5JAt7h5HdR8KgFoDd4AYdzfC1hQKpskmCnUr9cPdfeTlHz9i
REWMTyoBLTo0vXjlrpE+A5/h7ZFMGbcSIIllUe/K0+7UXsfmCsICuMh1hyrYOukW
60WROw9n9lCwvsptThck55CBKe8dzyGzaP5TI9uXpyD/UGgLkQwu/iGkR9FInvfa
Uux3bflb4Fwwo4cKAOnHnNBGpQcxFg2b2zARDUHjjXrx/Ns4jgC6UR+1Dx5IsIuI
74dtZAtUmZv1F///fCqcI482IHyEhCwjLnPXH1Se3Y5NKxlFQ27TKBm7kUqLh/fq
ppimvJT6VJi8qWGJTlZqfXWWnjFRI6QBKZiEMUIMoeIjiJXw+kmMzgJO0XreZnsn
/nPdRiqI7TrFZgWmjJm8GzcuxfG7F50cLhhyeEhS/SJtYzPn7u9ychvzIgd8fDKQ
JhzvB3UheG7UsryHLCbaDgmkhEtDuriOzS5w1ltXI9c6VIs9vVrpaI/Hj30GEG3M
AProT/2YCTRd1cgha47d2YzmV3DaZQoeKvR5co722/tds2R6wD9TvdGdr3nTIGPH
IpJAWzbpKStva+3/4FUhmePf0FAqyk2NA5FUIAhgiWR0o8jT1Onv6cIgimFiXUCp
1L5CrM7S8R3Edlc8GupM3P41FtD/BuYkZOiLPJu0JJ9MP/rx46PTURBmbjm6rfiv
ctqkrXWzMqPGexKv65UVsnEWWTmhwPgv/KkUeXu6TqGVctdXRHeVkILf2zrdK3l3
66W9hcmNS99yHOUON3ccs74tcJIB6YuG/vFludgs8KTk7tA1TPgnh+2u9m4kyY90
D9dFoFSlR5z9goQtnLonwtBjCU0UQ/XPznjM0wq4dwBAvldZ/H92pZ3Sa0zVXZPG
/ggpxhe9aeKmnzrl6LYb6ATrjbd6tcO2KtrtXBGWtxjt39jZ7+TCQmxk1Gezu5yk
7Ro4geg0KX8H3q3U9s0PTwzakm3b60L39nRgoifaw4qvADUf3R0aKtiAkjG69sFY
f95B3WwSy9mfAdgPhYUz4kMxQKVFo4ITEf6wQnxuzEl9i1JeLLO4lTSWkHYYoqOD
lSZeOTV4BpLo2KVO1ggpH56xbHcRGFCEgM6BK/j4uY9vgSnthOCO0s3MJqHHoRtV
ArLSLfDdNh1ntr+gWmEzHY0/4G4UEd1S+dQOESg01TKh5McGJGvdwIOK5r+9KY4K
09QOuTgOh+3FhnEmFqy0IfvXgbEHaqMUgzWhRni5IKNHnD6wmsRILloFDavzRTFX
AjZREo5kVu2BwFAdrxOKt+jAEzm+HC/b1acKWvi/wBxMUlk0L9OQFp03wdFDf2J7
JgGJ+k6arroc2LhSiJvKfAftn79tNsNPJedMLkhxUmx8emmbxDdOiEy7rDUF93t7
Ld5m9msHwzAoS1uQ0fUvW4q6C8TGrK1c8dfyqKadE/JiS8SwgEsMRzE3PkAvriX6
+WCoa3Go80ikfj+0zy1nrhHzl3A3a4ekQV1bEtsm1/6fRPuS6dQFlle69ARZ8Aw5
5OnSYSPxAw4nvEiaM2MqMLhTanZ89Yu31p1nYNhwZvdLPidRFDf/5QqDvB/fVfRs
Nin8NvwSCLJgBSnFuZb0swSVe178ILvLIjbe2QfAkOv9Lt6WIti7ZE8bVIYgISyq
8SAhHprptt6ZglbqMhk+P/f34CuDnOdKv40WtxRPyW45wt0jHoetjs3VgX0Y/VR8
9dEPgJYRqZlb9N8qyPsS6XkixaT5xmCjNYrqaFbSDu6rh0HYR2VwjtnhOK5tPFq+
U6bA9dM/99pUkuMO6mNTcDYGTnvNP+Qd0rEOz/yjNGdUSqLZfQYgjQtnVBmdek57
bl1Asifw0SybaFQUrtYKRGuzvvsVhb48tLpuDqX+97RJuTWeLpgVGJ1pLSNTvr+r
EwQTM//pmgWOVIcCHW5nJRw5lKx6uadwvoxdGzZxsHK1Vb1bgvXLp9ANZ3emi/i+
9U4HA8U6D9knC/RbbtHs5/EwovPxdptZ+PpIAe5QfbYanxylLpj2F3CNiwUcBFWt
IBr66kDbm8GXCw+0H0YcJzv98jnN+lCCgCwv+rJMDsdI6U/HUGiERH1/i0eWRFXc
L3HBLQLpOuvg451nG+/Xf4EB2oEVzbAYdn12//NblR2i4WmDIh6g/5OxMYUh+1w5
0OLzkYD/mxg3ePi0DLL9f/PN1CK5hJfOhtUDzSXEYX3k5EOISJX0ZExfvrs3tZ6d
Gl5efWSP7pglGTuvWYVv/0D/fmzr6eWjx9cgNmEStYsS3jx4UQwQS/qCGNkhbj62
+IcP+GdZFTEWOTdxvsYSttGi5EzjKNf1A/zdJGbU3sS2fqy0gWukG8gc07aDu7kt
cipJXAlsJ7NwcaKL8BZAJpG71J8QN0ReHgPZKVMUF5KFXk4KrC/U8GR9OWN1aGUi
rnyWaxrpeqrI4A7KfwncFb/IRJ8BRwYcqzsUWuWSUaLlNRWuiAn7oRLarV7slNIJ
a7QHc/5RLderVtZUZTLuS2urUvEf8e9nvfFf9KgMFCAKdnqOoXsBjBdbEqQCenET
NejBeBIhu4LlJMZPfxRkSS0/UFSdyShiqbDIGeczbFMQ5P7Ebj8LM5STEue5M/3J
OQ4bLhZFCrD1YOvK9f0ov0FtUspd7X56aJ4NkDvODc5RxjdabXyXxpuCNoOzahF0
bis0O0SGKt7la2CV725gBOL0DO+TZvyps2XeKGMwmIvtJWdbG8XzR7GofKGYkgNK
4Tp3fv54UIot3qDL8Q5RwEnkEuX5GaiLp9++VmZLLWcEWDd6PcTK8Aafbz0uSzSX
gOnQrAP/MLv5kLg0Q1zuHp50/MgqCcaBVGPv+hEvJZ4hjXuYmotBU78/ThZnxusO
W5Lm3dMcsMiLRBrrEijo17eZ4Q6U+c8sACCrD/6Zu6bvSYidePW9hlfS8p8wtaGj
Wr92Ug3557gcyFR3MWitBDb3+G7JWQdIgru/2Tw1moRPtEqY4Idfofzd+wv7VZX8
KddcBSVtHYHVFuAKZrMXlGOh+bXB9aiw8BvJL30/ps7XXsNlC0yyTPXhE8r1ulu1
32LCV0aPjTtw0whIrDEDe1DXsICOYjH0m3A6VDkSo5U8W8LJU0q+r38dH2Td6k0q
G7kUtmgDb+sD9hBSXpkZ//2zELbP5JBzR9Pe3Q836jpJ4ZQ0IT2LVLFh0V7rvDPv
XR5CeYNxsA2dF5hpbKi9L0fw1cMTeG/n8AFAavSFST3UURwF/axddP6wp3wPAo+K
vPwoC/n0nN09G7FUM3+7ONz/TjhFIJPV9gq86DP7U+ro14OpVPxkrLDxn+o14zq4
gPirvchLM0YqMpG1j5fqdqjdXWkbbxdSiDKttmF9GdduhkHmdjpEGyQFvMLYJx+b
ntaqcnaRFm4Y/MIzFlUwsf1vOxApgSdLnB9ZkWzuz+JscMU8n627ADja6sgMXqNh
R8mmgCw3jZmBwwz4pR+R2hM3BsIfBtv32BGCU00mG2ooOCVKmEKZ9Ab6flpTWc30
XpKXa3cefr6i5ck0z73B99hxWBfIY0Qlk9AYFkydKqHQmsABZ2mP+pHzLT7vVx8w
hgRi11qQbm6Vn3RhnAGmxByTgnix48/RItzutBREzvN/9wIUBMC6eFJuIhcz41P9
QjSK5GZDkcJng84t7ZAa9hfBoQkVyll5iKDIKYCe5reqrEm8COGfJIhvIySGtek5
M3xrrrCgaGFEjt+VtZkehnXIVfPtAjqF5cqvZVkJG359G0QjY0SHRnWU31Vj6l3x
V63AkW5Fc3YuXCunadTKSLNwPLvlOu/gPA1mGXfjORAm+wBTa+M8WR5XopaQS+vH
LUhpNBySJjehfrMZd6hgdYPEghjbuY9DORqtejf3C2mjiLoa73w8ZZmpghrTGeQq
+sv8g8G6A5fAjylapjJNwsggk0IAhjHIwbLnHyqLFDUziub/RkUOyy2TqYNiT8w8
S/qfl24QCdGnvgf/1BsK5Zzg4VsqtTeM+g7Fbsv6G8kuTJ1Werp4w8lUQ1kg5xcE
4ClmBND9Ju7od68q2blwqAjz7gkS75lAMJdP6GjebNi3LzC7W3H/uq4w6veMXQjB
XXLijQ2tdZvP1Y1F2gTsAJHQ/8523gkHnKv1C3uM32dIFVDi48VdRZ56UZMYiFEH
UGpbwIv1shmfT01p4P5HsubqvZhc8znbdeqXhOriSGerysG8wLQO19hMV2yrjci3
2yG6Hdu6hXDaucr5jblRokLQJN/YwryYUVtxjEddPD2Vt/hnSTbV69jjZQV+y8Q4
n4KWCeVJBqXIxGxAqpObugli7HT9dQszc1eo9dhP8hT54lveo4A4JASS9iykZ2iD
1zYn0p1C/gFXYqoqr/V+HiNblx9u7oJT/tV7WA67P+lWU8VoFJrnrVwRfDl9jucX
N6Oeap9aS2kdOE0HcTNFaywJGqgTDmfFY1TTVfX5eVPrSFEK0BIjq38IwUqHgFM5
Y6iZhcaj33r5M+jUBmKxKI4lQ7QW4b9HID1wwy/wWNaGR85c3iYI7M3TEy7HD/Id
LSbk+M2nJngaG270CQAQKj9msOFNh2SIX6UiewrjLLq0GUarccO4qWdqBjONwMdl
+7HmD5g5rWgABYXi6vc63Ae/vW9RJVMSUdYlgjZxC0RIKZGTCAx6F3wnosxDbX2w
R7StpdVYwF5+0Hcj8ljHES37C0kje514VI0E37VNFCwGN1C+tTQqiweNQNqV3Ofi
tOewltE9jEBpQTthz2sE2VAzrT2GRfkVI7ay5eGSFCiZMCRLVji/nahdSQrw2p7T
xVexm4GrC2UnksxKmU7YWL1fri+NJhVFChy9QIgAI5qLGgV0OuUL8OBxz6fLY7j1
2Cqh55Hxo1aRqzI42cnSkz0EispqvnTlvs4UEfiHsgPwVzPLB2ZLasVrrKNmCP1l
6Wo1zzXFkphSENlKM6WPpColTeAM9DIE8KJ4WxN8D2nrm9Y6yitmrdOl5zaRhxjH
ny3wYF/uTaDQj8QUPyMr0mrMwxOSesdFez7t1eVIT9dawTeie2wrlyOTdjg8JpQV
UaaXq/241PGdWpqAmg8vQkUqizK5vCSFGiVyXkdvC603+fcY5vDVkx1u3ryk0gKc
nufhXTxuuS8XbK+KujePjomcNVekqb6g7kTQWlp4EDyQFvOnbskfa/2naf0bAH+s
y5K/rbY+gphHo0x8nD6bmT/14va1ci1hrQEtoLfvqsXz41pADmk7K06yekgeb9Yp
Lzsz7VtoUPUENLh7qAYVU2yIMhvlMArt6zpHR5Ay3EWLvXKgFmpdSKAK+c/Zdq6N
Tp61DXMNacCeTkdKTwwg8qJO+15eUCpdHV6/1CJv0MrBynC3+Vmu/9QHrTyc8WZt
hykEQdlIpyr0U8myRalNDJKH9w06f2jNkb2LkCDJEeOi2TA1s0A5GQgjF6fWwKLu
naFaYjzgZGjs2WkUXqQ4hp9u3S5uiSR+35FF068P25PRU/ffeAc9PU1NzKpXueIX
hCQ2Zqc3UFgnp5+UUUtrejGiRt8j3QBliVhYSeVjEQnqGO+xd4vJEnWuJQqpGwcT
pbsAU91adLW9j8B0zCDEtQBEdyo+cJejW8xFhabuwf3f95VX1XiOT/iKDtXUBItj
zv6qYOh5XCD0ib+lU+VqFd0xJkNSi29rAJd7IEMqSRMnM7Yz3PrGW5joWWz7QqtU
o7WGMIIR4olvuqDSzIhOgypqhhni0VB3mDQdUMZzp2QAgZlMj9yfZ79uprJmmG87
r2JbNDLnjaElYun08xIUE720OTbWoCE0Zek6+71NRobETJA4NJ6gZsvGhYo4FJ4Q
eh+D1RcHJpDBObM+JYaV1NPH/Zp6BtwleiP1apcJtGkmLjV5X9M35GmGw/N8R9RM
ZsLsd0z5eTapTd5NANMtpN8q1w9xcipV6Stj7zBxSgLS3uZyWw5sqmwyv2kqNFvj
Ap+uCxdZCvx3vxdGklqp7nihvPEVvZAsFZE2FM+0bszjQ/9yCwy/fKIQHr2MYaBm
xBdaeK2IELvhsMaozcEq3e61jo9bBi8uUtMehsig3O3SUYNtnR+vvEDtj3VJAuFE
3qn8CymyG1I4itIEQ0+HCKlNFpSDiqbTKbLdUSuyOr805o3q/FLDlF2eKZAp8PGA
Oijn+5Z5olu68NkE3fdF6O7FOXcGo9JwdS5QZORA5HqB1MGY2xN7MzWg70ItnfZw
+tehE32aes1iM6bzVfAc66VKhiPFleFPIr4ncu4V42uATGvm31Opk8dioTRwAPMZ
fl4ajTXj+tSXqCRrF+PW4ML2nRqh0IqVrUp0Yw5xC64qp5amdx7Kbr7u3UdK5yGc
omC818r7N5UEGEnjMVXxOuC3eVXAe6Fs826sifGOkuMjwkwjA9fkLT5IrD//kMMF
rsiq9aP0/Aw+4Dfz8Qz8NmGOMmgAfZ3NghtZNhFD7+//QNmEPjlU2TPPkUSSddli
BkyT2GM4u1vnnb8mr4PdwD8vhK8lbwfKAK22zpxtYAdESOA5zZQrAZXkozynJhhz
JEu4iFh2BolUJstELOGd1sGWF8YOj2Pv0WEmfsY80t1kxCehmhQYjeZKe5MMQQhp
Vi/u0/syhDJyzYWGtbmOoXsnIBwI/E3AfQboiMPEsUklfxzasmYZgC/Gon69Rgzf
uP++39Hp5bSoBYohfD8ceba73szsVPB7c2PM/UH+DPXw9Weje5tFUcmObkgvsgu7
5irzMde6iYtpKIFbqbDlYIU+7Ig432+Zv87b18VnobumeB7+zvAAOiQOP/fR4LZj
AEIYSbuVIj62nznGFCbfty/Ot7jf/AwYFdMjXfIK4qnUkB1P8yLDGqeS19To4Vqh
su/7T0oIBFp7v6hweO81C5krVz5p7enDHcGX7h7MftpRivdDH3QucqgzZlWC2ATA
6LD80aGwQl2e8L58MXxACRVrB1DxWKACN7eIS1p0dTGZ2DnSY0S8RhmA/Ir2rdDA
6NSfTWXVIr0vREVunQnXWxAjsuPv65prdyReGwAvbpzAfbQuvWNcxIJLp9NybOP7
S5kmzx581GCeTdXn3aVlQztYWuY21hSW1SWcG2dwQsHnTbZDXV5A/DH8lnNzn0P/
2SYVk6iedCC1OiGGtvoEpCNMxYqVOAoszpTq9vCBy+9e1wU/1cQVzk/5/VKgsqAM
UP8kfm4ijcd218Blx+KmsscWQlHCPfLiPFapPtUI/czCDZisejcjiKZ58UXxw4uy
aPe2BTF6qLhg9ndRYPoda1Ro7dQ+AU0Ht23VBmsyUo4/4jUd2BROZPuk19CsNXYY
zalEUE910Aj3gmMvRFntVkUGGMf7VRm5FpEy62/rYjXikO1rVlHvHMQipaQUx2Na
afRbvY8JQybyRVCmmTEDQ9nz/zcrNmgfqsaNTte6d/qY4iLL0xtXg7Vpus1SEJUP
CqLbZpuNlQf9KpiRgJ9B/dGyAkfmoDjWow2bdRCBRgCNi/0ooqFpNenSTYNCseFd
aF91j++UwpZ6vD4LutpjFyHsbd1aeFet+AEOHLSfZOWzppZ5ZGPAo1aIIqNUcAmc
/7yN7ufKbeSI2zB3aJHzqcJ5YtxuAMDDli/oOZFv38SU9Ljl683YKg5ftXJ9icL0
sZ9x1AlEVjPVArsI7kwIFYejJWqoPf32TneV986na4eXbrLsbh8EMCpe5x7wtAZn
AyOtzIgpLLCM6aJ0r3LvwD0IkP3Vrd6TIzG2Pv/+2QmZV2wErgRDE72iwERO2Ayk
RZwx0mfOJRRqDF5u89ocKreAcvNoWvj7BsQlw4Xj6FKHQzOuwUn/ObqnPdhaVMzh
fZyVeA16KGNIolOeXJ+CgMyfE2rTdWm6Ovzx6nc/2/A6PwT2Ju7P7pZUYMld2mJD
WZg4vS/5mI73VWyEH/aQsZBLdc7LcSmmBcjonxlEQvMHD/M8Rdvuwp7hoYlVmqdl
pNxpKSoT5tPgSD6CUZDnXyZMSONVa3U5aIsmY8Nw0Y1kybUumCqsLqrjhh6jhCA1
9KlWoePFeSNe3dyMH06PsN8oSnIMOwknIqF3qmv8WK70JGBj83c84djfIj5hPQya
OCYaCnCN/EZtsXMlD3Ct41WMJcq+YefDxNIHFcHWaPXkODS2QEUxYPudjWdIse45
S0E21JVez5qJk7C4ZQy+2XKOrc9BZae0BYRsaLZljxLXHb5LGtBkXLRo9wWVy90I
I6bclcQwspJ0RmujTGR4wv/0hX4I+tpyJSJaq7e6TvZYXVEJwNmJr87PpxsJ6e3V
0KThxivoxZlUsGFuvlyIYWYPpanlVX/UaymvZ14GCqfYhS2B2BFFTsKWFRF8GAj7
xpw0AmAM2oZQG7hDINkb96bSOeXw+TGmXJIP8NKROfMMWApPhgceTwXg1fJtOXXJ
ZBmtDvptAp8KZyddoQfV/Dw6Jxn3BZ/jpKEMvUXfid+4T7pegGrSS3NofBeEcgta
VN+OsKoIROCy/utAfMMwZiIzLv95DVXKohV68foQOeum8217sxIN6qpeFOcAWy7l
XznwkDCu9TkrqpkMA1C+4mFHgiQ5b5FigHJHrVpP1racwJxoszxqXYuAlg7ma+Ug
7w/0b/OVj+kJtQu0qVdLjbWLrsYUWbviz98iWvW7zKDLbhffIrmdI5w9/URnBlfE
nVwk6yuEOe0wZQEraLDF2ykBGKulNvUdwhteXSl6B8acUB4rHbmZUFudPwDxjN2/
m5uCvzyCoSefA+zt1R0tJKrvsqCr3Ol7V//BDe7YqOihBIY+BdgtcVOsWyKWOn3q
ErtzUBI/IfB7Zm8Mx+is4dh37VceB25UBoKoJsLvNtTGQLqLv6JEoPAo6v9yKNwY
0hUD68gEANf95Bp5ABAUBTWxFUd7s5ZaEdg4I2WdpjU14vRd1Hr5ogoz6ZEWZRAn
HKmpj8a2Aojm+MLlsRdlmiiS484ieUTNqsEARmtQansKNMEwp1k0f9WBi3PjC7/A
qzQQHlS3iaJXJ341cjFj16NlO1BQERzSG/7pGOCqfgjOvYJBLRLvypWL6D+eBTFT
0sFS2gr+gXcXSFydu7O00XWwqyOvnZlccStyVR88v8EsFBY0N/T18ofjf4WzlJRo
0NkmhribAGKgQV9/mk2OZTJPFrNUk6H1OEx4I5Ft7caNeVCwzqgDbXKaUP9QiO0t
5CqVassaSw0Dl0NwBS/InLK5UnYio/ESHVHVqAfx6l9KCq11KtOl/fW6mQZEd5Mu
gWmYagdN3b6WW/5uMfMpfvIBLdQaTmYK5GYMgvhHdRg8jZ/O4Qe6PR99X127SMK6
JlcXUxUKfrgrUOm0vvt5z5c0/RG7VK+J4lhIyGedjCYE9brc40If203FNQZ2hFFG
qxEkhi6Q3KPQWJIOdXnxSEu3ZGVB7G6+m0sNwy/JUq0BkSUZhNS8sXKTsi02G8Dv
JGcXUpY6QV5G9IXwVbVZoMRkDcibezR+Ojitl+mCi6+A12s2AvqAsStQ8o+SS7ki
ReDx372jJiPUU4sR2iPjpo7hHMcnBCXTGfzOHa7nyJZv5s5n8NF8OexCqCl1RZUw
VqamWszmuiQLUrLu4fIZiS8rxwPzqhhkApTfm1eSFVsO7ZZqBl2IS2eYHSWhzfQc
tBSQ1rMC3gHiAOK0kK2ueC0UwXdXnSpYjtuQK2dTCdW2lGqppyt0qFK13TM7ROEb
yKu+5vufB2BfjjjJ8cMsJpZCS+o5wPFf8xkhPSjrNqAEabrZJ0RZsyjSXQjgjjxJ
sP5Fj+1j6TysVkHf7XssW321Dc4tk4Eg7S9BGxqeCc3373kZUqKLMZgU/vR6Vj6T
FFFJsHQ+6ELv0SDNTreRlXwQOsJuUPZPUx9ZirF8PE0O1+VbUzmhOjGbKkktFzwd
rZc0vZwJhROfjZ3s8Ka6q8oFj8e9cYVbk4XLQFAitk9V1iNrkoxoFHedN8Md+Lmy
1v5tNXvEdlktrceCS/mvIZElFr+CWSZYf101iU4KoZvZQUw0RMn2SAlKhz8K6yFp
WPoJpCy5MvIo1UazAWVup0TxfRIUjJ+4Ps4A7rOepoBL7TkBnMps7FTTnvVynpdE
BRy4+taT6S2jDCuwAq49+YlvpPDrKJCOC2fmvqPvwpKbdCrd9mJHFsx/laLA2fcS
pPgoxIvI13MHiHQDoVhdNCuUkAMDMSrMW6+40+w7Vkg1sF9OgZFCXNP4+cC+foHs
OXeqKzHC3/r7o6vz17/Qb+wEwxgMxOe4sUi2tKR/BPsLgCOCSEAQM53xXI+tzwWW
mE+NMHh1CCkd4zG1vRFvuTGjvkwE1a2AaVJ2SQWb7/BDaEcwBsWDn0SVqPMKnQ9m
UjTwYeuQVIS38HxoHhzrI6Jy2+XbfSP2eiNB2AUMhMqbFw50IkcF6nx1NAhQNB2+
61HuFFV6MqVhETjDNn+92Q2DXYrA8FIW0CGqi/c0iIjqdqWqLTEpEekx87rRVVcb
UbdJ1PH39wSDpDddILn3PR/yV3qv/6wT/Xb8VEIJxw5GrqkjZCsKO2bpbeLCPRUT
oBlJc5JdEGZ7WxN7LVGrZPJnOMI+EuyxtNhGlrfR4N7fuwmrarmVU6SbozF92MCY
zkax8WL5xFozKTJLPdL+Uxd194hQIiTZwEHJmVvyE3P+0xlp8yDB7SXgWJ9yXtCV
JIQKZypOkl3ARwiq5APLrpU7s0Vjpijv+HzKirJkrhc64IB/t9HWh2o1jEucEC9A
YADIvNChACZvJ1eYA++AMeVELsGR5nLFgmh8mWoz/JFH8n5wX+hx8jtBBLyq+hJ0
GWrVEFE05yJ7eIO6w4mR+9E0WpTMrEl/qNICDhjjUXIlH4Ii8nqE5aTdKjoDZmvR
xip9q317wATdriccdbdkPQLL6hZv4C8tp8E4+y3d3nMqjawAJThumOqT4jxFq9XS
pp+vnwE63Ek4yMf15RVaA1ucRMrBS2xd6t1cp9cw+iM9FgvFnYA3JwQGNmMjqck5
DjSU1g0l5xjwKH8k3Zwy6RXv2M82Yvd0fMQjpWi4X2KUU3+45EjCaj4LS0hzoZcQ
kCkHFd00ak0zdm0TzxNbpJki3PIEo9QdaMKesTP2g8cSlgNXxEPkxywONGJ2Im1g
2cHEvPLBg4C3HmbdbGgMO5R0MSSzlabPU4cw8ulH3ndAo2xZE/N4I4TN2I0EptVT
WNVDSYx+eFwOM4Wu5hvasTTedTJdLEUbSWvBavHzSeQyX/3jKo6hELw+J0L+RqA7
heUhhy94XZ9OQOvcP5bSPMURTI2HCG2JXPiZGkVBDQTghNlc9s4dFlfa3SzSnFDS
oSmrpFnTTj9VJLoY2S0fEdr/6VjxjMiPvf7xx8NGMKxs/gMznW2IhhjHRRDQPva+
O8tJvqsMAC5e5ErnVrr2Qk4uhrWomnIU74M/YNzAAWzTMa3TeFSBDcNiT+VXhMFk
MzQvkXEMxrAyRbIeIkZV0qw+CkqxQ5iGcx7H4LbD87hGJq3SaCNhQRHPIy7qs4K8
musONHGXPxlWsPBcNZp/ag+aDeXfsNv0d7QYhskGiLAjOz+xl8raYjpoiFFR58Pd
9+OitLdJHB1JYVxhaI7k9hC64iYlAl0MIwPstanMhj15M/tPBlV3Qkt0Ie82n0+8
lMr60RoCc4aYN3unFmxCQnQf28kvvAkW4VuSzI174bKLUyQViET6IgvZAl+SaB9/
88uAM+gUVs5vedYhJlYDUFDicIaQB7lcSus3KesHeADceu7So6xnTBPM3wrLfWbB
R72XVEwHk6d+QVMsLXZXK2ubCiuFD7mqbQ9cBZgIhlnIPuIAq7V6SzT6sj+lXlBt
CO/8dRJbOWGgD33X6n5YbyWcPiw1z0icV1bMSmODLoFzgudxYVugY1VZrJQBNfK7
pVEeTNoxvwrZqmKvBrnYTjDzPcdvlivLliOvt+4F1J+MouJ+nHCl1iCchSiG7pRO
/CWGACkn5cm7iniEhYX8/i2W6sAnf7/ZSw6ov/xoKY9t3vopnZBqpBIilnTm77uB
zc8hqgKiXI8BeEgBFcNLy6Z45uJ21FUzsEV8QGIramPEOstSJjpdbtWDxqjK+nNJ
vnp1KCX2wcxMiYrEoQ6iRoDBvygKFN9WDbLFgtC2ieVAx7IosGqeNfA5OM96rcyF
0pGx5CVwkcVcszKB06MsNqnHeYvXryGEdAIMqKGxkSk4pTX3/q0tB+US6Zv5e1pp
ty5EM53W4q2lrDSz7AAt3LZ/PGyU/+fv4/8T+7mJ/JQhiK1pmwW0xs3Ddhk9DkQZ
HZ+vj+Jyt4PLF6Kid06szq7HHk/b/UCWGQioOFfgmwpN9gd8ku/0JbxdVQ/qyJqG
4guVB5+z7v+yRejgzNal0XnC7lHo326T4bRqjqA9gye4it5oT5W00Yp9WAWgGtY8
IoaeFx1JXl4W+1WHxvwiT184ayctmW10HFkqUA9C0d7rKPY+he1I6W7GJ7TDtKte
FCRynTNlIqjOH4BeYXtNH30JkGydLRaTABM71ZLtQNNwIG8QMtiY7/ic2WN5eEmo
Qz14dObrytFkYqhCQbBx3bPED7XF3XL4aLrcg1ETjClUS5hDgrLEFALg0n0BuSx6
MjvNQ/AjtarHOAax+12RJiCKEpO4XVNTsrTLZCkQbNTUSeWKog8U5XxkV8lvt6uY
qNw7Lz76L8VsrRBToQix2Na1cv9uR5f+zFZt71p6+Jms9jjAkCidboi8KcF4e5QT
3106oA4uCghuQ2CsK+EsEtgdWR7xnG1TQCjtMVRWARO6J7Dy5KBe1duzoVXELMoq
AcCbjC+Q6cO0B8mIQHUifWCtZJYEuNqmWuz3dP9f6pOJkh3aDOApCl2AJnzt/atB
WZDd8BBWrFfS3uFYkdYpWTD9TGl2tBA6aJ6RwhhZiMx7a6PD79j4wznQTgDDw1OS
SLPc9DZmDiWJo0dmjm7F+Lb5GOUjEI1eyZuPY66xu5pQRe+VKmJ3z22tCniQYF9h
Sq8g3JOgiQbWjfon5K7HOT6F82a90CJkVBcQedZ5m5Vhyl2irPHcrZosvDrkvB+F
Zs8WiiWWDiE57T3Cw6XX0J18JqiEncrUeLGnKRHJ7o0SzWMIP05mKvsR1ILlyZHg
AnA4guNa5rh1XgdcBK5JVz9IEyOwbsSBhTjxNRp1foXZMvmjkx/v6G5AEo/NgNFH
DF4o0cRwG9MbzZ6GnI6E2s+O9QnMbOFFr/1oUFGR+Fxz0p6C4jP9TCD36GMUeD8j
bBycbKZK8OTFVg+AAPw4I/Jan6h7RyBMGmBNaegVSr1SAEsoeudcN/J2c2LdT/5n
qJQeeVHHkyJ6RONi2xawibtHTNtjkbDJkhTYGy4ULWMY7BZG5qzV/aSxcZvLXuEq
Q9aDxsk5zHA172njflro2QPlUr6/R2rOAmcASob45KIcFPWN9/3LGllsj+3kcrpj
DQjWPPDqzsnpN5P0tp2PB6gnUmeAetgn3D2993uG46mLoTGycPeTCEAg5KDiyFgd
oAgRMw6lNfNrooGRAOFOEh5dychiRzCgdGLkY7UfaSVSVsgcOgtFfCGBAavZlXQn
edr906j05q7pv7bMJ6oGJuDF/wECUPKJKOkwymWRoO9I5Sq076J+UaqakqAtAX50
/epWXmjsztagjrKpn3TBkSFPlwokps5B9Fl7bV+borq1xkw69UV3ot0ds6+o+8vl
OMA6keakzTzQVLyTlk/fuHh0whIZB0mPsjTZQad3IyorNunms7xcAWtxD0EcMvg5
UUUNEek+rz9s8iH360yUtsKKZhX6qsj9l2DRbZDS7Jcy/5Gp3FvRBzTFzKxVu1nK
aeJ8Kf62E10Q8JLWYzIqNd045Yi6GEwjRXYhAHcGwrnKvTktQGVCu07qc98tqYeb
wRCF74zu2M/vxagT3uDZslXzBwE8DgItqNEe2btkAIMbPBl4nJEeveb90SHSlw6A
55Zpg9DnWFSZ1gZireKfbBzQLU8F3iWPYDS8xAeA1gWKnyBiwAonDyrHi1mufgp9
uK1UPqgrDZoVRfOr6rtFv7iuUJhSJ5vWbHv6a9ohMrYkBaDv0MQm3ugLL3+fhA+9
yym2pfz8HzC/ATq87ICPfjv9WAa4YE3UJQWV0zJQ2yP6HgKWY6Cx5G/2rG+Ee3kZ
8UQJ1moyEJo9xoYjGLkUQnirGPCXGiO2CWEU32toLHTArEYlrEnRrhl0+ylmNK9k
pyeaaMpjwZUx336uUM5SdPVIQaCV9/MEfvMQYUaP1XbVOO38kId0/ZYeS6kVmJRx
1pTiigZBjdaQn5zR5AejzQw+ZiQlKnIjmOTV+XDhr3FVXQmNtdMmPk8qdezFIcrI
hQW5err3fjtB/4erkHTut94at1w/YmB9s7URdc4XXVqsY+b55NO9kjQ12e2UEFip
JlakTzepJgRBOwB6D46y56s2tARTs8WZY3Fkz+E5U+gD1p2HN+I/KskpeRhKv23B
T/YRlgM5R8oroWGsQSepKhXdV51RXB9nm0wth0oPAwvlgM+Zvwt7sMxu274puGzI
fvlfwuPwqcAPhwZTthD5PBAkB5RyBX/gx5DWqNDANxofIU7Db18LfE9uL9KULyH6
KWl6qO8gvv1EGociCKaFJCgK1aaC+cLq3qTjJhuXTn75osYEJ/skwfusV2OFQ8o7
qnDOJw1UW0GlaFibJcLyxA8G4DddxHTFTt0SSiuCnaRk2xUdCDwc56JeK1q9p8zc
d6YJrGKgv9lcMLEGraQ7IH5Otof0vGrblOKCX0gqDDl65hXrjBF2aO+ksOYTFSTB
W1SRs5uYyhRqAVq29m12gK0BM1KRrK4rrlR/ewpdZLTe/lBZE5K8TvKsF9vnSNQ/
12huYI4x1KHHYIOWCgokcW3FRwAcsl1qTOnxqetRfi5TAljky+DHSWz31l5oT7+b
2xEfccEEDL5+AWB/yVerZcxFbxAxUWoeR+MCSycSd5eCJx8X57B4E5dPyBpPZxer
jemqV3+Y69RvJXylKXYEDfUYvE89kqq33jdpSOAL48eQFkmjOC6Is2Bibo4rzEe3
Trvsz8BAwzuL5BfOe6jr+rk976EeQ9ZIxXEigdMtWAV2tdDekKktGNx5l+9R0enN
yqwiIYqaX0lq0Cgkb/cPL1jqw1w4SjK0sMx5ApQcSrk+4eflyuXTadQf4t6Murv0
+o6oNK6XCqya0jz6HXmjXgoIDABpy3Eh7GMplg07QkUD/lc3Pq4c+D2+r7aiGgj2
7ut9mB8Hyr/dpJyV6cAf5DfBRAboyPvU40Hv9ASLCQsxuC5NarX+AtdkFnze5/Fr
yossMplmNMrUJOzXTYrIDLG0I7GV88TOArKaleKm5xMwwNaagl/UqX0d6cmapYwG
OQLGtlM2dt/yg+LTsKur8sbJOz6vTgVq7tkhEDqlB1jet+TtZHulRX2HaQbto/9K
QisVm6x/3oa2XodvJ6yMG4XzF2OMpV8DbeqTdsQLUuPSuoK9avQv6bYzw7TtbwGk
2d4Mk3Yiymz7Ko7w6plR/K/R/RSjPpGfpKUflWq0mhTlEDfDPVFdjMB4QKCdCVqH
/J/8A+JCBsnoDgUm5i7XRNqAokdGSXJynUChHjW/qc8WnTQOQJ6hb4UAmvlRCfV/
rvSW+/nWEKo3K7l21NsjM+5bOIhQNGQanaBEmd3nnXPrIfBY9JSNVIgpR6VBz5U2
qaPrJaccgp8NqVSPNtwqWEBsDoV3f+MtBXUXYjCKr/ZDU6k2v/+LYMbOIxTSultt
fTrBejZK0E2GO+Bkqrv1fFagAp6cAIATEd3kmmB0nVOkR0lEB2NwQ8Qk2gC7KdVs
pJAsAB2l7IY6x4DhGSA7865t/NPh8Zboexf/jL0WVt9FyDmiGZc9GzPfrsoASK3F
K799xE8jHGMsIXC5DehzwZ7royAxU1JmBB/+7lhZfxggowciJApWeiJCG0OUppO/
+5+GLaeLvBK2gOfu5qRdIyToE1zJZ/jCmzEbLrpNQcuJk9YYJ7AX/P7IpTCteg0I
2G48kRwmz4HUwUeKal1jWgQrIjqfVVffu79y5VZEU/AyFqNeXhBC4bE6AhOebAl/
omOjfuXYsuo2NYAsxOMrIGp+NbmKh1UncaOe4FYCl37jAOdmRG5ZA4KQZ8mh2oW4
4I0/F6aPgmhjmzonhTZ57hflsnKbgHOLKcPucl+KhdsukC3eOpshj2Am42N19ovm
PquDVedc5BEV/qmtLrnv8qdo8mis6/sRcsK5wRuc66VabcP2VzXFrdcSo6utF6EW
tR78todd8MfQxVthdIdYXkjI1dA43tI7anMBflWWpGsG3NZVQSfgqX4IpTUT+Aex
ZUCt/CZwqhqUws8o1EaHQsn46OOtVThfwdHXwXgXhJdqB0Y2RkCmTvEenU7FyQ4R
hrB+u6n1alcfaMJ6C+eAtFtJ3a9osx99E5Egmda76j7lDcTMIQLx9T7H/mAlJJO4
cku6h3rpilzd8CzXIEmMCKIVe/apO4a+RZSJTJp9e9yZHfa5oSdBzBbJt5cYsWE0
8umhCVlKgy/pivkwbtkozfCl5tRHVUY0Wl+iH3N4oh/yae3Xf7zHrKFJKx6OJm2g
7AvvJvUjCVxNHWvUcrQClJNuI4FLOSvg8x/BDRQfbcIMz+rilME4xI/yFyBanc3u
2HMHkY6V+g+4VTpg0Nyj9hzmlXpX7FGvRVA53CJbZ86PFgQZU1Cis7hWwcOzuOfy
0wDhm4Iv8R/Ma1Ejfwp9c71WOxgPqa7S4XjFj7MynJchqGTQzaAlrZRCrX5Lkzq4
e4/V28pJqBPWQ6xUQgGJQvaaOl82k93Ae6FBjWhrgdJ277kos6wRM4nqUQ7T6CXy
nxiYUiUVHL2HtVkZIf3A+B24FGvC9q1BS05KbYWi+i2GHL8nVAxGNCbkQzEhHet6
GZoYjR1TPq58x34jvd7gjulDL3uNOQ1bgrnlFvCpUpVcPEMfwIs8QLN/Kd53nJ3X
1k0Z868buf2ET7ZXn3vuJ6QvkQ5ocoS6WdHlom8wMMJrorDN+s4tE3aH24/v/Ak/
6+RL7s+CCeMswBQIHsWV8ewmATpzH1gAECDVQII3+Woy4kB/hVKCr/sGgWL06bha
3OMZJp/e2/YD7liEGs+2mu5MmjuvD/RP4LuWkpPpCJjQSPmU71EQCv2gk81x0JcS
HA8Sg/EHsSQS4GfRTTSTjOwyFZp3iSFVxihcX71BuZGpIzdo9vcLFy1OUaSSq++9
kRWro1RILr725AJfvkDhFAMSHgCLw4QY0n5I8RkaVYKERRLDE6n+Wm3YaYlrCxfL
LyX+JlwUeD2scP7lOa4nAkCcpkSnP20ezrJW1hFqe6xwmh3K3scBjB4eB3mZ8Nru
yU72wJEqt9qXM0gfgE2SDxEPOX98v8h6BIWZRMRqtoZeUp8meCIXICcpMgeUUQcR
zRxRIdomD2qOXj8bCuHNGrDjurBAi1n3cHHBi1kCdxdjm7CzXJndj7xTrUWRYJzC
9SZAE1xRPqqzv6pJur7L4qqALttCoieXB9oyUv8FS22cjkVySH9clJOCbccX7dBH
`pragma protect end_protected
