// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H)#G?Z6X%@&I9K;E[V0B\M.!RF[3QCT?A_%I?*?/U[@FZ]ZOKHTVD0   
H<^1"'?W)"%M13]W2U$3#03'_OT#.@<QDQM!8D1>#>6ORUW,&EP KKP  
H!&#;AW'XW8)@X,A<Q0K!>F#_BI%W\W:)7H,IM]>I-\',PSI5'>4]?   
H'.W Z-*Y.#83X]_5]86 "?]T:6FF&<A[#?UVQ#>&4+$92C/!%EO?]P  
H7VC^V7A)H<M-.P_X@+9J2S;DH\UE:/SR*[H"81!Q#:1VA:'(#-*J60  
`pragma protect encoding=(enctype="uuencode",bytes=19536       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@HI"0B.U:]<90F^#/2U^_C6_FB;IC+D+!"B@2$Y,1+"( 
@1%W_ CB<L2^GOLN/*U8RQ155BVYHK7U^J,U*[#@10;< 
@H90$1T 7 ;RU,FG$Y!H\Q-Y.73R86-$NV(L?3GS98U0 
@8:$+28Q/GGN%,NBM/LIKZZT5/WU1U80F)R,21V?#KH\ 
@M%#>#LT3V?U]"/(9]4VY@),LP00DLF,U1SSN6QAW4>@ 
@/%"NT5AY"!V$Y H0-!\F>"*GG4D*@>00H2,Y*<"LH[4 
@R\P#%$#-VP2<X]C1E&L$7B?Y:AXW@7T+YU)!C%!4N7@ 
@FE@=(\C0BJ$=0S">K\:4'(D4\;A?>[P%#&0;"7:!L4T 
@I">/0**KSEZ?,C;,MG%\J#Q> $'S=J@SIV) _A =*P8 
@O@],)<T*WN4WFG.8-EQA#-X4C%JK9>>X<89D_+/J$<  
@+>ZAW8(@W/S&<WYJ]("J!X^@#OFIF>PCJ_!P"#P5T[8 
@47F68MQ]QFFN!P>0ET*SE.ZS'5O87E(JXZ"R$2N#MND 
@Y 88,'(),%%9Y5V2OK?WM<H]).PF73F@")\F0(W@U>< 
@'#DGZ\"4ZD/"446,BGD:$QC)K'X9*->:B57^B $$CXP 
@EX#IL#'4<:=BK3M:=P^1&/)*B%&4XZ<I)%1V3A:Z"_( 
@.1R2, 29_E<P4*#4!PG9G&L!Y=DBNM,:DX@L=?:V#<< 
@0="?(^]QO7[9:Y5_E9=?L^(:U8%?ADJCBD$?2Y>E63L 
@M!-7:6&U-3Q2<RLZSORQ6R8'&_Y<T,XHK]/LD1SK%M@ 
@S6/@[O,A&E"$*@.M^E0<R[NNJ\C5&1$[W,"!ZUH2KQ, 
@G2S_-M)29.:G*O4J/SM_ZU/Q@W,^W?9KC4;O9#Q_7/8 
@T3S"QD]3,A9UU#36_7"C+LY [@(S6OJ.P+ 'OJ.-/;L 
@IUG$G66V_O-$0=H!\]B"80YGYKLU]P4A>+3P%KS+0&4 
@([D;,PL'*;-+I$FLE]4BR"TEI@I0P'\OBJ1B6AEDRL, 
@DE]AKPZ,WTO9V5$CC@%=O.+A@%%;!5!)1O[8#@XD#^P 
@& N>P4[\<?XJ"8X"B I* ?=F7GC6:&^%9T<;FT=TF0H 
@20U^OC<GRM :%S;]!8-)BL*A!B1E@"%,0>QV5-'TKZT 
@,:C82U!6?+>KY+6$V 6@Y.>2K?H^'C5LQD"N!VT-"2@ 
@(A8RO+R.+>JW0]5<4&Y6&S?L$@% ML%9)=8;]Q!J!D$ 
@E5'\&$56O\T?AW.G,[Z9\I$9093:C6_\@/._@Q;:<C4 
@7W@2T@$LK '+*1N".L!*^U$HS'T >*FX;"Z)/G3!/'H 
@<>ICOU+( PCEQ\>L;0!$7]+J9Z7RK:ME8:^ PYZ8L0  
@)H/6M/U)OR-=G-.W]443P"GU&-<)^F\]2AE,=\SO;\@ 
@ZZXC_']V3^I"%$=X'Z*$N6U$MSQUPLR@ %>5%NZ R<@ 
@ V?H(/*)XF&57'9TB9ON2N)C]!?59 OP4+F ZI*4P9  
@.SL,5^TY46P?_TQ&;]6:7D+EQ$9L;(L'6)*((8X8*.L 
@(]XOP$U_OY9*_O)(3(,5MKH2$?PFO\6W'0=)U+P#A5< 
@1^*PTR.]RF<.]8>^L<F'H4+WD#0UH9 /Y]W.Y=>CK2P 
@YABB ?2V/FZ>CF%C BIS=?D(U%QY%M[1AB+=Z6%H_H, 
@7N7UEV.*#W)-I&$E013C%Y[M:/_ED>\@' =,UA'HP?D 
@*I!1.31R1X*[#;[S2,';Y'$U DE@;X(0P[,S6-^SN00 
@\:?F(!2I*9I;AD[((9Q?#H,^R&_5OB5>$[J+OURXZX\ 
@1Z5-32+O0,K,^7 9YC8!0E C^.YM=;<"3 U LFT1XJ@ 
@ 1Q5ET*_KT4UHKK(W*>V]U ZL)J]W;]VKW.*BN,F(7, 
@9RBXO!FWZCV-$7,2A:SZ@4^>)P\,M+J&LP6N=;65?/D 
@"\^1,QY,Z@Q2',X&^$X!X4^FT_>0,,.6.WT@4B@?H.4 
@CL$:0J8V"?@2D 4=2W5;&IDZ!;IKGJ[@X#6E:HF8&V0 
@.^;X2-LY^L&XS1(!A1*F%D%THT(ZS>RL#H\$5?)=;?  
@A "3($]IJ#E67J[[$ZQJ?G8O_Z^V/FO(G:;LZJ9\UET 
@@HD@;K&^N"A2!/-M?#@>^9)R!FUE8K+;)P)F "#W+Z, 
@78ZZR\WJ?4@*J9M*\CVAZ$'FU5J8/++A\8KIEOI]DQ4 
@.?V;OS5)%M23[4^45?RCH1>X5L,'3V&4VJ@L-XP.MP$ 
@Z/92,CS="I):=!MUK]:7RE<1DS^<&=RBL8$(K=UJ\JD 
@Y<+Z#PX?':$%IJX]=K"3F_CM:3W0TFPC)6T]2YW<?58 
@'\Q+T/NC&_\$B^H"-*]2=!W2Q+CL%,6TNT_?C6[DM@< 
@$*TY"WD!UL!WZSSCOKMZ#?3%J2J+!S2]K8WXT;RQ.#T 
@I>1]U8]S;Q'[1SGZ:7?0/BO_U@L&+ E]7L*[ZWH!XVX 
@QQ0/>Z'M@R+TM<7OA9V::2->^5+F:U32]X=C0STX1M< 
@^4!]H7LX1=;#&8$5Y KW.80?M9.+ZD1QXVE_FND9D"D 
@-4"E&L^=2H=4U]CZ3+"IQ4AEU:NNZW;JG3 F@"O'>T8 
@,)\)8P>.$,SRZZ1G)6++T<737\!YD2,NKITZ-;"\H2@ 
@S=Z ;,Q+][P5(7NSG97E<V]>+>1(:(+L9/^)/+?7J+< 
@UZ$=YG20B:J(ZQPZ0=-YB$%2+N_//]"ATWI1!2LFM:H 
@$_<GR+)"E"^1>9E%2D-=/ ;'SR60+]6H.7C^M*!3W9  
@,M-Z6H:$;I@J"QC@#!=.!Z&C!:[R+Z.<*J\\B9!T7=  
@HCV!K;PQ6MRNRJ%0J^W4OD5C7F'LVW_9R_M@"R49_EL 
@UQJO6P3?1*T;GQ4?I^:%8%%+WRU")LX'D_A\VF?3PU< 
@;T<&CI@?.%>F)>D63<0"WZ%.X/!USQ?JSO+)SEDD[10 
@;)-*^9$E8=9"X9F20#7N[(>]=<UD =!D1)^+PKC1/?8 
@8KKC=@"@<:</)]0UBK9$R)4-=FUPW[V ?Z+1W&/P>I( 
@H^@^HDCZBWZ(Y6VG (6CXW36H#!J F>M25?0( (G>Q8 
@OD$AMUJ#KWLN"O62ZXLR@ E,7 "F.=@/K[@31 V2['H 
@'<WW/M'7"66TM52;3B**LN>%6BIFUZ9 TQ443&V>GY( 
@^GN/#(N-!Q=\^B<:LWUR#33-$U&"MMAM<),<:'/P@FP 
@7*('MP^?PQTR!SP@WGR6NX81(M"*:<L#86?1S8^1W<0 
@C><+SW.*3QY=BTWH_3(!8QMKFL2>;IACEV=JV[0V]VX 
@U_<2@\.6Y"CS$Z3RA#8P;/"92'C\++RB+<[!Q(-&>R( 
@" :![SUAE:4S'"\R,^M883P\W2D$N=0KV\Z5[V=*B!, 
@2I3Z,T=9.3^*D=:Z#)\AS^X:0%L*U>0+U$!BH^4MP>@ 
@MDQT G>)F]! .U/I3SG[J2M;<S9B+YAPA6KQ7L!EWL0 
@W' C #41@75L.-Y"SLC)Y9?=<+6G1 >$,59T<4R\#]\ 
@_Q:XJ)XE,4,Z^02L7TU#&!VTDZQF*GR$,,T;=3U455  
@"E$BR_$+H>A$"K0@>CV335V_OY7<P+J6ANQ@;.O%$KX 
@IY4;U*_(&F9*%I" 4]0ZNQ(B4&;.HQKN/1 C0_R*$?4 
@:3N@PHP!KY2^"<B[[ID9?>=YV L%A[K\!V(>R3,6[SH 
@_@U<A*33I@^C'4-L_6=]@"$XB<2 +JGZL"G!D>:79=L 
@GD,ZAR;SGR6KF*V8G9[4=FWH@>#SH:.P;=CO FB(_#@ 
@7(,I7^&?Y;3AF@?ORXD>Q.3*AQ4A7GJ,]M?L4>3Y9-( 
@G*?T5$+4KF_!!+S:8-;3^'6?]&=0&3Q[S92,X1\/,2@ 
@9I!XDDZ*.,^.(L?3MEC8>T.Z27/NMHWH-E'Y/@:H7DX 
@_CJ*!5=H3=?U7Y 4NI*%BP,!-25BJ4CDWMAQH!)A=HT 
@Z^_)$:/PP%+A*)U@J\5*/$(P0DH F!/(^0$YW-62$OX 
@S\]33=E"A.#KY 'L[Z5_F+*J%:@O>W\@H?!IF8+)^7\ 
@.+59N0Z<F.-F40"Q)=G!RVR)S-25#!['=^QJ#%(N9 8 
@[2KM?7%OTFQM_QG?,HB.$?1C,HXZ-=S/8+S$MJKS"P( 
@>5>_4O1*XS9-Y[OP:S??[&A&GR,X3<'H.-%H[37IK H 
@:T8!L[[P[%QTXIH6DFD6KX5)6 3JVBN:U/(YFG?3'_4 
@JG:L;FD%M@RI/1QA?VU8SFP@$V7W37SY,F/#[.X-/B8 
@ @*9Z>H_)!_27'3<9*MHU>Q72VA(;=U-K8HP>U-:%LP 
@=OZ%1W*R]#4;#JFV:8N6&@*ZTB53'>59240\:__E)$4 
@<C?.Q=E3IW(*YH2#MMU8@[4MR*02OD4R]^O2QI2PG?H 
@0 ?3""XVJ=DL&D#;1?Q]0%O07EH L&D>Y3P"Y!-4&54 
@;_T '/>]]0]_@-; DHN+QO K#D9DH/(=@:V@<LAB,UX 
@F6%BPB41H6*WDLQ:CD(MK4!DB1, 8@]YG!QKA?_J4GP 
@N//ENW?I>K[R8JMGAD9@->6P@^1L!&5$JTX7[:,3$]$ 
@9LV9"S9"S I:#XT3G\]RBL^]:_;7/;%N?2":>P;&^]\ 
@;+Z*%K'-!G"]B#4<C%[@_K %)DQLW<"J(MX**J*69BT 
@<AVF+LRJ[@A&(/TN,E-?9/Y!"2QN<<N-;=0 3BEZ_4D 
@1O9MFFJ),MNCD0N L@ ;M!<L^T')\1L"$QEIM'81)L< 
@GR5@SB-6<.0+V2GGCI!] B%=(% 173I@L!IV>>=!)L< 
@.'Z)7\&,S6NVL6!T'B=!)T;B3P0E39Q4:HTE-6_S;Y4 
@)XIH7]4N8V_DKW)8 VEFV6)+-,.WLM@^]C?!NAVZO7T 
@=U@+@TF[_P0#^NA4LD&3E^EH9+97:K<30*AQ>W]A#7@ 
@;F7AP^"3%ITHQOA.DN=(SX:!X\YL!&36U"UCS;G:+,L 
@]B .LQ'QL5IB=WO18K8]YP,EA^2CKU$E=[X:2SB45P$ 
@)U&9 R6XVET[M'[$& Z>(_*&1NM@B=-&A9Z,D-'Q5?T 
@@@ZY%613$A"9.G6L"UT)@YXUK\*!M"3E01><\6&%KUD 
@M_R17;FT5&\>RD354C)7-7.22$ Y ;2C*CP$')E?E38 
@)%7@QW5$Q43R?>X'*^/_Q:HPD-<LKEXS^"[0LSOJS)$ 
@_$J>$#C+H)BFLUTTP#"+2,MR<"P%>"^2Z5S/?5HN7B@ 
@E=4S"8?\F*\5269SC>L5Q!H0+8DFKY4[&<WF5.VO=7D 
@'WW>CO3KM-NGR>"+\81XC5DT<*A-Q^)B:X;XU0E8+O  
@WX9-K3"EI'6A_OX@/UI92D"+OE[?ZDT[D\=$,;R4Q9L 
@SXA'3)L<V3R,CQ#3SC2VGY?$0GNPT#?IGXRK\O]\)M0 
@7N,X'-)_D1G?Y8SM@YP'M,HH$2<TD4OR8HA'!;AX5V0 
@L^=%"'RR\W@<.*9K0"(5]*/G2N!6U,:EB5E,;A"TA@P 
@ZG1_>;(H$?XPWRC:>>:7O0D7"2,\>$PD/.NO\="@*0P 
@XE.C5_SAH7->-7Q.]E+X]9I:ZRR4V,($-ZH3E,G6@)0 
@@U&".)M!B8'EM.Q9;S/J7Q=KF)_S?>8VGNUK54PSAQ< 
@+0;W7%6L%)(E-OD!P::,C7SV"R(NF='$R-;'FTB"<.L 
@,UN1DI6ABW_U])>T5+!\:]GM:$M2D]D !$D#!;DP@O$ 
@.K=&\/B$K=_;M1WB+85.(,Q"_J@-1A$8* .*VN8:K:L 
@+?R/7$DP >U0#"4B):R:<:T&1 J]AD"]?L[EK1*X+M@ 
@O5;SS&-A['=LF %(ZT8X>L!WJB2PT3@<CT+C@^LZ,Y8 
@AUCK:X( WJVIFXZEVJEE?SR]/B77B[,I==9;GF0()U, 
@D+(LR>1BUS+JQK@L=F+8\H)BQS<R[S]:DM1EZ%Y^&M< 
@8944/ V%2&+1*+/,[^]&?2K3GLM-WF0;M)XQX6H"=<< 
@TO]>Y8AV+IC#H\Y-3:^9BOQ"'F.JD3+_7YG+< 8FXA0 
@5Z>HK:\;^>M=U[?]6L7;^FCZ;].0W$ P,%]T@H1J/=, 
@28$T>JG\)9F.1L>/VYD79:50G0'"L00E3 VA)C42@4< 
@GA$'[$M@>!LXIU:G<!S5(^-:0SD$'%?9X^O^G7.,8(< 
@4G@WIWP#?:F&X1Z94_:D#TL6T!VICC@7#Z+X!QQHO.D 
@?)(L_8\?[[C[/1H0/"[J_&DP)+91AJ_]0AFMSWI0(CP 
@P(5!MCP5D79LYLT791;X1"'[E#!=($?:)O=^KC+(1VT 
@F4Q@U+%RAZ5#JQE496(G=/>[2N?4E7+MF9GCL]:VW)D 
@H7[E=F=^$!*QMV-;9N^=I/H.]QX^3(XSS=,'2L34T+  
@MA:KG'IE6KY3F.V!CNE:; /R! L?D*:OQ/(>^/_>*0H 
@G#_A0L82ZP0ZP>7,.8;-CD&U ; ,*B:0B+J#,LG7>#P 
@H9W%AV]>I?:K!MC872!&):DU?Y!%_"5Y@0%-QW^J"YL 
@TSS0EXF2WG1M;RX LFC$ 6;6 UX)KJ?.,KF;H5V"E_X 
@ L:[#UFLST]8-!0=ZC>P[-_L(JC0D+W8-1R\<&VO=\8 
@4%!I,RWE_(:KNS"Q]2^TP!+V?$O67Z\R1%]W\S%C[VX 
@: 7\3G":7/6<LHU+XZ ^ >G?9#/97[/OS@ Y$=D,=@L 
@([HQ(6XRY 0!" VKGP2ZY/C92^%R[^X^X[NB]34'2<@ 
@4*RM'7D**@NYJ;VX7W[K8>VFR.6<Z2SCQUI?#BYTLH\ 
@;@P9&/"EG0EM]"EP.#Y=:^&<?$=?&W9Z= #;N 184XH 
@]FM1M&E30TT/DBPFRNM8C:V^^-J=W!$1#PY?=9:GI3D 
@T6C-/.O)NWB#_[&7B2D)+#R(M0RV5]9S.199FX+\ Z0 
@ES7#YS,[<;17:X/21#>A:&X]Y_;#WKB"'6T^S@YJ /L 
@]NM=4,7KBZ4?%QJH.$;D@,%?L(C&K6QW+\X;QOZ:JYX 
@Z\<B>UA<-@&^?_IDUN?W7"&@680:V]'(N\?TE0& ]M0 
@"G1*]-ZN$CV!YB?+TG(%X)TPKM2#9V%#\(\G:3YL R@ 
@^P>^6<C=X<]2V06=N (>-<<-.JY%\"HZ&J]L@1J=)F< 
@0ZR@)'IY0:LH)]PZAXW?  ->3F0\S<(T-Y(H[Y\[S+  
@,8& UIIR-D]?%]E&@_B30.;$\T;KZ3>F%7 =6IU%(-@ 
@DNAC7%@-=)2_X7P9YV0TTXE@&,:2F'MW: !AX@B9?)< 
@LAXZWIJC * 0K$9DM(4'MY7PS8MC4\, HC[LC/:KT\@ 
@YICZPDWRB=/AJ\H0WIC-+8AB)P*M\FM D)T5?'03TR$ 
@.03E9@,QZ-!ZA 2%-I&K(0Q+-T.#BRV[)M8TVJ2?#]4 
@,=+G$H#>C6R0B@ZD\T4NUC&6[V'S* Q=%5];3CT\0+8 
@*=1 6[)QN2\?TZU.7"1609]-"4CW)<A>="Q<M7^9V<< 
@8(2!B(TFE8:SIENGSN/66HY7  :?LD _75AO,161:<$ 
@*V9UL8Z+TD77++!73I,O2)T,/$8NM[ ':F,+VS$U_@8 
@S8\1#V9X63W-P8#T69-]&Y65&. OPHN?L6<*AMYRF%P 
@.*N32_M,4&/U\%)/$GYK3[ZV.'DPK&&+%4P91FT @@$ 
@?--:Z[)3(\L/9P1O?0IGV*N2#3M[^>FDR:-R#03(SA, 
@MZ->'/UL0-V_DI"DW&&X;L4*29I^&I\6*"T7"(G]7K< 
@N%E8*D]N#7M<+7\+Z=WVACJ";3)R"G"]MY^SN?."I&  
@IFUU(8V"I=E(S"I(S+7=HN?#!=2/J$3"ET3HIX >M-( 
@CZ4C[-BU1UOO=2T+X_K"W898$NJ.^U@*5SVCVZI1Z90 
@S*-Y<\M0V0B"KGT;!=^F>JA(BRMDM(?G#N<P];*""/, 
@V;?\[9%GMBN.45-&.IRNX./H%7G4,$:_[_5M-E-.P9X 
@0WT[] M7Q5FXCA?05Y37/XS>)AH)9/*AI!VP;8!%]CH 
@GDSVC@UGHD%0LLZUO(PI#ETG;__&*4;?MU!%98R=NJT 
@52P3W[GG7=&ZYOQ"#J;1&22PH4[/DAPJNJ*%#!BW8], 
@UFBIF<YZ'(/<M_UV__FH\M8M]1WN,, W%?]T6+6-8W, 
@X=X'6D4PJ,$C/V&-O#Q(H1][,R>=LZ%2CP4&-95C9 , 
@R^X._(S?_QV-,@5*R:JE)RNF\Y(/&)DV":U:"9]NQW  
@R%,.&JF,MXXP&T6.)K*&!1'K_]HC$J=J*'C M^;+WTT 
@1MPALAYTF"V0HGOI<;"'^J4;K_KG6)<8@#-YEN&DT@< 
@/*C(E?=4*3:@%(]$CJ4([VTC[QAC983E#Z)+,C-NYF4 
@O8 !.PKX^7;[=[_U;L!50>3N-1:]MRS%$ND2ZYN"32H 
@3U: UK[E'8E*(24 HS'S/E>I,!>D/&1C0+Y%R\O\;Y@ 
@@?<Z7R0Y0\J4DEH+PZ.[S$OX+\B-I[STET.7@=J-A=D 
@D)X+R+8Q2(MRT $]\&S%S^%=:!1Z;;B\KZ]'/DM?2A4 
@9!_.33>K>%%?-3<P#^W)T^<$.\#V$L6[=,\Q>-R^#0( 
@<CN97@)" ^N(@?OB2 ?.>AD>'ICG,]/C!Y7TMW-P3Y8 
@G$'UY:C\:[!76J!JAHHXBK6%3X^R0AF42R,]^"$8A^L 
@GI5]D#NE%%"-4;3#>#'7D\ZR]3WYD>DL\^:;3$$\F"4 
@J>/\W=#)98@E>@!(Q/8 N=SD=?!Y<C! \EDSX'\7;I< 
@*E/IY\.=2$Q9>3PM1]Z1E"-DO]4'=J_&I=MH3.3GO,P 
@KINZ(GB^TK,&$A0FR[V3Q@'0RP+]I]@1Q<T\?IQ.%VD 
@'[Y?%&,*[\<H!A"2 #&;-*<"Y-*^GA-RV-NMQM+L)/  
@984S/U["E5D^9P;0'LT<$5X&<[FJ?$BRM4CX^YDT'X4 
@PM@,]#M*[<6&'8J,,(#,L^.ISCDR07FPL??S3>X,!V< 
@JG7AK30OG*SFO+FX]GS#,620?(H*07,HY5RM/%XL5.T 
@1W0H#<J>;YTQZT?9I@HDSB+HFAZ>G/E;(TAE0J&**%( 
@<]XD6_I[D08J6*M(I !AH7F8X]0@C4"$6XA%-7EM5JX 
@S'Z@2(U6D%#*EGQ@P1]<'"24TG-86E(%_BSTKFS(P5( 
@NN5C1 5R106E!S3;IC:;F,X%#UTLS?JH<,*0>I7;W54 
@'O>U:W#1.MYES<+(#=V"6O/@"8S U(O3/2>PWEP&VM< 
@8@;4RE,GT9U3V&#*_L.'<<5F?$D#R?38&FIY=U@I<YT 
@06^%,7"_)?#0)!X?%/R?J!FZ2.]F:X/TN@%@EL:0(S\ 
@/GU-J!=-O"NYWYI:8V3W4["!;#J'B%82<O%[7\J_-3, 
@<BCSP.+LNOALK$2&(>&Y^M2F3D,+3GVAFLOAA_E9"', 
@]1NGB;PR!\JP+IEC@R*9O)3AR?'&)UM]G6HFC,IN*.\ 
@!-JQ*82>?<DS@ZV--F9YM_J3-6..EOP%WSNJ[K-'X4X 
@22: E\_9"C$E)SD1@P6S)?N3=Z:UU-@_*,K =:*'=D< 
@Q\H#[<_?Q;H4:"UF.\2,+AJ-EIV+#L@PI==UK,G5G20 
@L+$V-LQ\5Q]EK@JO54K9)[.=E=D[Y8A:,*.FJ[U YA4 
@Z]"4VQP=HY8[61)*5H+J(R_,GL^_H?7.6E[/Z0@P^TD 
@>NG Z2<.;;ZV+7B;!-%N^^[C"RVIQ3;92L=U47/"'?< 
@8ZFOM9^!07"@KG1RBFKHR?\>= J>-1O(=?^\"ID\6[X 
@OWK\+'[OEYL0C+3'9[4UL&#;'&UP B[:KPRW@_F=HEX 
@FZ 8*##XB_)P( 8&D@$?<5?7ZLXU&W%6_C'@Y#\DO70 
@;38(MO,+2:./+S+)IUOU-K45<S;&_O7-'(BI1MGC2.  
@E'LY@AU ZU(0-"F(I2H 4R-@=.TV;+U]X/;Z7 W3$>L 
@(G"060%$LRLBZIOQG_PQ2\]5+0FIS(F6!&4TG93@%"  
@QQ!EBM0XX8"MMJ65Z.CNC@E >(C3+2^K8=B75TM1XG8 
@>EF9#)3M 5 N C#807XE7\Y VSHJNN2\QR1W$N$VEU, 
@CA+FWF&B#R+3DRIP4#*8P.S#/-\]S+F/SPNQVI<HNQ, 
@TH(EZ<R*9(;!#+7A+&#UO"+#4%3J_(:$>%Z&]+GY7O0 
@3F<%5@IC2ZJH5]$I&L/33=90 [B:&:97.&P,BPP8T0( 
@Q2(LO[EJ&S<K^,&DX6,CI$HQA#.&T+:BD/B)#:8P*"\ 
@-].O%W0&&.-^L3H234Q,PYC^*M,5\I!)'T\L56;&.,$ 
@^"ZXS>RC>B^'_@DAM0"W,YVF=44PFU$Q/0+2:!G8Q%@ 
@)K/_;"'M,\OEQY=OH,VD6)=5/J)G$[64_:_F7F5\O\0 
@S[FA<-DV-8PVHP$XHTOR?L6BU=69IU@ET3(CCHKIT@H 
@.MB7/9S"L?=E#Y1DNAE;WPYHU8Q+RYG[M"I^4,4I/'P 
@*,6[7"=5@>(JKEO6T:2V5X3K4<M";K\$KY68IP<./(T 
@/6)%&))\;(HFSU6^&AXS1<:7S=0<Y>ZXT,OAXF3G6[8 
@.=<9Q0X<C5Z#X+ K*/:H9N$1*:3(><JJ!XR+?G&L9C8 
@..?AH)>I$H (C>K3T.KJH-XXYPC>.].E15F&?Q!"'^( 
@[9D?PG5R!4V_W+N-KA&@3.![;3Y&F#TH>33=Z1/IP"T 
@*SG=V^TH>\RB*]%ZA&( =*M+O6!X08Z3O+!C:^JT\.H 
@"D F7C22)RE6^AR7H(J^^*X$9J+:EM0O)->""!=H%IL 
@Z?WXP0?&,Y#YFCV5,1<.><@K[O$C068-ANBVJXV6_"$ 
@G\*"0T+W.885"YED1TTYS<" ,7P,/=GC-GXP>C_-<#< 
@LB(U=5>S0W QE?O'<G]>B!:#M&GBFZ]BW[V#-^=-$ZD 
@M1YLL3>K0Z4XF7:BF)*\.1/^E'!<\ YQJ7$HZI))G=P 
@Y &985"+&V&)?%X+JB_OWT6P/V/: #RD2QODL\Z'=U< 
@F)]V]K=,,B)T0;TWDLFK*]7XZN81J%2J1V6#+\Y!@0  
@^=;?J?'PH(%)M<O]L:A!^VH0'\44BP/SM?#KBJ[YL]T 
@)><CGJ5]-Z.J^9>5BPO2CH%M%MB._SDM#G?;@"472GD 
@%WL'E!4@A6GZ4,UI5#,$WWN1)@01Z<8 /&Q&C@W-]GD 
@@;IBN?8-Q2N!SVQ+<+2YG3UPPYR+PX;4,A[8F(YJB+L 
@*+H+B*(Y=T'JA)18SA-XMV&/-M19P8G91G_2^@;8LOH 
@R$^5N=44G,JT3]+Z5XUN9CVB)ZYQY@\,P3LN@:1&'D( 
@^V=E84J?WF5)WA4ND@W*Q*@2G-J?3U'MZ9J"'I-C[N@ 
@K$6TBP[!Q/9[;AM<>S-M@UWM>XN6<F';G@S!5%=X=P< 
@'<T535\>Y[JW# 2GJ/YEVL[:"244SCF__2RN#*"FI!\ 
@+CE$:TZH,#WB38VOMB&HP:PHC **:5UYRE.=\:<CF?  
@0:J<"K_S-1N_7(PJYLGP-L 1>]PS+7J>=(K$.K+GKI, 
@U8D,#<13+)#X]RU_Z,F V?:6UKL!9H,4DW1P8[ZW9TL 
@^O6IMLPRQ0$#CF;;5)&ZMW"NZKVM4@2B:>/2N4'SPW, 
@@ 5XSY4IBDD30\7VHUP&,#<#_#H0O=^B Y*B?,,\8/( 
@+DZU&FTB$.:VY&47 %!CJ6$3=TQ-'0T3ZBC?@^^M8LX 
@TO"05Y!5?H70FUYD3MKT1Y>=V>L0/&YH)DME6WG[D:X 
@P>0COG+O6A(@CW91P\_:7K>:#HLFV\623C5^_'J.QIL 
@QV-&1@CR+7W]COH&)(=M)QD8B,:*]A-GH!'L3U:/TTP 
@/&BPOPCX5X;%BR*O CBQ![BU2_9]N4FK$ D2\8^PW>  
@G#@K'?>[LY;;P<VS$#ZTK@$JN:,#JY]G-\SNDI9+'5< 
@!I%IN$HC@Q?M7>7L%Y6/%T^3QI1(9IP<NOAAS<9"2B( 
@FEO) 1#(9.SXE*NTB&*T>)3VS/E/L5_9R*EVSH2V>&@ 
@H+6$9J[45ZJ2AEQ$_BSRRVC=(^_II#:CIHP-MG='2Z, 
@S]H '>";'[RR&27&64.]MC":Z@VR"#;5B&#C2)!2V+( 
@YY&+9;ZI)OHS;$_/(:<MU/IO),?HT75=^E+$66@[]'D 
@LFSXY-'@O_M#13UUGH)YY"^IEX '-RAL=G4]/A[N)VX 
@)XA2)//#L12E>^A]D!9:WN.1J3ZPDE[-GV_V?]K012P 
@X19OK69VJ+L*^C<:L0YN=<FSMXBE:;X)^$U'ZF34@?, 
@9"L6,/?7-]/)I[:62 !J>:FPI(1T7E$G6A_\H*=,090 
@<=W8X<R"&ZQE!Y"7]XCZ_-E"Q)T&/JY2A-,B-*ZF[P  
@%ZDJ@,L^"LJDE@1%<.V!BRUK/9F$&PPB"M!,A6T']^< 
@28+NJ;37+BWT!J"GI:(.6SF=$QE N\^@;A9?\-M+OFL 
@TVAQ!S# W*Q'J1-DF+L$2MLU,#[/%YCIE4%Y<BZ3::T 
@N/7 -&2Q.2/].G\?D4KQA!Z&I3T?-2\_$G*$ZK)!&$T 
@3& /Q=8O,((]'@]\R_7B#%!0^B2?VZ9FN%/"S5>9DPP 
@6N!@%K>O5P<WG#2,,4]>.AW;RP!!/]G35:67K9+(U.( 
@<0@J#:?H>K_\]5&ND[:@C&I;(!J/^N\ZRD9BF9!T_&T 
@-.&EIU.<36!#BI[<>"I5YLH12KZ1:SXHX+=^R^:*&?\ 
@[+6S;[?F7$UWNM-_1EI!WK0>"Q8;=/>(XKY8O ]0D*H 
@7-_]9+SE[13C@U18 $.KTY5/2J#WNJ.D3W72]]^#C'0 
@NT@&6?W.KBZ1%F5&\%#\L6A\Q)K;J1UJ5TR2$87\%%0 
@Q[$G&81B)K&&OOIHTJ[Z<UR'6+PZT+ 7RX)-MV6T8(@ 
@E EDV6 !2JV;8/GD>%;K\V 4.ZOG%G+'F@(2B_ZP9O4 
@$.DW^!D4E"I4 ^BT*E9'$H_#DP8*H8'04D,2ODQ>12T 
@T362F> BJ&Y$D#3CC.L-0M)O%:51AT3?LCENMBCQ+-\ 
@%ILQKTN%KIVF%9$:VN1!ON5'J WA2 \5K*%0)S96)4@ 
@5#+[S ($;0!8!AFY*K;.SS@U!RHVI+*K(#6DQ-+A]UL 
@@&B S"SY*[:(NV<MGFX,&\"%=Z_%$7.<=&!M@LB=LP4 
@'5)J3S4)0(NN*)Y/ FE]D3-KF\P:FR?MAN%1YL=7RZ4 
@2@E%ENP:#T!>D!GXUZ/UK+<,S'$(9)EORWL@\]W#%&( 
@YO$6M59\EK!;P7J\L;M;(/= MQJ!?RPY)S4_4SF[<[D 
@? F,&FCS5?@2]M9W)Z_][H(<557,U35&!//T]BY%[C4 
@8)]@AO%+;72RM\WW7RIA21L<NC58>+A,0?9BC&U^ &@ 
@ 1[MRQ#F\8J^D3](\A>:N](&IHX+Q%IVU21<WG8$?&0 
@&:C%"WYE1QA!WN(]O6Z#";+^B//U?)YZ@FI*/_DT OL 
@\*51"F49Q-)>H/4D5J HS&?9^+ \GW0X(A7% K1./KD 
@QYXQJ$0!PHU;H-@=J/N/GI#1O@'D@R_:L[R2RR.@40X 
@@ %W5KNP(H5HR;5WND;R/ Y >?U=IZ)*+R:+XY<:Q-$ 
@*V-;F,JV8&5SN;/S.8-A4"DVSX! /D-8:F*FG< D.!@ 
@=4H%H!70(JU53=B55O&'RJLY&H14@(K4/K4G&/J/F\  
@&= U8>A:8Y52Q,QLTO'X^&!(X\"'2V'V-*0EKU.1.OP 
@ICWWYO_H%.34G1^)6,=!\S#F. Z5QU$6'WCQ;F&@?:L 
@U(69%MYTUV9>OHE2F>'OK=,HF(RH_,?[SC8FBIUOJ!< 
@;P3>3ZY[8T7M#.[94)<MWYE_#D\PN/_@;T*#JV=@%,0 
@EO:O,W]%7//2;.^;U*VL".(B\Y+&;7!CWY]4H<RKKQD 
@[KDE)O#=<1[L7L5U 0(.(BICH]V]7$PO+S\7L'D;_,( 
@>X]5*K[)ZV_2?_F^SD08:!&;1BE(-C;@)JX<G&%1<%  
@9"H$A;,@()&1A.;Z.3/4/<UA83\O1P5?R4 D393=@]< 
@*&;"C>Z(39R\';YQ?6P%)?^M(_()5Q00KL) SC;\&$, 
@3S02]@P# >33 M9QK=F8=;\1R1S,(?K&[8RU?NG';#, 
@;Q;>_."2WU3>3Z?SCJ&;4\Q!Q>.X$DXD4O%_W/_^6>H 
@A%E#XH3_(4)9_&[;;FX4.F&$<7/%=SJSTN^,Z]2I#WT 
@L^*U9B-GDM& Q5M[,H*UGKY;[+%%(O9*1EP,SPFIN-D 
@P2-DU@GDDGAZQ76\KO>F\&V5[AT=P)([(FBJV$TYL.< 
@ HUADFV0)((U37=R>&KST-I19V<_.[!'7V&#X2\4RW  
@ZXX[PCRA8-X.@ITPWPKC5TS3=08)1=C[5K3-F 1>-,T 
@>FU!M*XXD%(3EJ4#5$]3W4$;$/$L[P6SD"'07=B+SF\ 
@ZPH:L](GKK)A ;L?5J*LHLB!M;-/N:^2;.3NM@=!?'< 
@X8-W%<D@N\!L%H#^ECL8/8OJ6B'4KYRJ[0?XD])8<@8 
@6'4?6,0]->C!M H[MK97$VNU6B4U?BVX H B_HEK-Q0 
@:/:SH\5!ZG4K#'QF*/BL_<%<;97$OJV/.;)&ZZ'O%2\ 
@C*S-M7I6@<!=\.H)1,U?"^D\1=RX\9QT"&B/-SLO&K( 
@_[6J9X/AS=@J=T7A6L\>U &%87#G-I^RM05DD_WZ<_4 
@BAV=AX#D<<]2E ;RJY0I6,5?I,0%E-&<8<==\@=T(:, 
@H+M^ZPY$=SU_6]?("9)2_:F(8: OUYHETJX7/(_=NL, 
@B6*#.+<V!UXB\ 1$"5(3%MJR_8T9C9$R[%/JHOXJYKX 
@:A9%ZZ@#-H-=5R[);P8;FVH+^$<R8I!MJ#\K\Z,RTE( 
@4GP7J^NP%+8/3YQIUT Y\?P^\@T??0]"Q5L(%;SH<Q8 
@1NU7Z[VC:ZJ76]FZ#P]KZH%=(G\>Y9_MW!\?PEN!&VP 
@!A?7_"5-O(G3=D,JT+U()P)&!H6-WJE6+NA27-\4FBP 
@=XBF];<A0B(JVX;: Y2C5+OB^*?=RLS#3"AVU/HSNWL 
@.W7-S9,!K_$H2+)*A:/1J>K>;N*[EPWSV-+)>D*Z:E$ 
@GJAN8#%NZJKZ@X5*BUJU9*\\62<\@X$GPCP^-0V(D3@ 
@B5LA/.';=@Q':#7F(\T]_O$&H?"_+/CV<YO-O1+_(/P 
@5CND ON@MD&@Z?G+BA (1M--\,8>;,"\J@72F4J-7*< 
@G"B98-CT^".YOK[+-GB?NMH[Z.(0UQ"#$<NO1DD4^@  
@6]M-E;B+OK5VP=MQV #S')O45U[61H-"Z%](ZQ%\=58 
@IVZ8WNX58I++0XB:2P.E_*I43IUH&MK,H;GK0YM#X!$ 
@1M:U.  21UP!3Z4_X4<.#XP?JU(N_;&:A(.-/0#2E?X 
@UN\+$?1L.-I^DY(!NRJG4\$]O( (U+*24 3TU[1B=2D 
@3'K )S-J*$QEBNINRB[@>E;6X;5I5-$"81"+S.!#$%T 
@?!ON8:WBD,%NQ6+8 79N0&11X9DDW*T]\W;J4>1V$[@ 
@05IG2@EMY9]-8JLV"&D'A=I("MI\F<EZ4WF5SQ@7+B( 
@X+'"O.+/L7JK">&RWW]H.ZEA3K(,L;E#$DT8=/&VFP8 
@!3G=X@'B&Q]Q(1IN#EZ!.XUKB#H3 R*06*-9#;&*W'@ 
@@?R"H[#MWAI.-R5R&@O@ZD?@(A-F,$(?SP[#P2\@#X\ 
@[Z^"1^Z?/$NZ73?ZTL_KV" ^74531)UQ[D>6EV@-=?$ 
@>;KUPB?P;BK 07TN8Y.L*TC5,]1]KF[UT@!;B/N/G#0 
@P;<G&;]/$?(F,1_X($,>Q3T =*#I!(!PA)JE/D-NE , 
@VKU(K&L:F>Y>W:5ON8ENR^SU0I<[N93=X:<_-\*4.T  
@+H0!7_2B)S2?^)FQYX&61!<2";JQKB1GS0*:#6%-RY  
@QAI3CS&\Y-HJ<&2Q7/D>==?7YHRSO\ <+'M^]:%]S)T 
@_'59/RW9@.V6%@K<)O HH>DWO9%?[/##PQTEQH4\R$4 
@5O CG)Q;MU75/%%'BB^DKVO'L-C\VE5K25N%+HQ?Q.( 
@UJ9&Z2NS.>!<#_FD%)=.BO]U(G1MA$MOU5H*+E\XM%$ 
@DZHT?5JRLC^V2%'/>QA;7V5ENST2VFL@@)!$)49>8<D 
@!8MP^Y>ZS5'/PDHQW^AEF]DYMC:#\I01.3<7_F_'6U< 
@]HP5+/[]2[W.,E;Z/";$CK0P=+$T'W]5CJLW(*;M?H4 
@V;XYSTRM*?VY"*>ZXF['[)<E5UOK3PI.9GL--,;G%3X 
@,9I[/O+(CY_Q#6I4)IT1)U-O-J--ZHL58TKTT@%>G(D 
@GJ9?>(<6T>12FT:_"1.B)H@D&%@[$ [<D."$MH9XA!0 
@EO-9.MX90OVB2R/9[O[@-K?/&,<;GU\>XQH@;U$\Q<T 
@]MDN,8MB#Q!B%99YZV\6:'?09]#"6>\!K.F3O+IQ3FD 
@Y;+M9JMVLFY-7F7E49:,TRZ6<N1IL$^VX3IVBQ'D"Y0 
@'548-%44\P3L/8KJ[9F10QDT.F DR2O0T:Y,Z1D3RY  
@'*%,X-&JYXZY2=A$)#)SBES3&]Y2B_6P<^<M&3J"+38 
@+*C7+3^P$'#"6#<36FDLO\7B*'O)H9+8G*IKI9>T$3$ 
@?/?D*80\TS#0UYQ&%2/</\ZZ*JQ$UQ(KJ.+FCI#?1OT 
@H(4;54!4@OKW)';4:8"4%US:'J!:"AH<R\\0R=G0H40 
@7LOYL>6=^^-=B($5Q>\1-L&MSVMPSO4:6%1A^+Y"$GH 
@#[,K7XW&6P,5W^L/\!*17/C9GEWZ4O2+*B;^-)1 ]2L 
@K8V$;U31H7]\ ^P=<=HJ]<3A='OP9XJ17;9ME7(+SPL 
@:9T,=M%_%VL'&YW'$'I"SVYHSR5?Z%SK)"'Q]?2/UA\ 
@IYG;E97%HO->Y"XZ):ZA#%H#[JO0!$5LJ<J68C;I? @ 
@(;,"(O8?"I&\-J3S-O@=[9X+]5*QIT_6>OOZ$9%[D:( 
@HJB-X5]QB1=FIT@K/W[8&;GMM5W-[?1 ><EGZC*5(&4 
@N3(1+R:2/8:J#M::+E-=0G;'@* EF'0HEZ=7=+))8.P 
@FRI;P_$8Y]1TYS;(>G>3E!S6+RIGI3 ,D-(0U0?(YT4 
@1OF711\K]2);,6+,EYEZ+S>.=M?7R 6L#X07&F-&/-( 
@+[FP^F](EH'BD;]]&\0C(+JYZ]J!%#(.2)B3V&\#@+P 
@\M*\!.XE0(=7'=LPIXQ.CACFC+UJ02PO< "\:9BH6ID 
@DZ?&Y_QBKW*0ABG4>?/R,[EN;!98F9$="A(<N;PV3LT 
@X@?;GSCXX>]>Z&Q&9?- ?._6"K11S,LB8^D%: I?J/, 
@@D63U!@FT->B O@YSUIJ[QZD?<G:W//?J(4('?,",68 
@:"5Y.8: ,W/6$!YLYLG>"O!5.<"8\@^89#&*U ]B3*$ 
@D #6J)M6CLQ1*'4#:J.(-WT,_ ;B[C;/"G5^A.@OBV0 
@F$-MFZJ?D2%1A4_BU0CNE8K8&8B4"X@L(-..P/$X7)< 
@92 CE?VK*^#Y!BGP"[(1S!Q8TXTX&*;83.KRL/@Z]%( 
@XQMNBN49<[*'B7+N/+B=.WL#T.NC5V6P,8SN!FQGD]4 
@'1MFI#DU660%4G434%3ZBUU4<H@:QWJ=[HOZHO8<ZSX 
@K;_/5)DLTB3K<((5!N#[TF*BL94T^I9(S_4]L&FS=>X 
@>%Y!,0CTA4=UQ@<ZZH,PS+LSN^A +@50M[>G*^['#+8 
@/-3,$464IVOV+2!)N&G%! ;*R^8T('IV#7EAN5F\1VH 
@-^LM3U60/Y1K+Y4E%ZB@Z?CA[M\V_SD";X7&&QK!"B< 
@C7!^BR)42C=D8!.7G9H@)GO)<_82=%7O=^>U)#K@8(H 
@T[U) ]0KR-Z/N$ZS=UOOS]=P2<$D^B%-R0-5\-*S0@\ 
@H'E1 $"WC:+;AH 9+DI))^?PCR^4&WGX^L]#)-\9A@, 
@;89EA8DI0M Y[0N5@M(#I*A_1H!#19$8]INX%U"D_*< 
@& W\.!OIAA*__0%[X7#8G31]#,J+?FY^_R/W>B5K,U( 
@9"!R#6_%21QNJN I*!P81Z.\0OIT(V$<+FG ]Q\$NW8 
@!\Y-FH9W&@1M @U<ZLU(C@N+U18*CG-_JF!Y@;.]&J8 
@%=UMX93>E>BK\==SM[&$&26*E(;^4P6A9BI@D\,)7.0 
@GIHM=1=G".P0XZZ2F*$/VEN1 _"]Y"?0&4Z,#:5>ES  
@^ -']*ZXIYN_'\_RX0I%S1.3HYGYBKQ6+(OHI.D/I,4 
@HC-[&6(IG#'Q4Z>[><7:Z2T?4R;(YL!P\!>C#\$B$^\ 
@Y92LX272:*(ZO/P#W^8"^TU=B//=P[WPF.$KYQP#O8L 
@GUV% MDHE-1#<W#L IKA5['"P.*@A/(RN-W11]S4O_  
@')D!KW@UZ%)YGAB@&;VD_RDU\)/R@WZJH?#,9)]%58  
@M7"6\EAR@;R2XH! BA]!BS  ?6BE(\NJ*L*C3MO(XQT 
@O@>-=P$6F6L-TNM,$6IR1\%F@7D<>/R/*202<M?!"4\ 
@)!];V4IDK"9 6,>EEB48@PK[1CD*VP6P@^Z4ZN%M5]8 
@AT>?M(6O+:K?]G.@##R/O<Z$0%' VY"I["SLP?>J;,H 
@X&[89'J[3]FA<[X:O$+) '8Z @WA+S<H @<3:.G]/6P 
@<WX((45(AL">MZ5-/;PMAZ!I?B6* .^WN>X.F&4M5Z( 
@ .IO%8[3)<HYYFKK;;M07AKTV/B"[DK>'5MOR&0R PP 
@7*(IG0;8A"?>37;$9"^[[N$GA5#%<N9)W.>>I$%3W-L 
@9YA])IZ%.FC9"65E/3E^[/K6P,BM^692Z#,[<!:ORHT 
@N\>2QL6ZIZ9YHA8?T(]Q1;H253FP!<ZE!?/PU#X-U[( 
@4H\$U-W6J5L*X+P?27M60,3^# 4 YAH:X+RIQHYY#Q( 
@X3W1H&8W:3;"HPMKHZ(^FVKEM$MAI [E!3?+<@)8(4< 
@PBQ1[7_?GC6F@' 8'9X'F7,WDF432Z%A 1;Y-,E1?I( 
@T?5L'LU?<K]\!T@0::L?4_JB=V]#PZ01!J\R/L1K:O@ 
@-A&K$*?5@M\V'RP_/N\Y\%-VH"$9A9X_\];34#_+6Z( 
@A)M)U6T6L7N/@E\<$&["(][B:OSAIE&2=WAC98,7!9L 
@^3<TPM@,B!9=$-*.^25W=V[/ZZF7HH8CLTXKR#2W]P8 
@SC68G!0V:O00"+2CH!(P>VS]O6L'1*+=G[99V@E*=R$ 
@= ?6K&):'&!6R<,&EG!-+2<-L"!]FLQ0:7C(G9SP U0 
@*<PY9X->/V)XX0%E\#;V.HV\Z@^%6H2Y7M*]<M=B;\\ 
@#T5(^G6<7^AS6-F4[AWJGT7I=\-/Z)M209AX 7?X>[H 
@J4">IFO7J^ 5$(O*GZ>?0BDURV<O:,1'$/92P$8E9<( 
@0TN%<AJ.-N+U5TA\D'EEFP970X#3N D&940_G7K5;I, 
@SZZFMD6*[JM"T6N5&-ZQ#&%-210>[S$"D8LUS*F^0-D 
@P?&E)P_>M#JN2TU\GQ31##)+?BU:2^W<*L3;A9.W3R0 
@Y#,WAO"I$/K%"%&A_YB.:I*!@M)8K9Y'I$@3(0L?0^T 
@@0D1\O"GN0E3,>QMEQOQ4G7(X'&F['481!.:RVN"\48 
@-!T-JG^X"URX'1MFRH[C&U>Q>&L]L]T5I^9$U>Q#7T, 
@1^(68#/!"BG_;D49_%3]ZZSK9*51*H"!KN3*17%@DA\ 
@>7V&CVOAU'MZ"HVC"NDMVN9(]T!M%E7O@[[G6AQQ 0T 
@AK "+%3YLF\FQ8":6F%Y(OE:ZH14CY5BG)E9D2V>;U$ 
@Z8R6Q0T$ 9<NV#]Y,]'.W0(3.\\&#:6\]WV:)W#V]XP 
@#_Q6_,JY_:D-@*H>8:!@+L2G\\KIF-RW  #]O3S4RN0 
@,GF@YEE=M4,5X(Y(!QI3.X=/&!5G<.,7EV5S0V95II0 
@'Z/Q0@>FMUJ WP$R[Z;0>UYOFO1>V:;!:M[;Z':KDHP 
@OM\RWSS;=>=9H4$;\4CZ/5/H!*.MSE!&E_(IJ7H_J?\ 
@M[O1GGL/_LC!8H![N#$>4O#N*^[S0C1+8ZL7?VQA(+< 
@FQ RWU1C@&$2JL5*AQDPIE!,H(+1/8_3+O73P6U*@YH 
@3R;L.E2EB'6:I0,FI.[IY=+ ;%"7=,'O((]4\JO4)&D 
@+R(J7@O:%L(1)=H<4&1@-'85'W"VRML+X"<CWA\#;-T 
@+N64+P?>OS\NRN%:C-Q96L"_GY8LUV2O"4DMSZJ!BM< 
@"")EY<[@XHAFVL)]#YG73_[WR 5XPV<N5E?6%8+6&F< 
@JPTL*<7HF$V7YXGM3OWC:LK<4VMM."_[UXIGN.K;OJ0 
@<HYH7+FO=8^[UT$O)#\#;.2_G!X2_-?L%EVI &NN-RP 
@7,6!=F*6ZYMTN%/RUSU=WLME9\T\C60A^Z9 OET^4.@ 
@0)0Q M)R# WYSR6(FL)$^<PT8R2 E')/K"8,[P_J"AH 
@5L2]8UZAY5Z_<T?[H/9M@#7ZW<U@7?MT0@D9,+C8C(H 
@Q F' 1G]-\II*^=3E[3%XH_A2[J.;/*/E"VTZF0%0BD 
@":S/-N(X(KI>CUP.9"*CPKL4?(OS@L*?)Q<:"D8C&:0 
@\DUWB@UJ!UAY= MX*!/K=8HL$U5M^:,%=PB*!<;W$\X 
@LH.]WF<NSA$$=K__*:UU,_ZVM&RA%A79Q.R>%'BQ45P 
@85L,27.%-Z(EL.%]Y.Y!I2%;R(PZ/KS'NK='N7  ]G$ 
@F9'D!8V_,G# LKR5^Q30RNBOW^I-B$NA!+U;6T8@D#L 
@*K%TKG?7KS-5O&9=R,&FX,?]F%\+[BV1H#'H"M^?/J4 
@)+U&2$[!"%-E"9$W125^0HOOEGPP)-:D'.HN=TBS65  
@>-K+:M')G#"]?>;06-^9-315H6%S]"M15R'[$I/,L2\ 
@CQW"?_BC:S&/E+1YJ1X][Y0E4:ST!V-QO0U]7-!$)ZP 
@#.)Y,8%UK-@@%CY%BN5GZ#ERI\:9.T+HJ80=^-<P^/X 
@_4ME&LRY/-T'QS,>^BSX</MY6_A(O8 WIEHAN&\ IJ$ 
@&5O U( RO0-K^B"FR0C\I)JGUT,K82&.I,G=2NDPL-( 
@AOB2OJ>9V"'=>E40G$B6^M )!<<'I+/T'04I8^SHV1H 
@7X@Q6OI*#HJUB7S#>&<6,#JPBS/0LHMT]C,N3R_DN'L 
@=$-LIY')@@8UQ2(16;IGNZAL+"OD,(Z!))=B'YY&@DX 
@A/5T5)9&5@[K)4/8[W#%7SL7\^)9D4"UK51D/F[J(%< 
@$+RN#0@*)6&,QHLA,00)BWI=?@G9H'1VT1OR/$86M.( 
@PH)!1^&WV[4;TB0.5$&3YNT/_HW_BL3H?\U5S:,%1T$ 
@+L8E%CT*]5;6\%Y )AE4@G <*![G2S0*P_U$ R]D=JX 
@1\6Y"!RJ?KA+^2CZ!LO>H1S66:95M-;U8PW_FMMN#2< 
@(Z%X.U^9LZK6T&;$?+ZI<;>EX\NMX6IP6"QAKT8:_N, 
@1&U_M#PP4IG_#22Y1_-]:5T!D")4&IS!T1T8G"0=RG, 
@[2U$$-MM_6D64V($N5M>)'/1NMT=:7KMH"5U (CB.R, 
@Z1\/R;9[X*=:@6B&@OYE$=*1\Y2@K=6>:>>;5$7G_M\ 
@57N@)VYHRBU>!X\<I,&C-F!; JVQ16X4+[$E-Z*- FP 
@08T[&5,LWRN 7*1+?JSRF;8R/]IQ.^?20<%DNI\0LL( 
@_Z*2Z-.N1>X2F(AC"RLT.AKUOA_,0B22\Q<P+M]0.OL 
@T5A/29KN@1R0?9_%Z-GV]3L?=6Y1%XIB3-1R OF/N]D 
@/)O>MX]I1)/:S*G<W88Z6;H# DS-$VZ?&;N7Z"::@!X 
@#$O;T*2)UW]O2H>E%#"ES*A#(<N_CPZ*<\D$2?]*+ @ 
@FM8F\77UO_K8&PWE7O7P+T*C)+71IWK2@M@:GM#Z*S, 
@VRP[(9 O*^ECKT_B6^SJO[TD\/M-I@R(Q[C[MMK1"M  
@3LOP S <G^+)S\*#LQM$Y)U3^I@V$2*65-K\'VKY; X 
@#51.S<$!_J!IK,BE96]"A\\UXV+JET4.BSJQ!2<9[ZP 
@FQ.1AM/ [K&HP>N397>"KI=UG:R/Q"]D>T3@&CH4]$\ 
@=D:*:2BAJ2AL:+(HB.A!W6G[FCPBO#5V<N@;?:Y96=\ 
@ G<:L[CN*_W .A!8Y5AN$RNYZ"V)O[B'D&:N4W)YH0, 
@7_1<7DP7VG]:*HQ#(7U25Z3<X;]+)W3@'J:=5T=R\U  
@0Q4U+**D[>NEQF.K?_7>%O2K!@/K-,MV()D<0QI:]'( 
@.J0TYT->*39#Y9-2'IQR<W\RW&C61ZG'-6Q."6@LLC0 
@L*'W]1FM@91JEC-<0W T%#,>S=&2U!RI# )EZ#(^O?L 
@K@)DUTC MD=]M[@<ZC&5.1YB]MF]H,CRUS%:;_2F]]P 
@8/>%IBSE9GC,@!TZ__-KZ;^AGR]T,JQ<#P]MZ:_QY<P 
@&T;8U#W7K?SJNLZ".%$=#L$T7)FGOMT&2.YM WEZ&HX 
@BO,;5%FZNR8P8YFF,1/5U;IKA-[2ASP5C\W&]]6$W#< 
@O;RYDO 7GP'D'A".>U56BCJFL]6PNAA8;4=IGWPF9=4 
@!&N"5.,@,EF!-(Z1!O<A3E3KEY)YO&P.!_:&N+D9(WD 
@J,KFK# =$T^HV):-N"(^.:GK+%^EMNU'.<@IM:\_HFT 
@,)#V!("T3$";D<J(UFI6OTJDDIM1!>';4CG+D9JS'+D 
@B1+0T27%"^4/\Z_N%H<"Q(T'GRXT*N8OBQ($?9Z4;*P 
@\QU]X.O]K++)QZZQKW&FQ9 E (WFA,&!X"?*-I,Y()D 
@0XD]J6WBB@=BHH)QA8%%F"YI*?;_R.NATY>:X8G3(8$ 
@Y-,7EY@3"1-:7!TMZ.6=NU10>D_[TE=]N.Z+Q)Z@1 @ 
@XT/FSEV4S#  )+ J=-(/ :F?=9VE!215D)%.-WQ[FY< 
@=33AE"P16D<-^@BD+KDG9SD>?4<M&(5*:R"BGC!@5)< 
@$N!6@2D*U#'QA[*D7+;YI$T2H3O]EZP?8+ZA.T5P\4P 
@" [_GE=6/G.:1C&FU, 3Q7C2E_%)]-:C*N-H)>7?)G  
@%5YQ4:.FM>)M.R%DXN. 5&7**C+@JR)@R,Q7@0-^]KP 
@S)KQ8-X]8 8"QC!2H%S*<J6@>G-0UCK.G0O@SY><%-< 
@5"<QZNA-,U*/=%.'B<*OCAC+2.+[<]@PBRL#QBL8%'\ 
@*H\ T>KU)08Y+HJ!:5@Y6!^[B4J#._EO:ZY>4(#C"W@ 
@> NL3N5A[),DY R[E).ZLZS^6+3]&5XAT=!:.Y"*+G( 
@F_Y;1AC.;M\4K6 !O0[:*"G02I+69#I78?$[0>8BE0D 
@-&+1.^C?27O\GBARFCY+@^'%,6"<-GE*A-]FY9WHOIP 
@U**@_',*$Y/#]@YP$SZ&^&TD6&\(54A7NG_P[M[B8!( 
@692,/>U-.IBOL;;ZVPRBBUVL] +>U=GJ%EVVRF_J7LP 
@WKZWJ8G+8*\6BUO132TF>4F#D%>D+]M7P_8#?%PW$?8 
@$'J8F*W!:PW[E68A5'?\_"!A)#H#$VC'OI,^MSP&;-T 
@@@P,IE:E5FN/#(<$(&#HT0C@E%C][LX>ZQ4G>1AIJ&D 
@G=#_R)MD;O +R/2>C2-VD&=@N%.@C6N..CB[\Y7M!'0 
@7_.$Q")N[T^,@HL4\)?DYE^U_1L5$DF[/9<K(@[)37P 
@-8"RQ<ERIL5B/B#C8^N1!S?:;GP\0YS=8I&V0!!32:H 
@+V-VKM#2SDAI_=78C>U<,)HJTO5E8/A45L4X\B(WL#T 
@ -_86PV6WX>'03XW$,^&ZTKI*$O,G5BL2<9(CA;2)2$ 
@W")/),$ U^[DJUP'"!B='AFB)6158UN<B14/I _<.(\ 
@P9/+WS9.:KIC.^WM["/,L<A>CL88$(PUU].@>&9 .FP 
@&?,95>13,N([)]?36M$>BH;Q.)D_X4?>QQP4+SVVSC, 
@SV:)U.3XHXUJK_RX$)' G#QZTTWY?>ASUW_V^G14A3< 
@$_V#W:?3(;7BWDLV'8TFSX5B>#M9MYR1$)G+>*P<)+  
@E%6]*X&E>%S1E?K#.06A.T,'DJC=Y.LN]AJB9CUX#>\ 
@2;8-SU$T@@><L9<=M//C%8ON(1 XI\'3H>*<A)#S[DH 
@X'L]>2X[*\H>KA+<LUR7WJ/I>@$:6*":EU\M@YJ==Q8 
@ Q')WS2P-WBNX4:6+!&XFCY+C=[LZ@&2(TLWD IM#N  
@87.D$R1)\J-2&#*M57+O1&C"+-VOA;SP*1Z?V$RR+JD 
@BHH]Y> >!TO>9U(70?]0+^F;,/@_S<C)\[K"!07]-I, 
@ZRB^GI=@$'H/_2,Y=_Q/-_I=91_0)2/T=M($! .N\R< 
@AV?&J5/%BUAV<BW+Z[A&:PX8H.X_NU\F%%YYI1YXV60 
@_&WO@MT"4"R!J%>-.&[]GJ:HAR@FSVR., 9<%K%/_E0 
@YOD&(ZPT%T2G(53/<39'M1:3WA4O"U=0D*\(Z6G.51T 
@:7%38S; $Z\NO!6#"#P[%2YW?4-QUS:6==R*PW"01K0 
@@G*Y3 @%H5&_ &CY/L12&SC5%-=]4KSY]!"QJE.B^#, 
@_J]_4VOT\$:0_7?93?+2$3BPQFEZ02.I9N*JY'XIX!D 
@GFF.>'=PR#7#M<B%NM-^&A:6BN99$"HG;UX=D]92[WD 
@V"VV"H:%&F&8RKW5ICJ%W5_:=/1Q.LN0%<A" @F(^D\ 
@]M;NV*#BR\]<9+!3 >[-O:]Z-+4L<8<WQM,5^=N%Z@\ 
@9>U]%X/+\JDJ*VX4GC\_/(RL737AQX5[&;<VHME<(H\ 
@@5'.,G@F=_H1_U_'61.ODRP^YIO"]4H_OKC1O=H#+;@ 
@V@DF^U3XJ2&5%9DGHKR]#EW?))5:-'W*I"=P)?JVC_  
@%%.9K:&2H^OVX^&VA1W:H8)% U,!SM>M5D7O7:S7+_X 
@3Q"+1/\S *0_"\J\!+A:S_ ::"FHR5%>3I(ULXOHJZ, 
@W8M.WFP'+Z</L!;8V[ULO6Y;\SNK:0E!I +;;!QRU0$ 
@ G>67#WUYF]M\7*B.ABW,-GBZIZY:IA7LQ]<635UAG4 
@-D6<O>55H+F-5H<=*88I267005W-6VKI+@@6H,'U7DP 
@]TZC<RMX"9N7F!#]:]\:*"OIS)Q7'E1%[6([.6EPE., 
@K)(5,!*HXJ^Y76^266D+_UVR3 ,2DO:)B%.OZP0V4+T 
@&RY: P)RT37>O ^0Q_0BLXE:?("+T1O:+*+$^!@53'L 
@%IR7'9VCO_?IM;0HE>5NY[Q.&_SG(XG9/IH0YGM-'@\ 
@.8;B55!"D;/T_K.X!ESRM7&614;)RK(FC-VJYN@25(( 
@^1<8,RYX'D;W^X3"#VUC>X "4S^V?"-A]1I^R2"UPCH 
@D:P[)S>T040$L.W#,!N-)C^ <=8/T\FC1SK4^TB0$]\ 
@J/O]Y&[9_!)5_(V/$>KL$X$05L&+'+'-TOLD1)<<+(< 
@^R*F[?-8;@@25GWPNYP64;NV>=M%%H\HT6QJ<8FS+?@ 
@>!AO&+, 1Z(]WI-U*-TFH4G$Q7<$PV"W?&W V>E/K8( 
@K LW5+O$C3G-FRVG]C+>]HZ.7?IRY+A@3L[\]9+^Y\$ 
@6\R87!4(")*%UV$W?D?D?_QK"*"Z;J]WK2D@VYS_8T$ 
@>3I6]&H'=I4I]#L WNX/0=E=/]3A>)DW0/[>W/!#^2( 
@*P_ O31OB>6(_M"WU/I+KOWN!/PUE1U5"3_747ZF538 
@));5"_#4RF1#^S;&A-_]$S,#_YU" WH%%>SU;$_#'P@ 
@2^9E)3I6(@%J[&[;Q!KWTT#"[3V U.0&!77(D.M]6XH 
@D%4ZA3_;ZS9]4(2'.P5^Z>FZ4_O/LDDGNC)\L> .F7H 
@O)?FRR_<I[!GFQ=BUF;%:5??KBRV#$1,(;-O))93,?D 
@._-TRVF5"J?VE7E\0+RD:6[BH#90LP>!!0*A_Z_J1+H 
@N/[Y!@+O26HJ/0QM.Q7@U\6?"HV-.6JH4QB4N6F--JD 
@0<X"'JY="P)LT\U!@6%5F)Q4/!9W)">F(ZBO5<??!"4 
@\_%1-J_RZI?T%.IND1=5*TR>97YRT+#=P9,+WH*#+Y, 
@?]8>#2<QD1B&Y9[^H!2+QQA(HKU8_THLR:)H4@M_I:( 
@&0Y!_/(?DCQTZDV0R&?[;$BOL\=U&0-&VJ:O03LE?[@ 
@AV3PM\US\R!9-1=AHBSO)U;X3*HD31:D%JNF(X3[+7X 
@BJBA5VG".!1,3Q)G/_P.(_'>1>AP];*5HT1^61V;Q(P 
@2DGW%J*.-1D2:PV/<CL6'&B8^/Q6_H;_%!-79Y-J!H\ 
@7S'P%(_6*0+M\CPD<XH+[4J@'V"/Y)((XKX>24QL?=, 
@%"6HJ);80Y P(6?[,#._:]303)G<]_SQ_>+O95C=:UL 
@BB)L;%PE#<V832PD23'B(*M,9SE%N6J+,_"*BUM''C$ 
@'QG9IG6HUV)136T,7,ZEHWFHV(63T6)&C*F%S._8.;4 
@:C6%'S1[![@7=DNY<;]9)E(W^6C&7 (&0[M8#+61.?H 
@M(/:^$G(@>HC6:S%CP.">JT!AXJ^;DO5Q#4+[83I%6\ 
@6T^*L>HUU(&W?@*T-DQ1_^9B!SPGU8.+'ZA)GCH:GCD 
@I6-NVRHO.8H!='_EO1?L[EC>F%B$^+5+N)?)D#'BXR< 
@&DVPT:&KX0H<IX6O?US[Q:.UMZ$:B.E]5]01#T9J;:H 
@DH_H^W$,@F!@ J3"W/WZSO6!HK\=12P? "->HH5A4*D 
@6[JU5.A%#5[3K8_<=C9;B^_A)N7KNPL2\#O#KGF<FQ0 
@=.$":#4">TY)M2S8;!S/^7+9N6 JB3:R>&WWJOT@T90 
@L^S5.4>FZ_ EK","]L!!$5IB#C=="%&*3B6VB4_N.0X 
0&.63\$Z+G2J,W.N;G7=\=@  
`pragma protect end_protected
