// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H=9MZ6^ ;;%EOWT-F\;TOUG^MO'KELB*F:BNWMK1*Z,1^_OP7Z*/%1P  
HOG"A,TAPH]H#GB,-)%82I,PAVLZ>^5!DD8&2P_T#T7YSR!2FX;X7/P  
H2Z^4 =(#926_R"@]:$1!=$ROG>$O3J]WO&K1T=@/06W79#"@_@D?/@  
HOE\QE#Q 'TJ>KBMW^YW5HA5<T8296GA9TV5C:X]=N%L76R,Z]P@_/   
HZ+8:3<.%G%4%Q[U.2[_GE3TYZ/2W$);\ZU!8*YF$MD729UX%*S]]+P  
`pragma protect encoding=(enctype="uuencode",bytes=6720        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@[U1Y[0^2EAB'1YP11"N%Z.NTAJOV[5?_EF('(W+L.%T 
@P(!0&P[8[DDQ*<>UCWL8Q<#$<='R8]";OXMN/T/^]_\ 
@]X_,YQL72P87Q@S0N>*O_;Y9AN=#RS2)_,R(NF0*;6\ 
@Y*#@XN>6$0V)_#-[;_O>;D5>7_!K;Y=L5C4'MY,71UX 
@Z\I??YLWU]*)(=T,<4502&!:$$S;AHI@Q,<4&4RF/9T 
@!\=BJGWFYH;.QMG7_)W7>&86P%@9Z$_%F0R31B*:!1  
@M=,3U#W]!?^I_WKZPOG@VTNVE[Y8E\JVOAK*R6^9JTL 
@'^(<)UPK\P8#ERCRZZ_E(A@+59'V^5@LE>HNE5#$@J, 
@OGGC5'ZWNT,D:8>-WWO.!AY  XP\'3<-V!;.ZC%8,G  
@O!303/XH0QNJUYYZN"*%=Z,\0+4[]991IA"%IPAFW!P 
@Q%PIW9Q')]19]N5VIF>M-W=;1Z 9O$!GHH'1N07"$@\ 
@]4%U+M9MMAF>X%S,0*I'2QZL!O%0^G=B"=J&'ETD<A, 
@9/',_R^7#IV/PEM4P,[IH(<X8,Z,(&*VV?U7#R5D\-D 
@DS*'I''AG;[R5:"<W%:QL&]0#[-ZPW5+C?'"TONIJRL 
@\M.,_02^!%U7.?:Y%&#I*D3@+O& !<>)2BR&D\IJN\  
@/3(\Y6A;79@?=+*,:3Y./8X6S6.=.1@\;<RJLRA^<5\ 
@/ZB.Q2.SO1!]<6*B5Q%I"."]&XXB.JSP'A4HX#!>J_H 
@""A^_&N+&;,[I_*Q)M)7(?Z0*F=P&&6R,TS*3#HLOS< 
@>J^R[;>]"37Y7YYZA3ALEU"](+TLWSJ[(XT']Y[/RW4 
@!<(=\6.C+4ES4RB/Q(P&/,)'M#6<C*]#5@@[Y:[KV>8 
@^ X\XXG&<&]7435CA(#B=5-W%$_8&DZZ0_R.X>P=^;  
@>$V-Z?]%-MFKN)8]J[JAX)I_V@\T3%<[B/7%M=]G)-H 
@];;KZTMNCR_]+>R_U\OP?^8Q\VMC%7=SY3'CQ61/0XD 
@S9@ /T&D5"'62$V ^'Y@40THQD/-,U :FAI%?!=MFJT 
@\SIAGU:=_3V0G#?&VV2B9 ?SKE]1M)R>HK4R0 ?Y"2\ 
@%//Q#-CG!OW,>CR$_',##]Y#.<S%1 _QTE!Q'#5#'N4 
@#)"U1*W=N^/)X*/*J?H+<G72=@$1]C8?;@-@;?:<PHX 
@F$O>Q2VY[$0QLK;MUY,D3CU^E''[*V'ZB46 6$=!HWD 
@\T71PQNXSFZ?>!BUJ*26/SGI-88Z/OU@NC'B#H/_R%  
@R?R"<Q]:J%T47\B[KX2V)DY,?B<^,)15DZL_6\6UHA0 
@B?WQS!,LGW'@"TTJ^"LR0H60\_N'I^:T&6_GCU (FC  
@Z(4NY5.=A*M#!WOQ__;H(TE5$87]X^>[G.,8BU2<5', 
@R&,G(@K@/3F89J'HTG'#=73I43M?'WZ[.RXC1N!@H$L 
@Z03QT ^2OIB/\N;Q+E8T?D"%&#Z(93!:[Z!KGAZ(#)< 
@SHX5_1VQR^6['Q7="N3O'"[HP7JE6@%5*5X[AM&T0CD 
@>.P&S@(SCLHS)]LROSV""("%5.91BD"DS"YSSO N9^4 
@N=V4H6_@7UZ]Q:8]K5OJSW4ZCN?5I+35Z=&('S1$4#D 
@)\FM>2UHI$D#K&-#T=<E*A@Y\^Z;HH<%UCQ"JMD$%HT 
@8:)!&;R@G+@,(R8M(Z-YG#:!RJT:_58H<W>1.PY9A^  
@Q5.G WKS(7.I$6V.Z(]/@I/Q,J'-',U&A0_PC(7H&NH 
@JZP<= (9L$\A[ "N"D'>>!:ZNS,?3A1+QLD0"TFI^_D 
@L)C^%KK6:$OKMU(W0B;&3B=]]M@YN#$PI/(/%3BF^R$ 
@4U4$F>A!>1*MM_SFT%*W_\@N*N-'M[ZK\FWH'<PZ?T@ 
@!:;"UHG2GMC81H14IC31L"<GOUV'TO_?,UQ6G9+8(NL 
@[()G!T><,,/C'0"BS396.S=4LE)P/,0"YND1\]UA(.8 
@H-JIMY@^"]<_A*9O3V?:@(6CPHDU'*0AB,\GB!W!*60 
@,%,FY]2Q6_LWCG[*_CH*FO4KR3(4S85JHWR_+7?^<*( 
@<Q/ LTV/XM\S_E&=63XZDD7>]=K,I-0UJ;6\;EKS$$P 
@:UJ\-*="B%J&U')X**POS&1%HNO8!X7EQEOY ZU"3=@ 
@3#K" T?>43PO5-S]L2EW6WD]>J7J-.CZ$9=I4&IQEEH 
@$] %]H=#B[(;1S3T.>'/4R]Y5E-(',1DD2,/M,I6>'H 
@=JW)(S^[&JBI+&2XF:)0KN]T O8K8Q,[OT#068!VEY( 
@X G.IHY$!1_PI(@Y?^:D/>6M,#DL^$I]&^T#V.IU_+H 
@0*PUI?7'9TEFZ=E>X7O?J7;FJ'9$5"B/URML3*' <A4 
@ PO: 3X8P^VCSB?)+X=7FMDX5@T3^$NV@R#5\H?:?UX 
@%J\[)@OXNY#91V)1OJPU+>]P2OY&2HC: ]HAS,#KU0@ 
@%H-Q@B4D<]C&E!1>[[,H<W=9S^, -T1TE63P3<J-00X 
@-,B:]*D)LJJA!!G!U70GAX '*5]<_;@@!#(LJEX/[$L 
@.)9':]1OTI\<&BJXGWOF;VLH?2^\LK ><"-?Z_??3N  
@'6Z?'LH/HE'1G,L*P<NDMQHC,SL[:>L %RQ9FY58UYL 
@&.;#4 9X=T4/'@_USS./6\02 P(6J&;QI L)_+[_\=, 
@FM'^V7*48MY74(_T;R+;F&_,I%)"_,])KUI/KI)QG9$ 
@"&GBDI=VL;[_'G] /([L0/H,:'-K68Q>F^Q;L3/<'PL 
@<KX(K-;MZF:EPV&J5A9;'W'8E?E.1,9!.]^,8$F),,X 
@E;E  ^NB:IS=!'5_I)<<+?3J<A3-(MQ$*MD4U,,;$W8 
@1E&GZU_*,9::,RKW;8<A>;AX(IE.];*^' $V'TBE,QP 
@. 5KI0@I7O1[T<L>( '>(W:B&"\?C?D4U^ES--/I4G4 
@9 W,+;I\=F@N4')7).QH06R@."]HQ/9M^MZYW4!(6B0 
@_$HFPU''!O.".=_6%]J^7G>@70!<=J'9)K'[$>@7)PH 
@D0(8Z;I33< ._NB-H0'*7_QO>=?R Y?I<&A.T(^Q8RP 
@ISN7I"VTD3JD$ B/8'_P-.:WJ4&ZWI@*29ZL#?W[%=H 
@SZ&]^YH>(C@BTFJ0;M50N*G(CI6U:I82,2%I4QX9^S  
@OL%@1-RXPN%KCUQG>D^*QJS [B-\@XI9&,GYGI\W=U( 
@R(H[W'*!?H)RB#5,-5V^E:IJ78REMWG]63!-ZY[)]Z( 
@ !7E+S.HR2!"YK?J.-5CZ+-LE<L@#$(%"%&Y ^DA?H4 
@&$[>_8421&2:'EW/D5%\ZA=P-^=7 AEV $?A@CTZ\O@ 
@WJ&MW#[#BN+$^D+F9VDN&+Q*,:[PV[ 6B)C4L?-]:+L 
@>N4DR&N0L"!\-PXP[;NVO]"25/RF=9PE06:==)_LYP8 
@E-WO:>/([F(#LY4@MW@"$DA^6&E"M,.[6$HM8;#[/S  
@$<:4TB2^."=!='54ATO)U(CL1%>L<EPDYVQAO_*W5?L 
@*L<9;ZW\G_86 FJ\0P8)[^WQHT^&#5"?6MA2XN$XZQ$ 
@>B;SS:P&-6\R+;G]MZ-G&%$@:( [,;2Q"-=93T#5D@X 
@6]]VHW.,'(2CV9DT4,&AO=(NNC$CMXSZ2;=="21:2J0 
@Q\DCL^Q<T1E'06^_"L(J@8D2 3J<BXYPRH@GUEU_Z-D 
@(HU"2X/<$3KL9GP'9EUR*C@F9U3F[WN,UK(C!1#ZVP  
@#9U/M0#8*7S730.I%QH0,SC/?X"*3O3.",,A_A(G.$\ 
@82YK?<K&.*R;2]&6=535U9^?VXB>P'C<MZYJ0QBIUDT 
@L)Y3#D0@9G\MKQ0OT/&XLKZ.!]6 4V9;Z;T;%-!0M?< 
@\7^.LU'2N *[J+Y[.6BLKG?3V\-\:C:38+D4B*_Q]^T 
@N"'G&3L=AO(H(X8B3E81B?H$:A\#Y9)O+Y\T"=&LH-0 
@[PF.F#" ;%=/QHGZ9]59($**RRH"0SB?)%/1@Q;_DYH 
@?-I\-&%EB_%;F9_4?8*H!6*VI>HM@@";_.[I:IOQJ&0 
@GN5]]JOO%.8E/X?B:1?L2&J00LINEPC3(=:TQ)% H]8 
@UQY(/R.+Z-/)E@Y>\)_(4*;,.'R#6RV?(MP9B^F$W*  
@8;Q**FWWQ<1P62=&KME2J&FNC?U>F($+TB: C]6,XR( 
@]N[W&@L0WL*IDOO-3EK9*TN.QVXI@$0(">+/ZJB.O(\ 
@4QZ3<!ZP*1ZTP-.89H:;Z+10SBO<0IUCYJM%K[S7JBT 
@C=9,D ,X MA]Z^0V20*"6HP>TW\"(J8FA7WTEPX1AC0 
@GW4=9'-;;N>LO;L9)$/"6G!]@BN$[#S3\]$:(*4A!:D 
@Z5J.<'VRS$$$;'F1$:&VMQ&/5L*EQ Q0&\<K<Q!S3N4 
@Z_R(SDNPTQ50,LY6/J!M,<KPE_WIP$7RDW#S6NC8^J8 
@)VJ@_U'(6(!DOC-IRW\^_$I?4JNY'K;EMSSUSY^C_=, 
@*EF!AJP;PKW.'@SD*KX;:^]*TAOF.O:T!?#[,]%5J<X 
@* 0\8G&$*VOE\%%\6L$XC?\C]P/YTZCV0".A?5RU%-0 
@B#.A5RK>J=,%)8#> PCU2Z<?>FFGZ_U H!C\9-1=79H 
@0?=G280(:NW"(>U__/'""FZ?__P^%+P$UC8HT]--P)4 
@ B(.-1%=-GZ1/]_EB-N+*6 -R9;0 T+!<YUAWNW(K2, 
@S>EZ/@F\D_R; ]BK9Y&A:%F(^Y@8!;Y3JR??#EEZ@AH 
@C.#.@'8QIHXZ^R&O VA6K6!_6@%B<P5R0 "9NJ;N<44 
@@3EYAQ%JTYWR\V!!F4OQ2)):_6N+'Y@M+^@DB]NZ#I< 
@&^NQ0%.3V4]WI7@2,<;,#<E##[!1NQG3[W-S["R/- $ 
@<)(58.H"<FTG&/-UA'5:*>3]H-!@$1+?6)FQ;@QC\@P 
@Q2&R\8,%-/IG10"#TSL_5OBP@!("&%3?(G!%-/=]F3D 
@]44"?3\)>MHTS;V>/(/\_<&#R"541>>^)JH"XG9(LEH 
@N,\-RZ\2@=4RWE:N.$?_B#Y;AAUH5V0M_B@V^/UC&T\ 
@I&A(LYOL$UJ-_AA7<\J2%/CD](3(G_ B>O=?-!%YOET 
@B6HPS=O 1>'85B=KWL?1SX,WJ3HL!47_2G1H&Q MD_P 
@*X:7&ESG+0'F#0[:*K];S\#F3Q3J%7[;45'G6F@1S5X 
@4@G0;=IN127H,C7417'A!@$KO83+5(^N%TY3^5K.\;P 
@HP9T)ZB0+L["D'AZL\.@V.27&ID][&JJ.,1ZXM J?/4 
@4LXK!3%'O,$X7%MS6X* I0[)P5R5&WB?9U4?)L^1^48 
@8>/Q!@MLAMHNPM%FFEZY(!=7=P]Z D[)^T5QQO%\24X 
@*J_Y7X7E9J/;IKLD2UYK[-!U5[ 3G!<WM\)-LW]RLM  
@'Z$+,MC(;DZ2\20WEV3V+WY0\\,'1;MLX3R<%4(#<LH 
@MX32%_ZG]0XG<"W&R<4%! .#+/P6Z\OKXIUQ:(B<]F\ 
@E;2E^(OJ(P>Q;#E"+8C-\F'M-I#);UJ"F97 4#,2X?4 
@5DL6X9&&G?H#.M4_ETX[CS@?ZN4<$(/W;<']",[-V*\ 
@X_[8NQT9R$*"F 4EGZ=T$^HF)C8V5 ],;V:+P].:5/H 
@'SE.1]6@'1RD=26+4YL*6L#0KQ[]ZR-FC(#EA;G3)X@ 
@ 0V@V_S\E^5T- (8-L78BF^[JZQ*=1_ #L^[WP1&WY, 
@.QKWZ==Q$!2=4/F+EJOH(/F&'HZ2II4F'+4@FLO6[J0 
@5+NT+E?071479;.%+^K[3"\;K/?U^#/NG.!*H5FTHG( 
@V0<RO0E#H;>]<SJ8%(CB8:E$Z6/')S5J9EXW\PF4?'D 
@EBR28N6S";K2D3CR#JR/#4PBA"\/V#'>3>D1+UM<R?, 
@4=7Q(UFQ5CXNXE[I(W"F1Z'<F" ?WQ8><7<;?455%;@ 
@BDJIF'OV^^6QVED#].$ASK.B1"HN=+7$2O/3CUSM9OH 
@=\9"S4LV5?FQF9HP$KUQK!3.F>*<7<>I6Q.I)J!Q-FT 
@C1S[[(40>C^EWWZ /^4216J*O01N[.[Z/B"#^EYFRT0 
@#7:4*I0'"W'0:=#7;P#_<CTHT]L%#Q0!:O]HQG;XMY< 
@'X>T7/2Y0)%0O/6RO+<GGC_,I8M5FIA%K+ M<W;S95X 
@S\!<,L2FWL,KH\$C9@E)YA'+=!O>(I6HV2FD_XD1M9, 
@NN"%Q)/6*+5TVT;MI?0J[8N"/DK9FLUY26ZNZFS!%AP 
@*899X E46<F$&H5$Y#2;$T;Z"EBV>YN2LV,P/W/+H5L 
@VP50E)/#?VD?(*PYD 8;;-@L/M:.#*\>1;#MDAA4&?D 
@# 5OU(P2I<=4XUS'V&T:L[;>]XW-9J!D'&_SNH"W8PP 
@W9J0R$#"K2"J+7,$1 BL<B<.9UI/'5J'4S:WNY+4!%4 
@:IG4ST(SB"EL53\K4"O3UYEQ,Z'+# 4RB7HI'EN^ *P 
@Z+68ONLJGE@/-P$J#[EL>-$$%DYK@24M\'D-5'"<3_P 
@$3N(%$9,Z^$HN6D4/S*AZKC!;!3XJJK$?0RE6;.]I3( 
@D?AK'8*$;G"( 24#U,2=8"\VF9H(R".FL1AB@(12)6D 
@2?!K0/JD%V )"[O M[,D FVM_,WX&+_'%7I')AGGM<@ 
@FPET;*(E9M#_8:!T%',4H".(4!X'*QOPW,*891T=]A8 
@F1N99!RMG/YZ8PKXJ8I#4[H+':_7]$X1Q_HI0"ZV/$0 
@);ZS]HWKE^24S&F_E&'%_L<1VW_72UU3*W%7)%ZSFD  
@B"=4N/N*KJYS4^6ACBL"IV32)1B;Y(YT'J"+6SNQ+W( 
@B]H_0F=S']1.0)%4'^>2+ EGY*SI2LC779QVCCX!A84 
@$A6@ESE^[T/%'+@^%AAU'^*A6F'Y9<$&L#/Q]S74L=< 
@IM^:V +9_7!OE*R-J !84Z& *L$Y:QBA1Y61[P)3!%< 
@ :^'+!)%32MIB&.I6HUP2)J> \2@.3M_)O$<76$"WZ$ 
@-A4#:]/,[;($9:H$[JDX2M#*LU*X8H>;83/<M&G!W%D 
@&3%<$3_&$@T<37'>8<<%.A/S4&7+?:OW:\YD49F,9W4 
@XSQG?<.%I64I,#8WV!ZSXF\KIL6S=GX<0<IP32@\-:X 
@J7?3#?YP/=ZFL''O@"130I7F^?1UK0KSI^H$>O#_X+, 
@@Q_+K.W[APV/"$P_]Z@ GY->U7$<<;@UI<,(TQ&!Q?8 
@2IFLQP=]:!<3O/TX#<@9O\'KD8J;!FC;:XNLET&$< \ 
@J'23_-:CO,LGU78X;$S]\T(A;T>B"OY!UG9\_M1! ,8 
@M26#8)=8A15NC"X_VVR:4]+J;)Z0/>P!]A6\[';*'@( 
@(N@.AZ=H2JE3:<)AHZJ[H^Q@S!N:O,*N:E5"8M LOX4 
@G3Z\51U1,9DT]D3EFJ^IL;CJNF"+CP:DU!J8D*+A9!8 
@8?IT]D>1R.$2^27O_K96"$\[_9]61LL8/9Q^I^=FNO( 
@&WZP@G*$WV5HIZ+ HLW=PHF,PTM[1 %KR8>4FKA_LC  
@2@Q5MYTGU, 7(SM_$]S1$BWCMH;J*<IR?C;21ZPH$&4 
@@]OAYODJ<8!45[U*) E*I\R^'MCZ&^L)@ZLV4W#'K48 
@YT+XO"QX/T$J:+3#">#LPX/H:E"!0BSW8!R&DSB/^'P 
@HYQKF$TIOL<Y*GIM\-!X?D""8C\'R%+JW?XLQBT-J]( 
@@ANL($1"ZD%BX  :G(M^>>Q@8THLY2:!)LVO^29*SIL 
@8(.V@Z^3K1EKOE*2V$ABXM^6?8X9K-*7KQ-4XZ4RH:T 
@>C#6X$Z/+,[Z &TF3%^%)&ZJH"(E8FAD7A927JS7["@ 
@WGC?VQ3B^'1V2MH4@@=<FTBL]L[!#&WMHYPLB A%L68 
@VZ4K2PP6E]SJB.^2D?H1?RS!+_1O6E?ZPADI5UY"]QT 
@=>P: 564Y26\=X?M?B89S]<3 HGQ'J1.=8P>[OZHS!P 
@T#]U_ !%'"/["-2Q-@3_V'@]<3PCT!"=8A261:^1E/  
@07K?F>.T1G4IIY@'OHT18K9@M+RM!5E9:^S?G4W$A&P 
@)Q6=>U^I38]MH,=I]X"2''C/.!>(E- VZ\0E$+#2L1@ 
@Q4G4TWEN"TO\^2\SGZ,26J/#PT+G4XNC8[="-W4]H($ 
@"QT  +NHJ2;"SI@3(>AO?J'GCU/:R)=1WH6Y:N7E56, 
@1O8R0?CD=L JT5JB/&L<,YZ:K#F-.%R&D,\Y6*:LH8@ 
@AJEVVU+FHLYJ.?+@C^YJ#D;J)]@.%EC^0"06%$-ZW#L 
@^T69.\%'./N 55%QA)@!/)5K!<SCKM'>)AZL-R CH=@ 
@7]4!K#/4_^U)GN_O6P2T:<RR5=BO76C(F'11U<U66-T 
@UBA['W?E^?4FJJV,^#C!"X.V)=A>!8 SPWJGQBWP\DL 
@DU<OTJV->C5,D^$EA8(V:@_UB_H*[Y_Y!4SY)>B2PD$ 
@B^H 3D&DDC?P#?Y$K5 O\5H_'B_B[A\_M;B!"9IA-^L 
@F/F?)_HFPV9"1B]HZ+>F813H@HL<([E3.$$?IX"=&L0 
@V>KJ+1ENC*6;[^1=J_?:O0+2FK>3ES']:B*+8-@F-5D 
@U$DGS+>;+HKX44QR<9_^@!>X)W#HL-5FZ7=3:0R[%<, 
@7+\LYUTXVBCB[YDHN,,5GK2^SD!_!%:/EB8598-*3-4 
@\"\IAGTU;EZ52_&3:W>;J(PTC<IY-_9<F<<GV0!&5)@ 
@R(S7AG+6<R>Z!"NAC">$5Y9\;/U38&58+/!KJ@+,98( 
@J4T]4X9O'0Z&A)NZ3..P=^^,7O@R"3P2Z(%%T?%K+D8 
@K%1BH;[O';?:5F B:'5YG/_&4#N?.L-2XY1&Q361F$$ 
@A-OYSI"BTHB*-D)?=Y8*PRA0>6&I%SZ^A-6.5# OB_T 
@APH/ 4J!2A.S\?]S6.M\4&'YMC*T)F3TN?KOIA!X/FX 
@C.44N!MPQ#S0RSN!&>QCZ4\M1$E"8XM2L['-OV\%6/H 
@0FD:MYWVFX^^]^J!#V+8\6 PENP'N]/L95/?4M)!)\@ 
@\DUWVRT0#UV0:'=\&**FV_X"J&&]6&_>808U5X\_*"< 
@9=M2ZH"S!<Y.W4+2I<G\I[AADO3XO>NBO N2,PZ1X1X 
@24[?!J@_!QW'%C;<E^.8@.S&]A],(O'D ]-+/.THTU@ 
@\?UT43P;[[K_5;M2844K-ZAY&*HPITB];#<^5!QW/?4 
0'O^Y [WI"-JBQPO"M5*_60  
0_8G4>.$6D\CFW$?2OI_UUP  
`pragma protect end_protected
