// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SmMZqkcw9vdx7ZF08TOj8IFssKQNYkTSmAkmxA0gCg2r7NhE1PQzGB6/ZtgYnhAt
gn+sj3q/3iuycP63RYwiO2+pDGCdGVLg0tv5auRf7no//H3/UhJHo/HJC2J3jSsl
av2TFkN77wGW4ZIJ+2xcdiyzdh5v/t9g39GsmJNcGrk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13536)
pqkAuIk51tJvc8nBqRuuZfxkplaTOqDpMvrxXnF+fAxucaUj39gCilgf47ykc1my
umziaw2xLsjLX9jtyDQLn0dbSQn2TXiXjemAjqI99s+hftdAD1LJkhc+/TkDPpPM
1Qbu9gmSNW05fpSXpx72vlzrf7Gm23CHNmWxHIX23AledzA1r+2U6OGQx/xeoBBt
OSJWvT1nUDUoy5ASU6Mxrg2UQ5+oLEDxAUDKa48O/lP/WDDMkN6+vxKbTOfUGX55
a4JDqYSkK3VDdK2JM3RH3PmJJnTNf/4TY9nPPV9v1pmN3/b+SVc568j6NkEZKYrg
0+FY7paQuM4SkAy6/oEeZNmyYjSdZzrCIs5KDbqFBH2pUvtCEhu+a6rbDZeywCB7
CJyYtOW1O7/vDdw8FVSdLvFMjeoHp8wo/i1b+cF8bO7r43+67lAWZ2saps0DlbNM
7CPLCVJzUNuJMl3VDZOl9qb57JSwZZXWr2z2Dk27chUWOn2+NXx1fjJFvUrH8qG/
kOk3C/SBkUQXnrLxUa3VXsVz5g+UVmx/wFrc7g/AOQWaJIHmjdDJYliOrPNqicVE
D+YeFxCMwSz+x8v/3mU/1JjHZn3R4o62OMLWpTvxY5wRcoKRnv+PyM+9uolYZnyL
1pok/hpIO1+46kb+62hSffZPVmnhzhXQCme+kQ5yO3N5auhhE+2k3yLpYta3yHFx
3c3KRRwBTswYH2iNweU/OpFv0l1JsbNHPzcf1PiE/s6qyliP/tJ8SyiVvJrg/zGT
lTshnonQdmS5QsG/CQVgLqq+jkruIm6J01nVqwFj4djxFhUBFBK3rDjHlDcjwEcM
CgfFXytx2M15MxTDKQwqJc0MHWcPw2ivm1Lmq3INXN6+hKuCitTRlgSQkyTBqbJx
CvELiIdJuwxwUvt0xkcjh9Ntb47FFRTs2dvO6/iAOT6enm+tYNiHbrrER2Pv9RlD
qek1GwLi5zGVLgSFy2REnItJ5phtmZwBZsNiKfVab40VNX+ReuvwyW+Znr3kShCJ
yb0gvTwOO4SUjqPhekO9z6dd9nC5XuDSHp3dxddD0dPc7HuHp7e2yOGUd4REAaW9
a3H/IETZ16YaoTSKtMCYG0nJCYW4qf4azqEyPfz1Jx8ZFT62O+U3tuZpp0X+v5MG
0w8Om/tszZUABP9xfUP1Zkh0NjKekscM/Yp5RIqClxTfhdRAQeJecku+EBU6ev3U
n3KXmbSXFGFgupsendXBad/rKlXuw66989D9JFLykyctHwhfh3ECyJssdDtBOdeE
Oud9HR+G+pJDGrvYCP2g0DFTOHXztjU0bmCnjTU2NGn/GwUM+OSuLe4C4jlz2E2m
Dp67AzBeKZvqDuliqbDgfus66wljbIfqgz4bu/br3cWj+iT05jyJWH1VP/8DGEOo
Y6jnEaPBFGXQXAJBdsHh87cNcXwDHem8m+y/zIb85J6wS1kgjUfWof1LCG82vqtP
aeEA4vhhoAI+b+t81sbBotgycbsELkIFXE9zfAnyc2lPLQe9tA5GCCvriFdiJ+ML
yo2NxwuqLJ4bxJN9rMKYlW49ynMM+UX69NCC/LxyFCZtGBEARQmGkf31wjLGVyBc
2C/Ojw1zVFma35l09ra0OsYlYzyn5hEloatwENt+CDorLNiLyibaHOsmf4mrT+Kc
EVni0K1HCKgJFpfdImOQtYFs98qlXNrq1oFMKTBVTbpDK028xSwPefzD8RomAvZ9
V2Fp5i0RAn681pNpg09yvs0Memqt0dYRG5yrbnyrtEX8/tS3jhaoT1BUJZ4fLbfN
DdgMiKMGR9+uSBMEyXq2sWR290R6c0FLxoloGzTsl4s4VyJSGSKLBTuQGwN9Sq0L
jyl7eGICuqpaFdZ7FdU+ti2YiM1Gs4nlv0/e7z0R0riDGjEbW7SIfNMAyTCKEDwY
0u3bOZNtc9OoG52Rpskl2V99s3opGYOGCq65rcz+L3kwTbDxkriCRM4nZE1/dSbJ
DvFgyETC3vlCfg6eqwMVVTCkKS1Ioio2lSfsNMD0twCLx30zGSqFXavTlJJwLdhv
8UjJnYak2SsLCv3FLpnff3lAgUj9ZehDpMCZACLhkSvHRi+VeklWeOfehGQnR+co
hQEqEbLQvIYC2ZnFUcqZuTOiLzQiAGiKO+mu56xV2RpKUxQqSce7UY0OK2J7D6X8
oZM+ZQmPM/amqak8oNEVrgyGlU9d0REO3kDeUg+sJDCoRHve5PIgiV0T5oT4ysl9
CDoFmtkMA2EX0mzBRumX6DAjiwKVylBHlzmx0exXMTdGYvqL4UuLedXQuaQadLpS
hMk4Gkpd5dgBRjVQsYQDHQ49niOYVGt5ActB8PqVxQ3UOAa4VdrrRX4+/8JC1J+J
oxfzAhNZ9zJ6e2GsVBAFWAGDinNYZjWaYn/h8neTRNdxVvze3YKOPCU+Ri9SR1rK
uJuQX2TPEFEmf9sDJ/np4Ryxuhs0O9OxoN13wlxgY+8GZSKCUCN8uTkBBaNbz6l3
kwCqC4SA0NHQfuOan6qPIxlI9DkOeWH+B33sWgtnRuW0corqszH9K7xx7T8tgjGm
aEpIkB032Fs39tlGPBeKS/yg/2OgB1kEQL8UF4Fm1mSm375/skmizx0AflzJvQ7b
K1WrrlYF1wTFeG4/P+Z0aDdUp/o7OKRG5+cFCheIVr02cw15CFSl7TNWIRaDvNT0
Pj33TnXHHRoP9/FnXZRf6fL+/XWZqMcffKEqzdLgUNr1auUICt1zeoQKQE4UDnv6
unYg8NI7qKRA3t12NKXjVgjDbwm0bU1Q4f7WdiMjsBYxdJx2AgS7Dh7/Jb5CIk4Z
+rIrWfwAI187Xo9wWnJ+zMCzU2LBfKepcLfF1fu53QUR2FqHVjix3BOVMA5/rMzm
qvrjOoSR48ALzkUxf+mxk6oxuEx1EQ8fLG6rBizQBMKKfiAouyj19ymqnnMBmvLc
vSjO847quop9tb/Can65DdsN7zO81mu1tRYyNqzZngnIZSecy0axHzM0ltLtnufT
PoFrt0fCUul9l8dAPpu6xX91Cr3gtXt6gveqYvb5zt0ODFdXrPo3vDuayUOb3Jyw
G4e2oo48XU9MtJlT/Rg7zTho7yWHn4nW2mvWR0Es3inmAZOT4gFkYkHLK+YAjV7p
/eNmtcWoIeSNch1+KsphTFY7qZkTCBDF0JOsnMqMdHv5th/dJUVRlh5PR/5QaAPU
siZttUXVAoxXqaZrCRnYSEJABbIn+Rln1WW4jvJLtyttaJwltw4F9dIcVmZOF8Jp
N6rQoZN5FV3atLjkZMb/hWlGcqgVbeQ353eZmjpmSLpgsoog3I2o2DvYXHTgIYxj
wNvPzJcjBRIPz3F1eZpAJEMXC1rd4E1Rq5o9t1osMqUFtfc8aMYcvk+yg7Z3dA9N
053anXWtdxe7AFr/7Adz09CigHGRXcOeULMRdyU41xlYBfj7V4kZ8Mmqx0Bn4fZ6
KSqOzO/0MVwg/nfkbL6B7Rmdq65ZTLP/1UNqvMTDG31hG+xEJ6A9fOdA5Wi6c5/e
xkDynfJ1v+AvdRuJnnNJ07k1Lz72aoaPqpY/15b1bbqP4LLc6JiwMMFByqjWf1Gl
T3g0Ho+8BAeh90VGGoUMcIU9CUU5iisqwIDmFrv0vlt2HjcuIgUDvEMgBJ+omAsr
kol0dkT08Su220jd9umkX8rI7uBQCrwtRxkP6b1kxEi7g8sKo8cUsmiVRiACdsy0
bjffa5YIz8oya4oEHEQ8wUkMXyd3zO+fseZHW0Iv+s6F3GEfPXe9WwOgqnz22G41
fh1a5ZV9llLFyWf8p5x1t82TF/v1N8RUCQ88Gmas+3REPWIFgTzctE9xFJyPevhF
BXTHEHs1qNEUIhlolPwlNe33kMMFT7P5k0B+vdWZ6J2VetOu26T8/Lp4lSqP+rS/
SBKpkKPGC6VpL6ZYbTFuSuLTSHhSUlq3ZU5Kg9yogvC2K6O9yd7Ubzu5IeA9JRA9
d/Md6986zK2KiUNynTyYHYaVP++w1m+jNLu8IOO2sYlGgcg6YB/LDLr5fnZtiX3E
6Gggt2q/L9ddEkxk4Dxc0obWRRCKu2ehYH/YBV6itdTKB5HKG6hWFZaOgtUuPU6c
Stp6AhgxfQe6+WAimab/Mo/9TFCNhJStYLgrKfQuZyKIsbxrfYzwcWxEUKfQznHw
qyIYNBmMQlO+U/QS6KekV0C0cyseGDtR1M8Hsf1wN7pK5ACgFFDJE2Z85s4E33MA
i93CQN1aB4TUqQR0vE7VXx5+2MjiXrghyrrI2gHhfKZEHV3K0cAwAOdX5j70QjSG
9Os6AVRKkos15BZ6UY9x0k02CzYb+ugYu64AShKLtz1ySGk1kmiEferkAMh/c5M/
YH6fTzqcWxn65ywBCKq9C3ObSWDTqceJnasHar7YmoE4Kz29JXov39d3wILwG7Cp
79CkZx52NR+NgfbNtm5uiy2a+/nDA71fffch9z+2jaZlR8Zsp58XQBDEZRGWXaN7
YWNNdpV23jIHwz4llOLG9QEnRBLCilcChu03d+Z24O2PBxY5GN+rqMt8MI7V05wr
t+WQ0mFq4eb40IGEe1mQfAzX2vYG6vlOaDrEhCpJUrRVQq+AKEzci8HdrvgoEIv4
QpfzsrMYWvzvXTMgkGsgA48P0Kv4VxD9jTH/dk8CwhDVqFS9zh/4u3C1sHvk4pE+
zGpV2HsYULP7wJenu4Ah560GZp0EsNHoK82uj8J55+KEV8lMBs5H/3Gq//I+RWJI
ryIBV/9G2BfomTlX8bFmSzNr8Ic4Cuv8FLmjfYqiDtlzO9qQaUWGXj1AbIPs2KrV
leYa6l2GdAd6z1wQfa6+HuQjMQSVUk3SXBj2zFlqQdHBVutyFfynni7boeVfi5fm
TM83Dt9d3ZS9PPZ4dx/hFs2+Pd/8LgirjNQypZZ2iYv60r7ZyLxwl60XAFrO47pD
69521a4UsI+qXiaKbaMyNVp8Hgsgp0+Mcn332mZc2h1Z/sTXZngqAFVzEXDfiHjf
EpnS5uWjUyOWpEQ9wYUvpEgPrDVGn/hYx6OpulTxjo7kq5Cugx2dvBYRUblWxU+B
On2C4a+3L9UX/A/0CVK9ybBBhR42HyKQHla1peLkBzSO9q3Ljvo6zCjSjS6jtE81
WasthDtDUELF3bOXK9J+aTTYMiUMn07kF+Z7imm9iKuMZzICm+9/FMXMoNrsB0W3
LcqwrnfKayWTtSo7P6FraYduUFymmISb246fXqP3rVl+bOOxQmcTHlFqmrNfP42v
Q2TFEuhNaDzIn7DO1plIlygpdamjYJDbUbWeFT32CS2YewgBwGLAWJBDtp6VaseV
JPbUgoQ6u1A2VJ5Tc62Gc3o0edODsNJwAt5S7wXfQ1JRoaEXaByeu2nv753mP4ZE
oDEYQOc7mDiMVBBtNY7kSVXiXnsJM1eBctMW77Rf4eRMF8fEiknYlm5jCMDN6gJd
b+jR8ISa1MmdKfnSKdYSXdJ0vo8XfPgDLYl2ykscs+iY83uJDFTIBxG1d7cyzJaR
h8VZEEaZJxgZt5FRChnI6WonXOLKx5Qo+R1wmjKJGmUCq09JZMOwm2ztrW0CG9Of
CJGwQPJBs7Om9sPmN+ShokCJArVbGr2X2y0VqMDcIcJrFML66QgQp69b7lSXtAun
pfWA+IBalBGStNzI7z8gtH8kTAio5ibz0CcvIxnefGcg1W8D4hrl/jpIar6/DRQu
/uyZCjvVa+47uXKpg78ixp+HJLS8zbAVxFJKcuvesRXkHds0tMUYVn3BsTZE4PD8
Heff4qeAQI6CfqPc5/diVdp+pND2GNgOMqm9MFSWuJXJs5vJltmt2yuTPJI/bjPb
XcVlCG2B0SiRBU48Z3ZZ7x+eXLVxmJNIA/ESNfqMn3YpWK+PRxgIPYgLDexIe+2c
+Lj+DNXgSkCCi3+Zf69aUSO5d6+Tyj9KtSFQ+iti3bJhjRIyWgVXxFFzVtfIPOrA
ejDNCKRcZjbBOEjjd4tn1wgt1C8si3LtLsjkXP4IeQpgKfSsoGNfUt99FpWna+YK
B+frGy6SxIjP4M8lIQHz1GEvdJ8hmRU+8z+fFJuI/YBlNBc/MpPJaRL/wEG98R5K
ksxF1NBdkUpnHKZA2gxnU2NeuzDwiK3IIFybwNLHgEHzAP+lyEiQkdyrvvSrySts
ZaTRBUONWNxavAL4iSSgvLi2HxeAl/G5HutaExGHZGvMxNKg3l15iAx/X0EGWoNC
jlHHkTYsLy9qNWC/Qt/QElkzqgq8lYTNEAPP4PYo+odAePtSY//EZuynyklPMxru
P3zFnOATk59ZGKXGxXJU2PBusExP1G4dGgR638JCV7VgPgk95/sDxenMJvKrpJ0n
cIj/ej0bvupmbORfOCGeijYhdh3RI3j+UAXQjMssy2dmEAHq1pAym5iBquD41pbG
WbpTQTK2WcIi4D3KbYZfNGYOdTMDS6xz5rPG7mHrS6QmmO0BX3d3T+nMK9xWDxpL
SZyvx5tnNSgV1o5mDsts4SGMq75Za2a1zaUU5ebDoTyhAJwlz9OulIwxM/8E3RI/
P8GpNtxA1eEhQtANswub2EE5KPnrn877x8UH1LqtOB3DcPW8L7sCILTLwBVeVVTA
3kk88EmUK2RNZrSiEszdo3/FQQJC13LaLQ46MTDzO4H/rvxKNouGbYlM4x2m+NVq
FkmhtSINxLFbEmQerDVewc1QFTqcpmFh8wetfJG1HsUcfA7BwJQ2BJ4EjsT2xKXK
QrbxkuG70hPJ+gQnzdsFhTPOquWGXk94uBUsf0WQKQJjCfOF3S8xZhKo2GbJ017J
8R6fynzMr1jaTKGPirT/I8pZ6BgIQ0kIz3oSGD0abQyqXWA7+LEvilA3101OwDyF
1IYXDBw9robFvfDsbWUF1kX+co0WM5uVCSygDi/QG+rdHMkdg8zjwVdSCn9AQ1o8
d3AdbMalM5EMZFIpfxsO5LLkTzoymroKN8U0lyESQD5yHSoA5OXkQwuJJ2K+XP3H
T05DVPLaWCArBhUiMbf0wz3mIjoo2TKQZZBgIfLBhfmHNlVpQ8xLkGXyqaiw+9Wc
aKseSye3iOa2z2ortSOGubf2tu6Aa8K0zftELrFAbxDUqnvZstQdmGZDd7pLrjJh
j/Tdv6mMQq4RCH6UnWfOsffuWHC3xG86N1/k0RIHrOV50nqe/U+Dijv0+hb6qToA
nQ6oSeBY6Zb07VAQ4RGcOynQzvBA2hymqttdwnbi6Lk82uqFIEZtza5kPJUesgmK
kEWxmVvvHgoMjwOE9KLOVGU5lhDfReSOnGqiMo2Olj1O6TieI/phXe8gR3FGFDxD
txa7fH3S8r3YtHyaGMm3cl9cFlRFLKEtG/xRFM+Fc52ELs2w9aL5jBz3uD0+SHjK
GLDueTf3gYxQ/mxWMTdpdoRJvAO1866uESfcTuykHWj36XgKSaSI65BrQsJqrl6b
6gjoxir+bhJ7H6bSMGHrEx8V/jBahlwU8M0Zr7440E0l574qqGo8IaU6RyO/KYLB
KyW+gIc1sSesEtgZTltMod15F9rMpp7Zogw2hoPaZv3zBr+9v2zd9Qlju5UNdCPS
Cwh1AZji6UINqrZW0NtpznKhIQxsufGauAmgXY5R+22JfM+rw+zuks/0BZ1dmoHw
Tq+Ue/LuUSR4kRRbZHjmRZjlrlb0hiibGkNbE0/AMGAsKXATyDM/MuPTtYrS0j3A
TspH2yjCW0RuSoEDjHCPQcZGo371bQbOFZrcY8WUkQQqTkKqyUedNdYlORff1LH8
QAhVQnh8LHp/JBXzAsrFuw1aDCTyxBp5ADlp7rbMHjQPw7sRFgM3VZ/ee3+KEKZS
pi1rYQ+8SqKdg2bQyvT5E/a0Uqq0v4h1l5CGjkUdD0WNtmLiTwgh373jyyBGXgr+
0QV0lkIIrzSxRTdMpqhoog7qavFQOszDfSlj9EsN7Kg+s+WTu640Ugv97U2ZyRtP
4JOtm5GSARwecLz1Oa23LRN/yaYjYs7LUecedUXcy3IS5V8xm237RKIoCvrWqBNt
06RBjhcQH+MjR0BuSvb+EI6A14vKaas5g6xtj840VAaNnpd0129XA2v5KbZpqUlf
FB0/GRl899AcRBsWpzSbBHQpbNT/MzQAjlD0+tQsAphV1VNEyxpnkkY53J7BpM1H
VdrKjqVvzDf2eXGtTSceQehhOrRXqnxidnkuwptffSB18i5bECAE/0VsatrqWC7A
tPozWxFNy8Wi72EgrbByY/ZAuuL29/pEEcS6GwNmw69DaBuZ41ZZ0GumXFnJFd5n
w0GpGRZFsAOl/JDOkfqGADCiegsvUrAWqZHCBT/xetlsK2zDEsYTEQgFH0NlN82e
GnIPLLjOUCdUm1+IZrVZbRhNPaav4iABblh9tSPJlrqyN1cdSafA6i4tzt6L8SA/
cLrOP/Yd+bDXhv9W9w+Z2S+eaipa7/g4/6kY1KqYN+LGbiZtfto7hyaKnh3Yynl7
sM0qxwxIb3g3qhhc2M83DmsU+USMmVCtiwqNGBzFNJCJJuG27v6Ka9SJdQLXUrtJ
pihst7ZLB4pWMaQH0nO1ILK3ge29ufT3xGvIV2ZGFkjfdDIG+vsoHJDN8lFapaOs
O2d3vj2tppPFuf4fuNrJ5JUNwvw4N9VUHjglPbZ4oJAjm56YCxi3FXmKxliFlU+4
XzwCZuxDFEaZ8pURkXdwWAJbIDdl83YSCRU1645lpenav+EDftuDl0hvagmoBAsI
6G9q16A5aaLMopIz2Jz43N7UcRquPI4WQRWpsYrYvS95/vnoxKFb6BSMBdB4SBMN
r+pw7/FRDqFsWNks9eWxSRYHcXcIq2G0m/ekQIHXMMyxDmz3Sdcl8bqsFtUDsYSf
fdWJuV5smMrHOHxujCHZRCvx+gDvB+By/NtHANNYaLqJpS1I8iugXJf5CYpSwqrU
/A8x1eLCYYtGfAdUUfqjzjLFqHYcYyZI3f7XbGVpMxgPOAP8VfNPmZDCKePCiMyB
F/RyjSbvFagd7alFDv+WCSUGgqjVmaN32DELvHttyVQtFqCjKn5Op7TRZPLXd1BG
NvbJV1juV1myGQs9oofbiaWx001lQxY/RJaiSOzlRaPz9ysw+vLlpnZFJS2yUgpk
45b3T0fXsEFh0HMnhAWi8jk8qqhw8azN2XaBEPeR3kjsPweb+CKpzTXim37ypG6i
ywmxdw4krHloDQB/J4oJ99YEN0QTlNVt0JWJLPx76S23grJrKZb90nip++xsOfbI
ZtaIzU59ZzGUAaGSAHDWHZASNPJuC+OOzfZbFggxIyJQIW1myP+OHRKaJF1B9cX3
9iWmMSei/aLVV2RDlJlFTmcVGjEPnXhEZu+cfPhcadQql/TQ6xnlAfAK5kJHkoOu
ggByTlaDAA4k9AydE4ieYMycr/ksDo1y0HdtHPhbTFgyZdPKC1Asy9j33957xRJM
jSW2anSqDuQksseH7gtjhunw3vo89GHTCD3N+ufWKVOoWBB5pKwhBGQmG0EFhEwK
FVdEufFpQYAO+z+BWpSG5omwD2xOOPttDYDBURgCc2qQd1uBSF3NCLJR/k0jgFan
BYCqT19WtWDYyrGfpk723e/Crvxtgv+C8VIrwt9veOb9+7sUDTuac+0oAH0sTl2O
QUt0QNxHMsWUq5v2RJEuxVjl52DEpJbNi1iMdChH803DhTIaO7xOZSLmC516dORu
yk4Vx2UO1qf9uIcrSLsj/90tqYuu5j0j7TwscmaErarZhfGjstw9Tm51RtwahlTr
E/Xi8icPRudmJpTurOvP67/dh//gp2Ns+ZbFPNBZ4l8xCJ4N2ynj64YYIzsHaYCu
XteOmGE06DKQlCQhCKR/HC5drklUXdpxdt9Z2Xd9Bb1vr82lWP+cjsftjWWSEWBA
eFrcKXDzGbCsfhqT1YNyZ6tz2bE7oGs41uQmNpAWLnlISRuQQ2s0XbdXfSqdCiUd
y1/TGbo8QLl9vWxeWDo4kWQ7Joj287uLmnFjSZ5IKCV2X8zKiAeZVMBo04sVM2Ov
/PO5JFuL26efma7GTAUSdMOx0RJ64re1jMVUQHIqqgQmVByYcfmMym4UOsCHA7Es
g/QuyC4yBXdmfPUHD8ZYX51s9EWzFISsag/Kn37nDRNux39eWELQvk51BAKNV0it
6kaTk0dGZLiq/q8Xc3ioq7cUhyXlgw33/tX4DDkoIwUesxCBZdpXVizvGx0vgMpI
NAfq/xk47+SMLu8xASOLD3PEIO5+t/ZNvwbo92lTU2PS2k4MLX1PCc7kO+dNRKTJ
mqWdUhguugK88hUQRJf7DBntX8pNTQUBG8RCiyYCT6aKRFw5v9M+heXQtMOg5KF/
IrgzUbnAH/jsXki82FqLm0HFsySNbOfEVCiJHfZ/9LwZrtm6otv/X62dHXBa8jgq
Z/Pr89uZHil7ZxMPOleSWvjjyEGY/H3YVhiHH92kNJ7iMys/P9/PenK8vCa4YJLu
E33nuQ1NheIuz/Oc+s+C1V13dY6dgzt1uH5sj7aMgkdQujfEFRcXNw6yM+EhU605
guLLjaY8SgAS1ofA4rc4h2/Dvx9FOfJe1oJxBnErzybrG2bJ3y7knSpeE4qf0Lg4
gcS181wm2DOAiSxQgMMXZ6xvFCmAuiaYNo563TRtdugt0maGJRC5ETctvyX0r6S0
kZbT3kzTcqBdtnrUsSEfmSIuZimWWWhKcgPHnPyteXlPkJ05SOHiSToSk+vPhaFy
HE117jgOlLGtzy+BpRqu99fWxNGuzVkyrTJ9KQDesYBmJzT33qULNRcsBI9O4hIH
l9WpUGHofQeoF/2J2Q5tvxPlgsWL2xZ2ZuW7lBRRtbNptltvs0b1xC1VI7vxRAb1
RBogYFu5BJfpsKXst6nxSivCj9SCYIQDQbNNkWu/xm9nKn6AB7ostOI1bStShtDX
fx0SNdz+G55J15XMstDmM/PsJSI8GRWwSaUnDXN3VwNzIwuNwclc5lFRLmNYs1O3
r5B0j0PzpZM9VldJg1mdrZ9soYHw8IjuSKulLjS+rvoGx4VNSZ21//SbK1P9sZpd
5XeWvKCeLWuoV68WhTJKN2UBYTO88OWm2NEJDLdq9bOVhYNphrz9O+jLAcFCvEXV
jPkXyH0i5dQzxNC0WLmIFf5XT/E1wiwfOG2TUw8lS8njyPZKc2SJhc5OmdhnH6Ec
uo9XCXcAMYnZVfVCsH8uzM5Q7NBLfqnJTL7AA7oeV2gCTbo5ipGIL/xLrIgXfnxS
qbe3FzsdrlufkdhhXO1Sj0j4IoLgCB1BFmenQtyjUPHJ2YIVognFevBNYRODPOkQ
sec4X7qIGaUkhzyXZZAeDJCDHLBUx5hEO+TSKyCOpuev307dTxdRMp51x0DJ2DZo
SUBRe/r4R+bHB7qTmAahUA1tmYn0HAzPVvL/tpPw/SG6wKTazyGigdHs7JgQYDgE
BjpUrJvXXHQjZVSMDCDPzRzuV4psM8/BhQbQdXyPbfaVJ9vF6LoYvgG6mKVBNMZq
nwYOtH1Nf/QMrrFd022tj0hD7aZnj2dh0wmttukf81mnASS6cUFJ7b5VbiuKwgrd
Ol7smqOrcqnTrcDL+B03McVIMew0qIZo8yN2ZdAVtDVM9WuOj+hMb2UwkwQUkmND
kF5T4f6vlJZp+NUbCSyiEN4H+RW0i12LqlX7QcvpXRyj+Ct4b5Pb2OFRW26ajMgf
RPcrh0RpmvDFov/8wwp8JO6uDA4NDXiYqS6q9s5ztEET4DGcZHUTv9EDGSjdx0k5
KYYUaDJM9SmA7snvrBv7jvErhTKGGfQGnVBdBD78YNCRcHKzq3XuXVDNL8ggUT3+
gpUNGG5ZAxY370kfrh6bGmY/5qmPf3YsgjjpFeosHvp+chcMgLV4EpXVPtsmRSqh
KIehLm7nCTgOAtk0jmPtLOqJ9BXlNu3l4oGNAJGl6r5ViRrePjyKAQgbEyB6r1Jp
Np5ixWbHTOPYoabKxWfrFTOyTOP2RJaMvZ190OHU5s/dG3ahCNt9VM+SO5YgUGME
w/KbYnb8g6CaAU/3fZtnjar1xnZ3UU6GgivVgMz4YX0j2k4wWchyelf38fwK3y86
IrSd086oxfVfeByAo3YKHh/kc0dAhHJLe299xVVmnG3qweq2IerVlqx43xEZekPV
pvBO/5Ar8tdOerCyJ421APzF0mAGdOPNa6wgBPHS/WEyUwFuqt8k+FnoEdM2O7iO
fZrAEabdfPz5UoWRaLuIjVDJ4iGuvg0s1qOAUv78vBqQh/KSCAMc/iUqC4ZaoFU2
bzrs0A4nBGCBnwUfsLmQLhGbgRNx1/lycruP4qo7nfRwWd0U2CQ039BaX2fwR5pM
2pQzQ1gDb2dymYVwmpTqjcVHTBPiV4kQX3T3nscM50FfRl/v1tOnUMHRhTIK9T46
735xYla3wCIa8Lofu8E9GnUJs7Yz4IFIvamNztnSJkrCDcWnSAN/K/qVz3X3+mjw
DngZF/tqsMGeJTcp5GuycS9YNTzkHzw88F0aAonUUortIdDONvGKyyA4pah345d5
CAbFdU8km1ffM1Qj6TPzZi/7dpl2+CzNeqF0jV9T1brG7dv6JfBJqoWdCD/2bgkt
GkQ0G/QuP9cAL316G3ZJZS72sndoY/W1wDuqobbHZ1RKu6ol9HOE2vPOKwb0RlA4
G62sjg9wbzsSDmcU51piMKaLVRaqki0cSRxzEFh1Xdx8e64bvnxCseU93MjPFGqY
nfqR6RSXcScz970m8GdwqJF1Qyz662zRZoWRVF6BHc6qtMijr9uvRlRnmmi3Jgqw
t1420cSj6M0zYgHue/9Xsdyv2usrF9TSv23DtmdcdDlijGML5n2lRPB8yLC1T/9Z
WLt8nSA2Gj1m2E+T1BUUyctsPa9p9f6NewHitXlkJCkFJhj4yypGjNqkZ3gD/6UJ
yoyt0LHycnkuepmIm78MIjpJJyd2ROI5CpglM7jIpbnIszl9psolECJv5PIv12He
U6eXRtVhEUq8kPAl6rAbujEw3aHYtpQjvXMzksEdBm5UrRdW3zjEfyuyiunUOib0
L4Q8t9CXrNezSons1kWXFE6kRD5clyTNvc9M7ND15Ee3mcOg54SW71+CA/y+IS8U
M/6YB8RWlWfpQRv4LcyErwDxHVcghnHzNtJ9f1OZAE5Io8adSdjrKIa3nJTYdglV
PUkm97ue18F2VxNbm1FxMBsyaUmEA/11dTxl3LCB64DEHfj/4prtknVAkVavgoTI
oUCShTdAojNoUhLr6mdtfK5z5L5LuDnUJ3uQwaq5jlOTWzVyFsfephR3pwRT9kre
zzRXGmVDbre4N4rsEYtKm/sjTB2heQ/L69ivcM7uqdvPVNyA5bV+G+DBEYXCkPnd
KVsgHXGOajUGG9V0uVsvNydYq7DUZNbor+F3X3AwCqt/1gJRiNnwkOG2I12EEt3t
3UdErhrIABhYtLXiS+sD/9yagHsF+PmafoL/l+liok7OUT8YFtKGQmSdpHG6WYKd
ycwC9o76cZ/1s7SPX3L7XP4Q7DhmvCvus6AyjckuoOm4JXwvYew+wczjF1qB+tJs
7aqn+kNqYSK4/b6SzLGryxKR8eBVR97zUBqGzLkvE7TjlzhnqOJKDvyt3scOgD/D
j+7W4cNtOZzW7UTtj/+q8tGp5ad/W228ghgCURNaeGNuRIILis8BW+OXvscIjNiJ
uDq0P3DZvdQUlfdMMieqFKUdpD359hJftsW/eXGw0TjGhqvyCO3MjldbMEalwb2C
JCTw3TOvR/rgAbQfoenhbVnVkSFUfRwcYz2OY5qg6BYCaQM6Ki5cV03X7Ol0iChX
Ac9ys59EcBJPM+bIYEcvVtlmhsC4NtcxN/TFquqqZP96ZJJjc9sDnQVWMhI/QVwH
4g+LGKe2k17PnLd+0nwmY5IESyZk/c6YjO1Jq6JjmEYWs9bYDSmOLjG75LS8HCze
hpt4kh0jlVGbdFkAJhRg4wtg9sEjoVmG9xoqZi8Sl7KR4HcMWLL458+0z5i6xyvw
r2g0ZUgyurrG60fpFsJc2bXrKzQEXjvVhEKrXlM5vgKwZVD69gHt9o43CKTzhe4S
9gfg8mD850GzS1JOOlfBK1RiDZko1icLEYkDWGsKGFbR3MhrkXaMFM9JB14977Iz
3fo0j2qC4As4WcXf5SxdqpWoVUZepQ9bLDEhJH7Pa7ZZtRRb6+vfwe8xqC+Nt1Te
scoipNWmMlIr7Hro1GqeivCL6q12FJSQ0/LjfIohfuec2DO1a2+sy5jXwtvvVK6k
8YAb0/wfb/zNfPBvy8xWtJHuFqxOgwHxMsH7H7c3ftirY2unIc7m2ll6+4T4ArXX
QLkTTpCFLAbRZ7XXtylWEeRQVVXhuYrPfaao4kJ98KQi7U4n/6QyMA2H+F/fjOmu
40NS4kZ26RxpjaEykaSvShHx2vmPHCMabx+m+y4sIlfuaoqg+sp622gB9ZKxkJ+3
tvZEjTP/LD3OtZtgkLwEdp3UM47d9acEeit+Fc3TugRr3z0z8dNIohQjUboyZXpY
R8xD7yxPJstKRd7pMye3Vu8g3RuO0v+ecs70Ze2oexzolnRKLrCzxq6LlsHap3Gr
FV7Vfv3zbDlg2BIMvoaTo1QUSWxuSVkvRP6mNvoWCrlEzKQmsIAJ84E6+Hn8k98u
I3qOhlHHfYqmEf1Nna32NSGiV/P/yZaH9cEr7rIDPDfPgXvo5Z6AyNHJn21i4adI
y/0OSU7sVUY3t7RYcXxbEVzY743m+HL4xlOGQK/f7/D2AzgjCQg+9oQ570fVzsJv
V6VBXz9g20L2N0n0lCixTMGwrigVYomPiuLnIzq5Pfzg0IRAS6T0FyDME73f9U1D
VEWPvTgFAVoNvdJ6MmnlnGfh5QFSLbfvtBWb9XzSje8bO+u1MGTUFGAc2cnEPDTE
OYusii3CKmJVT7Ln6jBFhnwRLwYU31oJcSabKov/rbTRTD6tyTYcuLv1rcjYOgnw
+ugqNJAd/nMmZ63Hzk1ekmXasbVm6QWRq7pp4TsACj7jsy5D1tncLDmiOcILuFOf
a2pjXBjOFnysAd0HjLYAthmwEU+4ey/8Qlng3IsFVhWEDFIJF2tdZATNiT5B82LM
+A9Kt2bItSZb/AGzYFCxpluZ7AU4+tnMsSz12G3LhDh1EIJkhCLwWlSD+qaK6K83
Bxk7zkJED7v2l//RLd/VtYnMcJCPo58wPjDrFUc1xqjraTo3CefknElT0hARI4fw
c1EUrHP3K4RdcWpTqv+TOFhKhIYfQ0FSnqhlZQXF1xcMlMViDVBdooTOqmULIxvt
8pa36ZUcpwm8E1bQ42YF/6C+ptUkXhMS/ShHjusMh+ysJGqFwZfPTdr1+2fMH8yb
8K1xDIetco2OhRG6gXb2mWL9my3ErGQ1OkjhmqfRk2jocTteBGrz3hdY4JTqlUBL
q8rx806XP6tGDgOy5yLPA4LEjoA8I/fJXF3lKNuiNxPrn7E9cgMCrv9cfYmJWr1X
WJmQ8VGqYhgvDmrofe7smVo72Ka/1MC+X9E97w627OsdtoNqJnMU4TjJ0s/bXSwy
snbLyGbW+kXR1njeULdYBddFLzfK0IQkeUysnTHE5Swyf4/Lq6EhKuPWBiFeU3fC
lSmi2G3GqEykzX9+YU0DO5OSNIv3O5NjAEq7uZLUU2z6F/5Xrg8VSO2nMHPQ1AID
dD0MdxX7I0oh+mBm2oeIbEUK9kzpOI6RxomChadfRsyqTKD5ttiBfOblzXzb4CCd
Lzjwj8guksToZ9mHf/nWI21NTU3xz/4bBQv62ZLDk87nJZViM4mf40VofDE0wMQe
Bniwrp2gjAmDVqvoZbMtKoWbHfV3BAovsnBLlJYyG6sgVzg1g89xR4hxe2F3wqGF
X4/kotWrM38sGJ02YixU3wiIZGzrq9YNOERdJIU/msihzj/+pphQOVYK20k0DaEz
oQIvKT/Hu77xMwZEujIaoOVUYkvYtQTxwvHlHcIZPbw1w3O0bcGDLsHbHQiiRh7Q
ep0xVKKgOJNDhX/SGaOEY0nMPGXtzP+zZ63yBN6Pf5Wux7b9zBmIQlHqTrdE2LuV
32RpKxvre+pneMFVAF2Yy3yxUKuLSbEM2jjL+bJPOQy8k3V8iONVz8fckODg56Rx
mloXs+pMG7TYKzjSTx9iR8qvV8mJdcHswge6IKaR1G/aCYSoGh2BmcatZRN4jwdA
q+7f/PW3BgnEID8s/6i5Ausq+Vcs5kjF13EN9IkJDAJUkfIVmltqxzYErhTzWW3a
gFxANs8M/XmytQ+r5KkwHzi0ONFa5ON84X60AVQIDy7EACUFwseqPPAOk/5xqxXP
2kENymfES7tV8L7GfHGEFKBqbC0lUXKxu4wQ179BY46HNeQzjiNtSPhyX7qeJ9S7
Rzz1169xiXz8pve1+zdt5IHvBEsX9nL4Ppj7gbHXTBE3/93fts6ra/H9CgJQGDew
+6OVJ5aUG1S8nxCz31PSJVMMOArKUNuepmT5Wa+PcnTC/Oi3Y2yUv+fEyvh+Dzsf
Ms5/N/y/vqYWD8E1zLqyjMBSkETRxQSBmVJUwyBvuCWbAbxql/ghfOZbqIwbufsB
Zkpb6y6OqqOjfnhc1Igu0NwM7iFtQJjGFSQtvPZxTC9TzoA68TNSh/XquWfMc4Bg
slwIj56yTEVda4yQSHMo45idVe6OEiaLlWImN7aTJan0QuaP3kLz4Y5PzafZqdVd
foorgy96M5C5lWdjp9ljcskg5gRtNiMsZHChrIlPV2gsBGRJGk7eWSNFWJEE6LgQ
RIiZ7gnONgEopzUafTdfbL3mee0DoQHBX47HTux/xBLxmQCufCgyRORwvJYtvxHe
r3pPrsM3Pc4gGORbJ6jG85Ar/o7kuzOEffwN22SYPCI+4zCIyQ0Y7tyUKmV5oWMJ
wLuo77EtW3TnrSG+vgh+aQG5XSQt7EaFgG8ZMp21RAYbzP8VZZjVrfoev9QN/z+y
9feeP7iU3SPMZMJID9CuUN1oZKGBA7OpC689dX8V5o4mGfneyIqvdRxAvSdogQrI
j+wGudXSSMThoKaO7tyoyDt48mfynBlnoUEH+oKOUtz5IKoWDsn8YBIoBJeQ2iqf
JjNV9ff/zdsFhtuYnzkiTsz6iM5I68eBD/bXyGSFVaTO30bT6bC/FOR2q07l9WR2
JdQz/t9MAyxexCj2at/8goRjXklP90ZRe8LF3eLiEL0zzdO0vdugMx3JBH0crSGQ
CsB8kTtnhe+ASpmGdYpe491dIRbMxUhQOWTHHIkBSE023sOnJRFqZWJcFTrI+tNm
pv+PXl0mBP2TacmB2W3nMdQjh76T4mXRbmCndKs1GhVUsPcmN4Ix7dPMjv8ZwEtj
PZwRTh6yKEYiNQSsZw5pxQk7DKkWeO/OewSjzG+HTMPCp7d8XojtbYKiMv3qq7w2
FS9F7RGSA6AdeX29K1LwKivuKkv1WFS3bKf+vtVtHRNtTVjCRPbDza5uomGvr3D9
x8j+eFhPei4Ofy6t00LIjAFGSwWhEj/gzUZD2CSd/0Y3NR5QRLqouK3vqo8u+bH7
q5jIHsn+KwfqPq51BcIY9aiVzTLaS/aJL3p2eLamgAxgzC/rWhTt3pJLmsbKb9Ki
jjkIsC8s7hF5Q6/zqRv71cXC1TqSxnGJ8X8vh1T2JmBx9DU+6JxcobINRW+z+Hvy
8GkzDmVIK86tdH7XishR8W54ff8660M71De3t28DmsxQjumlWBKEDMJRd7ngV5/u
oSnJbYBMsvmU0Mtl24OZ2wl6rn+mmNQw0tlqiBphxTysGHg8LQturyYujc1s9niB
odoKxTN34s/iIKIwSi8IJLRlRCYcg7/0s8zMwG39yC63HsmJtCUAT3EuUj9b7ing
FAI4i+t31vVDnk/XaHMTlXl/Pcc4TKrfnZF5VMg4V+lXHzzESRliMPxjqBgSYrEd
bEJ1VTDKQyFzuH0V+g+Kurvg3uotGF4dF3C9TZVdeQkv6+OUfBlZu14E3MPFYWWN
z21E25kZajXO/UwEE+1cfi9VW86Tz8AZcd3iXFViBNje2HSApyP3GtHQMspVvFRJ
CSNAj2CqiWLyBAGQHF93VvQmRNuV9B2EhgbtUjdKFNjnBiTM2R4Y1VNwQhz3Kp1z
`pragma protect end_protected
