// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:00 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ENbw1H5ypYpFWhDZVOLrnMnlFf1BbzeiWeBKKeKhPtIkereXdHHhzU1hXLyksu+7
zBTB2JlrQNOpdSWsVzoi44635YtjbDsYZ4rWfnI/cz7bXkUuyeNGnvH70Rynu8W/
Ex0weyodTY+2yEzAHgFqlCXZAAdG957vg9AKLSAMTWc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20416)
qE7xocsoWmzIXc2A2ShZwMGLUmiFWaz6Y2LGQFLwxKBgZBfzfX23Utp3ZPh8OxA+
THu2yO9IWjOxuvxkdB+9moqvLX/5c9Q7mZAUXnb4WEavXpxMcDOzGGzJxhvfnVlb
7qABm6C86Uua4TmM21GygEqB6J0hg4exDbkGgWbaPmeF+BzdYnvuD0GBqxZDk0t3
uRsxNx+FP9sbQsnRcCk7StlL2OZLwRYHiTVkE9XMDQ+aZ7RnvVUeZ8dqrWLPSSEg
JEnv+ymkIrbYyjrSXdsM3KeQKnTi20snfueSQfrFqQ18MiRiAHiPxbNrnbPxFJen
/YIp457vHDD4pgGTgWXnD+LnJ7dnF8EwmYqaqoLLbKxVJrybR2Jw5sTc7z39lHLK
I5lGjwZgd5Ow3ACA5+4HsXHUc67PrOwSkiPiQUPmz6MeW4yfwaHVsGm8Rt36/Bav
ZJMYbtve/+YmrcC5T6VSJwohILeTJbjDivSjBTbTLjnrTHGAQuUUzfTf9w5aPW1x
Y6nqiyg5xaj3jarFaCYfeVZGvGVyVnsp9iiaCtgVn6X+SIohFH28oCsidSVHOMTj
bUGprVKdvU9+9SejaSHDagM9cWMTlQBOrhvcy5XYTBDPsIbz57MOcTUOx+OWr/GC
j3rg0LGiA9KgykTS9xQELvVqLlyGvj54N+jBsP7i3MoM/I74lFzqYtgDyJoyo92C
yT/ADFpLQpE0Li/UxaOOUgo8+oOSOC0Bmv+Nwq0jglOC/P4ZQ/6ajx7Ot2LGP0Ez
vsvOm6g1b4TDj6OsN+zUpuK+CQHBRB55WFP0VYPSEFufUzziajf26kMxPUaFqTj3
1sMkOxKasRRGTOrYgnZLwG5KSX3/77t5mWyFBSdPBUTQEUs0QBuJxL58m4BRpnNm
cqJriAFaOeMnPNu+pM+Xn3jei8mBn1qmG2Bxrkz4bOl3TMVbFLwvFWYmBycJr9Tn
KZqptCdwjQJYYtF2KlEBAtzSFdIlIdyBvofJV3eFvlR4cbUbi2pbQWqET/JMsEAB
UJm5l+lNswPcDEku1/menvtbUhi8L3B4cm3BJ5cQIrCDQDf68TAO4gjboacpnFfx
SHuYjBcaOLePIRUrOuwWrC6v5SEPhhw7enp/VFxc+zd4OKaszH2TBzdbPdg5TNDr
DJuJ5+TNWrb0xut1E4VUtbmlDad7fdB5MmogqlPPlA6Zc4MKJFoVr4TJ/kMSxm22
J+wClyCr6baJq3SGTK22tbAj+FJsKMgFiZdLnB+hNOXBHVMmPkA11pQAIt2aiVdX
O9mZNJIsLrExFL4vuOMIQcgmxFyiIqhR4tI9WTAt3pl0cG4+6TupXRDWfqd4IpG5
mk4j9vnRLRAslNaEWFR/g0DT+Wvfs3jAnBx0kBMEbmeMFI9hXzxtMMEaiLVKEpt4
Mkb4UVd6FAQg8P+1QBOhPALcZSCpvbGCvliqqLghLI9U1mVYq2qJr2UUD7QoI+K3
LvVMegto0K018qeoUiN9S/WZbUo9+x6WMARomVlNw89LSoXSqNPT0uHlU1Q4fSXf
k2pTCWOEAc1295Olglh+OD8p7bqg/O/TORUm5pzm5shYfBe48P20e0QFw4W4JM0m
f9U1dXskVwFAO2r4eyOmMZODh9fXExFK3tdycgG12NxO3PaNyOVHmBQOql8mdi0t
Y0h74Dxd+snD2/MInnfxBADJqysV9BczMEpprhJuHyNcFKU6rPg3ara9raPEUK69
8LXsD7jczoTW5sCxO+Ztwe/TyFH6RUTDzcOSAq6fXywp0RMkkw4jrL2Csxne8g2t
pQqRlxU1UK/j/AUrG7NFWoo1kZRzppG3yNbuO3j+FLRM6Y66FaM3RhFD+xfStn7B
GdUH6pUwf8M5nsaJP6CR6TWLnGPgwWzDjca6jVYAzIcuNkhcw2amcvqw58fVtHB/
waufLmuA0e5b3FURjko0YuYddzb1KhKlEGW1NKA/qwMS1GBnHyLY2IfA9CEMSAD/
7xC+RznOSOQMTPXB0lYHTg3nHcZuYH5YLhUXfrqHW5ogZQqdAil6hPF2aWlKXOUQ
eG5yAc3EzQ7g5TEeNeY0zAq1cQNqNmb6ZWavCWMC9p2vJSqLBc7k+8s2+8MAis/G
IlMj3gReAH4wf8tj7fjpKaDpTpySKXi4Eii4oFNyWU1KDidVglGXBclNmsZ+3ge1
drrNrc3/oWlYhYzVGIiuY36uDOqZ9c/9HkYMRC+0k66JrDNhaaiwWD5ai8iBfckK
nChl3ern6moeCuYwDwpsRKNX2Hv06BLc5WnC/ft58m1ljU1suDYpZOpysobssbGp
GKR9rM4lOP3g+plhq7C7dXzuk7O4qRE3c5ebbKWxVyY/IGJERCHg3bItocyj53kO
S/kci6i/U5q1BAy3LN6fRNy//LGezFpdd+vbUUJdq2ekx9BXN3BaaXhhvO93w2fQ
OW3YvyFAMOSGpAyy/rOhZd0KVblaQrOstsSRUR20W/d78JGL8cZ7Lc1TtDt5enLF
qIL8W5LHEconYZ9QW+/CEPjvZt+wtci+P5myOKrXLOoncrO+2rJEXMHKyMZy9dvW
ix3Gt0ppsWOUhInZJlrMyujVJiaJYsL537roZW02Nch4TtIoun5bWzDQEsZ9llfC
L/JA6bMLk2lJcxpXRj9ahpXSmvXYjxcph6i5tqFZyqKtmrmjafA7P8X11MQ+0eZF
b2qL2uZg3Ouh0+94HNY1ZGbfDz99TIOR31nnK2jIT+TS4wNTs5YBpFW+U4GxThRD
0YDVpVyqMpxtIzWqhb6lVk/OodLxGhb9QgJg3s1sffXjfH+jLDc0WLOCtqjhl5KC
rFYREr7Ch3ZcIcF+qY2Bwdt1WNhbCj3qUB0cQWetXjysbs3/2QwATunI73j6d0Cr
fBhqTXhIYSHOtf6fSQGWXLkb3vjLX0Zql1Un9VGYU2MVqWlj68mbmMrAnw/XBu26
xSCIRU6xBWPXYwJFbJD9GTV/Ofqf9fR2/6b/Qlxd1vTL3OXlnVuDHMG7ctNJA5ci
dNRGXHR596uUDhNbsc4FjeajIFRGpfko2YUuGKWngWyqjTIA5w8imT4sCTziQDZo
n7plrwYiCGOjruiUv1mvExMoDZAtcpK3nFBtZ1YAQVAbV+1FRHAo6PhRMAbzz8hk
nFjJNOqBXkD6JM+zup5bJsfEr9v+gFyQHnsWawF4MDTstO/Rsb7temualhCDAxi2
HWNp9NUd0/MGlH73IiNKipZ/eh8GiTte/APedb+9LA51PURXosfUFJSunevCUzvI
mKUiz7X9qG+e0+uTJChifrHStbYs0hl5wLlx7UpNnmyff/Ccb5Xzd87L9RehIboQ
K8Ah6IBtmPhaeJGT8NghfFguSzZA0xvZXUamPM8AZoySOB9OizON0RuU7P0n1+w3
Dzd0xgO3ABAmaputX3fWsfrj13HueFpNk2ub4aq2yCn9aoOUM8FmTwUBdtzq12Sn
5wdmfDQJywVayinJ1GlwHDta3UTZMmUI3M3ozyk/R8k46762B2E8Drs1jtDLfP2m
P3OvAGp2NeB+5zHT0AI1Mxot2/USE1LOB+pGDp7uPuogXXCExpFGSB7LNCIH9Z0m
kNVT4AMuBoXTWcQBnqt5QqIos3HzseI3WuatMyf/LfMeusaUHapc18oGSLE3xzzC
3BtzhWq85UOFktk43LuYxGOF2WKPZDyUmFb02SY+qKPQfVSdZrJvBHLVOCYK4Hno
dL8ZZ8qB4xS1TVIVNs7rV4av/Xy/pH2CwW1V+hPaGeLboEMG1BAxd0Ii7YoTmK9w
bszuwNAsO9hQ2EbUX8NiTQIspoc/55ZVgedkmSe8YkoZwUcB2p023YLO6WntUooy
rz8hTdktxI9D5qebQnsfTguIwgVN21Q2RfKhYf/Lkky7NOLk4qiBpeaZHdI9rDyA
iuptw0sEwqF+5RaroDYmwpVPUL3bBIZo9Kk9MzNVnUMzkpYdDqeV2RqwW5E5o2/A
GyfoQeOniBuh0JjhrtN9+mFzx2wy0nALZouJatszOIXHkPY9FVzl06EIsoFYbBY2
i4UWqTMuD6o5Z2IqICxMyLU1no9578Jh0UGMOzN4T/FcLPdt5BFszyiZ3eMW6XQ3
aFCJaLmnYhf+VP64in37SKs+rqEjq20rgehVKdAD9sONGCABy2bJnf2uNaPqmXQD
XsFKzL5oshVZGvrdQL3JmeE/kWq6MON6305x5Z1kKZWVf+J4mQ0rDEbRLtQW0jgk
KqSFSIzTsbqcnUqtC0FnLw/rUrMXhfn8SiaSjU0jYqhXyckWaAgoX6i2Om00hp26
h5DRlAUXkPC7iO/Knj1pgFJuKyAO7zgZCNAKjR1Vrr67IGuB7l4YJNf4J2PHfEDd
kHwl8oJGMxnQcKiE8Qb40v9Oi4Ygi9yqLLC2tRzmakcmH265BMXnpQpBp5ZjNtFi
TETfdI89BnaV00Fc7BpER1mXSsTfpxk0pmRK6Wy93sBve62PtLervVdOUEvy8tb4
yoIiYk8yWGcZMFYGRWX2b3vl57VbmilEtf+3p/Khs8U9U9ahpY4zcl+LNja/skAn
5MnlruTl4FbhGGj1A6csGsoylg8QDE2k1MIxOkbSr9rGAZ5m9Ie5khSxYPrvGiA1
YzGCbSHgQHEF33dvC2uH7sPMblnjBymG0O6eMxP4/0JAr/BpFDzN6mYePeAJdN1N
hv56sSR2TO8XWDXuSrpUf0Cd9ZXHQQ+Od9GKx6LaQ5e4vMzSTdVBvgYrz7fLDfhM
fAK9BngVgB+J/6Ua0ty9r3BKEV0xg20BjffAhsV5BqRU8LZpYxT7DPcFx2DKSlVr
zElIY0joHY3ob8AgHL3UvfLF6i01cmHmSxtawf0ibFJIfh4UwBJpNGmpnLMqplIj
GAeV5+sRJP3arUOuXu3E6964u9HNYxMxJC5wcR0w0Y82EczSzQXX7l5KBjVNooUN
iwzKfsKAOSk4pc/NCiNwsrknDu+XsoxoFBP80nSlhl638BoFp4w/jmaIWgAKwlv9
mYfDKHPYw+GCTWgeFnoaTX1FijAnBBuk3n6DHdpEzSsir2Nolw48tyf48aPYcFsQ
NOMhuAF4OqqqjhGxeKmjWhvkqk3Vs4vYLApWc5jqkQmWFtKvtBE8Kr9/O2lTO5oU
ftu63dhe942k/kSo7jKkhjgtk8OIsbsX9RRAVYigRjOhpK/gub7TKuCGWXIwWuwq
LEIk0r1BT0JjheV/Z4Ymfmd92jHxnG3zl3r1ddw9aEYPOLWI8QHLqdQXhsVuVumI
qxKFUx4f404lK/9kTF3RMCch39wtWXPEqwLw7ICDyxFkL3G4E0TinNQwlH9ojcNC
REpXe06oKy8MzBGFwWGUivu7M1Kq3nGBEzXtIX0V4tuQRC+E4rYoZDP60f2WmGYH
agDAnrjBCqNAMY1dtwRISgIECcawICskmJunJXu1+MnejduUK5KoQE/6A6CgXPMg
EbRmG04cWYxs14CN57YxkO6F2eq7c7YSkA3tmDecLorXxWUtrt5cnkowUZ92ajy4
+tod/K6Cbdc8E7WRz2hVcC2gmyz5w1p8lHAb9cEv/3/wTWDIB05nE/nm8il9GktI
0McEyoRfFUUWsdR5rxfFoNSu6T/Y+bCCDD7R7164jU3/hN+N+tnn2z7wuE+Gllij
d+tFy7WC8eOCjgDJwcykpCNyWePQsOOIcaf5XQyvWaGOf5S5IwNFuqMw8Y3mkljQ
m3c8qDrOYudKZFudMZ/7MO4Hoy3h/8pQg/csqqyIBIcDAVB+TLZFs+BgFRVtsWyU
zuukIRJosphB8V9VkuD754wzqcZXnojujg+bG23FgDF9skVUHEu8b0vSJ1EMN7Eg
g+O0mIAydHeBBtlihu3tTHTFFLXbg/DOzJFKvVDYPBSgzcouAwJxXqieyuJKzoHO
nhMvVbxwhzRBsIuswX17JCA+Lh3zkYxzRtNByU73TqO1V4GsZ7vy7sAW5B9TVReR
72JNm8YIXbCeQ5rJ1jiH9uJ3ELnGCrUP1yFGkfhA/ANFh5wosnbSvOhjl5FM/J52
+LQ/ICVs6B31VAfJgQ+cd9K1ndFnohnDoi4pZPe7Xb56rcbw/Z5epOB21PEkxGp4
8r06z1nQRLNtk8oNOn3T3luZWajpPA4S5AjBY1eyBfTTvnHBvOWBwytGovx+l7jn
oTNZI2B1Lj53J8Q0DNyX1U/Fb490naW8SBkpoBOBAdLdAnuI9jkcAoUy5+QZLCQr
Dq0Yj4ZvtspDMDLsyAaaE9Qge2X7dOctOeEOQh5NUq6t5O1DxZRRd7TDAkUIIDM8
LQIWNvMAoyg2gCQL3IF+kSkBLEsBylqOo7cUxFzMbJ7L1h5fnqSwgOB248nLAP0e
hGgTjn+Se9XJER7ubjXS4HWwN6guVIkCNxJh9byk23HFEP9fcAm6+iosABNJqnnl
I+2TGa9lbVUD/WQlk0ZTsC1LtD7eWNkLW+l2G1LCoGlrF80orSkK6JjhHRDdM/J0
O2ByWP03RVbtmq6ZpGrON3KsRMmEUoygdQyGPdXiyQEZNKegfzomURY0BXkVvmRf
MeBijomrO60B6A2aVwzR3gWfSEmHJI61VUjzmQIrq42rsThLQhc5RW2+GbhlbX6P
ERgeptFFxrPfs36BUVnnBPckksH/Nu4vUh8c3yvqPSmfkZK+Pk+MQQ3eB0bLivTT
D5BEXMEMcB2l23XbFYE+pzGJ8TPfE/idgGUQoGhdy4sb50p8xQnDrjyuzi4pPWIi
HV5bTWyCGxAoYV7ROl3g4sa2GQmAgGmCzRuYHriRvy5+8mweVZAJR4ppzGHrw6Bk
e2yz+jYy+txc7zCJTS2xnX9EFmK0W8RNk1pXYHXzaZjhxnZQKvVO4TB2mHg4fEej
FBbShjgdSUre0TboaMwjKubXLs2eaRsKFITvJg260A/U9d+TjMirmzY/KyKr+ZFW
sHr4MFU39Q34JCfuiGSi7zBeT4J/Jf2tWvzTLrwzbdOiDg//1EzO9K1GVVvMPOd/
+i/deUnSGoPFpwAXmMHgKxIsthvnvvqUjsoYlo8I4T4NiURVrx9y0GojVJwjiQXR
uCbLRiYxXmnf7PArpBKwUm5Lc2s0L82fBXETJgeQE9k9U0S5xmFBRoLrStAUbRY1
Ua4PbVG4ayhIYidDnOCzsyF1rIJHMTxsQV30y3MmTVot2mggc7zLOj+yrwQeBDGk
Bptp9xFtb6iujQRFzzvx+mOSWyH9q5tVkblMMs73T+IXNFwO8+7u/+OUVLi8ACir
2QgCcPRcnZ62i1Qw30UzKycqGF6jkjcuPPaMUg90mltTE8EbgIQRKHzbfGelCSDL
+ZQv8hhemfg0lHp16HW9LOQUqkNGm/M0UmEUF0C8twyqbZztLSQpZhk+VdbIKMiw
pj0d5wbh8wUlEWA9P3y0Bgd519w1KtDwrILsMUXXY8Ady0HEsZXh9jAn1HNmO9sy
a95vFqm2I28zch/zWwk9Han6DvaBQVAQ46TF+3zx2Pfcht/OPsJ2SAFl6rXcHRge
L1E4B+pFWeyFcCRQeaVtgfeKX0vRWPUY3u9iqyte1es1sTYixC8tvF7haARAuAND
SmcxkbnTqVqJ5zoVeCTvGo7ylL9PYjbxdVNP1ZcIpaDeZ8DGpik9glVAbKP7c7mB
UMZb22SVMLChU75jO6f50UUejLqBTRdg/39fdpSERGxis543iW5LdFFvVkGIoBLb
pYP7l9H9juzKTmvYW5SyvBecFZpwDVxT9flOx2qMQwjGDtyk79CmGdoKayBehIus
tq6OQ+9CetptTkBXzRz90GXvocTEa7688WRvXwDj3ihJ18kTYuVcw4dInq/jPsoe
p6Q76DbBKyZEwdokBiTwIngz/sKh8ThFrK+/joM5SzJv4SjDFz+2QFyGkwl8/qgr
wiNWQm9n2iCuAd8reMPdLBjCzwzqAkxKA8Rrh35yfihnudRaL7ozWqb06IWX9emb
NKMkQciG2hO1TTq3KBnV2Wk1ffKDAAW7wV8hUyqGWPQidVN93i+gX2scNAFl/sia
oXQJgiiisB2J53SS0cwnuOwZ+jBK5aRoPr38DJo13cqPGhSpoR+ONRqHgBOI5OV8
LKhMJ7fGirWZCTDBvPq++sOmEl7m3g1Y5Qk1msU7CVpl8m0tnl8DXK2bftClkTad
opumNwXDQ2qxu1DkP4QbG0cvpzkHObuPWei9NXRpTC3MIBaIRtlWyrim1XMhVMHW
S4qLbIHZd96KecRGiozGXv45aV1MMqE95Vjmh6yggY5kJl5p2XpmSKgcdXVUM4M5
KfH8RIINKrWmLuVCEwf4fk5uRBwjL5GdcPv2DgNW1TYER/T+g0WDMBIw9NyvwCXQ
Wvm5WJ3y2NPJmYcz8K6YOaUzJ4c6F5H6Kr1agXBXkQZPQSkErnvnrOWawg/517cf
p7LHXju+tNnc3LMuhONlgULxOpvUCI3PxQr3Q0zywI7oxIKU64EECoRrGr5ASb65
831E2+2U99LfCaIjiztbESqXGI1xqKfIskij2ZTckI95/tUrC8eLk+dKEYYpeb0e
Q1h0TkY5pkLF+Y4V/ELJwAS4kCmr/gbN+ej0q2Bs0m6tWSVFQ7Q36wnM1i5Mu31E
vAUpLuPymZI0JZOAVFQZA8uugBOMTw8b1PPcyF03eCPqRgffQtwdTFjDI548UXK0
rrS5olahS7HMxlDTcVciyOj5ewLEOTh/5Xz9QsHsESaapaNgtGkKfqJVYHfI9Lmk
bLgnE+YSTmddpW89Kz48BM31A2hOiC4FzZaOfopyDBW3/OPyMUiRBseV0RBwxaOS
LqyTgPlznV3Zp2a8c3lSO2VDT7MKS/HPMLK/PJZiDAUSJevbwt/1ZGA5QyOafofo
2tJyoNw1AFYMq5f1akBmD2KlhSQUoxmV9XFqxfCnCsM8GqkYmDUhKnzvYSWd8uSu
7o/M961Sn+BbYTtw9j2QUxibiCiH3wrOZud3CZem35jmMpTc9OOqKo/efejvV0hh
nfJEBwT1+QSSIWeuWHhy4nowqhFMCkT5vO9CgXr9QoecHO50z2itAXvkPIwlwOCf
/PfU2BumRs97bZGN0HXAUkHZ12POzQGJSl1tZU4EPW38wwC7cZbt5cdnj9m76gzS
fYqU3fbedhQETQq7NJvbx3JydzYFxfFCK1786FWSo/YTJLFuN1lTsQ+cD6Vg22T2
9LqJ8hMabNGM9Yc7d/bRLJyjLiRiGrNqU23e3ULJbnqut7lIjnuofsxZv5wZ13r+
KTMVNLO4B1gFnidXRiFYIyNvcO5MEoD92oPQjBmG3UOQJ20T4QOL1Ylobw1cjaRR
EB8wxQMjf5OCT/xQyxrx+e5WLGZJnkHg18GtGW2ioNP25zEfFNSA32px8RdKm9vg
2SQTxMAVPtfRlgZr5c5czWq3rhRe5wd+C5++vMm+h9TO+do2mTcZHYGGt3L0x+cu
sBOQteWjjiuEcb0L8vAeUcZzebvwqtKpgXgUQagD/Y22SeJzlrK7/uHStWVpw6ib
LHc/i7G6W4b+dnsh3hIZb3/6CzfHtRLaGWBRQX52s/pzJrq2iQkksU1bsEBK7ele
vb7RDnzY33Ct4I07+wwVjrdW8yCZfgVeZ1NUoRuoosXmRkuie7fGEx/edD5iVvih
56Z2vp1HOjA+wU4OXxlcGjN0E0wHXl73xzlVgC8YZiugMJv2wf0vAfqMB5iKOsW7
wdUJZvtJigUgpQ5Vc0TYPjeK5VKwW0O8249e0VBpx9GkRXExnmdNaxvldeWnyinZ
u370BNFTvrY/oPXXwh35IGDJVn3O7pfST+J4JJ3BVfax24AKVFyfMNKmBBt6Brr/
qg6rhRj7YRph4/8DJ9QYbl7HLVjwGJkd2vi7sfdHvrqDyayAVJ3ig8/NpS+ZsFQF
QCAilcoVdl/v+Az405D/t4fmIby0oQqfeVV/Pm/Ih4ka60IPP4AG5CfTAiax7yXQ
8ZKhBPRb0sC+CG1glT2e8HEeuQxV6c6EUHYCtuEJUDzN9Lcl+NOt1VzR3MdfOpus
IAEpO2HUfb7GTPzCJardqK5MMMb1mSdMvmEUQ4+pEwrJsbeQIWL7+0ysGMxLs1S0
7iO7p/SDIleOhbXtpnColkNlIPIiU/Hc4KboIF5wZ3MG0UNaCPEms8UtbJEELUCu
ZPBgo5wpKEzF78tgttcL1lXYlRSQEP1f6ps9YXyEHX3/uk0c+5i8nXLFQ6ixKBGP
hBJOB0ienQyUO4jnqZhndkHwOLCaFBYvZPeEaVL+ysQHWBRfpVJhOFERUEE1rTwd
U9/o+guj9cjB/i60kT+w3TGEfMHigZ9l29BbfB3RcvwmtnnmfaNtTwqdKOVutJ8R
jzsJ66J4x9TG8ydd4g3svnkv0z2X/J947b78OPCsK1zOY+TSfOUrY1wnAMgsffkI
5TXgH/rsBD5z1YoSFU0o2ckSl4HlcztggewjM2IF4adbj+9ySf6uXngH1v9rYjJN
P6oVcFLLPfUVLmVxBTBgRXXVoxOuHHFmp0PrFPBnl6JEP2SIWW207Dd+kC1VSaUi
585VkdC1Yo7CPRHb1ra8EuHn4K1gUOBsdLsHkOPZAwQ7sw5XV7ByhKaxwetpefN7
agpppWD+RHOTPa0w8u8nBl19hFdNw5yiTp85v6JW3Qvs+gqSjuHCuGwdb+XDIYJA
HHhm5oSjY/x+k+oLoYtpcVuhMifXbYRXMeLGJNiJoZwf5ltnfmevhRmlHKdDkty0
+haNWgfToNV5+K/VLrvGW8xqeNwYo+OYkwdclyPJdRo2WzBO19xL2PhKLY4aRaaY
gc7Ds8Ej7unnu8Og8IyQ8wcpwf6RiUxQAd+2tHcz0Pq7lhP+Mioi38+81GRhwCMb
Lu3PavoKtG84ku339cVXXL8X5Pos9NICAZfPDP20IN/QGxlePIz9ZhGbk6calKnz
Yw2CyTpn9xEnaGSVvk5kN5FHWIU22uGkTCidZGTEwCDS24Ho6JFjIR9NFDOVktNV
ExgR0y3DBVVpJl5YxYnPiSaUbz8GQn95epjKJf8CWGc0gl3Gv2+W5jaN+7kw6wXm
bkjngSPk5y7PH9xzRrEIY0olWFMNUzJG8l8RQAaOky0zh72ZbeL8/sYHomKjnbS3
2pbZ2P3XNC5vtQkgl/HfuJh/iD2K4GuJmoto3b6KAROi+I1APt3izIkKwAqqZn/8
ioBfQjryqA/pUKypSLC6dtrVE8z+Ht8n9P5ZSVna+NikwPkqrejal+4lx/bk47GU
oNEUWkncTgj1MeCjnORJWgIijoYWsDOmN9LAqZGzftukxpN4z0vKc8woSjhRQTKa
cG2ht6nJ9HrR6wGne9m90Pz56+4DokHyK2IEn/RX1IU1z4WSLVH1AJMoyphycHe4
zt5h/3mSvBOA8l9vnaZ9tEAQqxhjMbT8ndWMJSb5C6CdFTXHd3yq8lfZEx2W9j0I
nE2PnIPwindOpxSTYy9sw3Qclr3DC4+BUhUMlZF+Wxcp1Zti6Yf4wLe8+qC1bK9y
qon81sQ48SRbC0zbcr0levGe0hhtV9+b2xhpTT+3UuRP9XM39ujK36sV++XBXYaO
Y1i20DWjmPV71fH+4n7Lvqtujk7NWKvMwz/m7diAg9H+gXkFrKNHBeVzrjjC14Ok
se7YsiW2sFoUHxOCcu1DSLColDNobjm1MoOHNxUO9Us4HNef6kyyzibaSL8pzBCB
cIjrazVszeOeBynhFWSIvnag3WXnTeVCpMF4af2tivVHQ15CkR28dMaM42btJNK+
Tw0XmbQzM7nYxN60G6ElS4+udmA4stM7HmeAZci3g2uhWk7gO1OfLeTp3dTFfdYM
4/4mNXcBWUPNcj9rJs4obRG5Jc27gbnrbtGf/aSw6dWMQr4d0g0BHT1OyU3oNfY8
fJ1PeGqQQG50BoNbGq0RFrIpztoQU6ZzaI4UOD4NsbYfOcW62jdlLt/T2D5enEAe
xc/n0fxpighr4Of2rCPXtjGV4VFLrBowQHvKAFxllTQfdezonzb/kVXNsk5sYPfq
eFfosjuY1dP9Xxu2D2hV4bL7k0f7VZ3I56I97oIkWy6pqY2YaTH8rM0MRF3tJUjT
qaED3pgWActpdCWGNsDCjU+6OQ+gn0R3lj21Rh7H2K71/uQdti3/Qax7BlHLnpjb
J2+IG8W716aH54BK26kJ7h1E4Tw316f4u5DSfBLjNPppENhoXJKsnlUojdaayW5E
VGJWrgZtOF8xTBjuCxgKAIF8Sp2clu0mONZIoaqFdzkZSuoqI9Bwd31srs+5SWpr
RiIWeD9z24t7RXE6+RPC47MDpvjeBUdvssxv+4rj2fpwCdYNUyGj4NXXC4dmje1J
9sCqtC2EXkNK9wch7wVmyJy8BVqLVVCM7PcKL2TbtDwZMZQ2SE9wuBj5UFFocpmv
oPhLWaFvgCwDX2jBG16CpZUA+yuAiG75nXYf+OkgHtPOtDLwJltTYkH1Y1DwLbW9
YqzaATP4mtP2qlLTRb6IINcwepioSHh7h0ivbFm0V6cD7+vw/EYe0qOD0V4qxjbQ
SVTPiPqo74uiWKOiLEwuXOGFFsx6C9LGJ7RkCN5PyZSEchZyoKHYkDZ8Z5w3UykU
QobXSPzEye8GKm0XD6T1jIChcEt2cojYwoEVoH8lFF6kVTnxBDRuS9K+8YSaOe8o
7miKuPXwQ2euDgNstjF+nCWyIkQObxQ9lLMadbWA4/1ztsUdHcYbn2EtNPoRYlk5
4Mch+uNZPTI8NDYbuIu2/ty6QZj+VU6oXlR3mwNLiEIqOLHq2fKp88DGlO4ehfWv
IOGT3mbEWZr/7tA/DUPtkI0qvEawCQ4VHIJNnitRNIo4IPbJJjZz3BIThsH1tVWK
Mr6lg2AbvbKu0D3X7nl1+Lw3dv3kLAYj8KZTSlrZm89Ol1hohDbbLgyiUO9lFx4X
0+KxmgNrv7X/bpZk/Exbj9FrC7IMUh1/9iLFK1PxVv+9/pCzhelA16hZf6PzbTKh
v0i407EFmYx7WBAtP2KVfCnVl8Aw2o16o6LDF0IdL2KSKYNy7bq7vjdrl95TCZR2
QVYb9sqWtKKXuxYoMEIeiMw+bZPDUSp9xron+mM+C4CNb5sBKqi3i6OPnMPQg0jR
agvtPaVVV5JTiiTcrQxkZQwGM5jGY3x2F9jgu/mAba4cT2exi82W0dL7rzJvldSL
v7alVMkPaulQOTzYc84MBWZ6KFsBQBwUWTvy1oK9NBcvykoY3KKIpxtX7auvG/Km
MVq1b0vnlCM7eFuViFFuY8oIOUkHH7NfDF6Y/prGHuvggCieoWAcQnwodtbYMFLs
5lLClVrr00tMy4soMwddT5nLFpGvIIIvX59EIpbmXazHmVl6i48pv9CCTEE7AHGy
kUG/oIPSGyIDjgDdrTjQJNhwRYoFm4373y/eNjbFJba1o9m6b8cHD5jb6caTKuIG
3nlCqwrkagNRD76XGlyM82/kke9MiY0kSRa7EJnwt5zxLT4pVs8pOzN7wVO7hrx3
ZLjtnTtfNjDvucrQT+OuY/hiYIU75o5ejAiVtbwCF8fDMiUC3q16KqRNgzEdfH4M
sQE+qgUbjFGLZoI2Um3H7N5ff07SFe18sokuq2a2LnzTNz7f4pDIWXdBwVhFpQt6
CA2HpVUmmG/I9wGCbfVuwIQzKWhTmKd/40GIex9OR6ZIFXdtX/oi9TEz49AtQoAA
xqTGNhA6f8s17ZqKEUuiBIExGhcRhRvatq4e07DYB3YoqpZ+mW5Ay3f/oBf8juy3
R6VEZGtQEtwMPaKs+P0SP9f+CmaVPAcJjYcAAKbwigXqJ02xh/PHwRRoGZQQD7mm
J34KmIveII56Tiv5+EBUBpyHn4lmJf5i5psBi8eHgjf2Kf4Oq3Ql/+lh9YsvDtSp
iBinyROe+SOpge8CrffHgBDmKzmDKiHehZGv4c3PfO6thGwWRe9zL/Ndi+mmLWvt
fo3Mqnn0e/9SlkLq+WkXtVv2kncfYN+a8Lje/UCzbkZdxSA9dH6jvDdcnl4yTtE4
4p3iUvqJSefpgLimu0wEVTOzEUb8GV4cyrsK9+zFqBTB+jXIakLxjyho+XNGJ+qG
qwC19kkxiD1rBHw1Va7yZYZxz5KfcixIQAsdLkZBn5FyoE5MZF2IMyApf2oD9rBe
O81qDAGqn+me7IWkk8Kd95pUOn5HkxO34kq0TSkCsf5/oyZhk3mZttG70PkspYSj
ToqXPi4+cI8zRZsnJnX3kQfNBlCcs3jGRz/fxo2+WQYAaZNRPtJg/eyFO7QJGi1K
WFtApq+0udMWZ/E7qw2Z4s+tCndQHNwX97tSY6A0Tn2J5l0UHzJCp5Jr+3aJIGwJ
qqPXT9x/7KDyYQ7jnpBEnKlEs9xBPqOt+9CkcCGY1QTLK22XceCMr8IN9OROV5q/
q8IQm4GyQiUEGiCuE+HR/UXDeLtkZLe2lqgPTvlP90tiy1M4sLAObUdJ9TU/0WF/
B8CfMZcTXBZ09qjRL47cZTM4xMlB1IdV2dPbOT9WBRNbRlRLkHysTgMaE2kmYN/Q
8ba87ImLu0ASsiyGxnTKSSBtSdnquTbOgOvnkoV5W6otO3ZgxNlXCeopMJaabSuk
L6ZmPjRUbEiiC5WioMZHeCJt818OiXVDEmbsanm+jNlmDxud9FKThk67vE7Mftvt
yrPFFpCD3KlpHRHEzdSR4g+U10s04ycPOPhV0MFDtLP4GRk3H1veui8HEDXF/4iR
jSdwKClIDDEdTCxPOIj8maIRtQs1H+8zawT55sjHbQW0VjPXT5GNdC8lB3AIswBi
TWVQlAMige7Ov1H86jv0rRCQukus9oxRm8+/RpP5TdGemw8h4IzLUVQbsqV0MLNz
oGYmGzYvvCHrZXDn8GjhSWB1NbJ4l3td+XwXjWAFfs/eUiXQZDVZkC7+4gsM18zf
aX8z7BmmTYMoHVBImHmzpNtasNgh3nJfBpmMYWSdViy0NqP+4eR4seAD0h73maIT
eGZpuorEjv9Ep0nPnDoD1l2x/GCfmgZQQvXLqe2Wf2aRlH3wSp4Zn2zDliE62yRK
tuf6vzLhxfLemzXyIYiF1/gmaRlJvPaGTEvD8dK36CFaYS65YFQ3FzZpbu1HdLWU
d/Be2uh+a4FGx4QCwHSZXA2XIo4U2bLV8eZP0ipkn0Sv1giZYDpYfCavxOamdkRY
9sD5oBSfTvbkB0lc448NELLVIJCgFLMfxMFL2H8efx4RLau+hovic2a3fY1lVtW9
giqFz6rXBnLQ6dRUIY0kKhc2Tz2ONmG03sbuLw6Zvq1+OMwOoC9eCdS0ftiMDZ4q
MwRJX7wSyTJ82fFyUwKQu6Qqf2sSrsvk52WMqV0XlcfdSnp4dqtyQHE2rlWKSh4F
zUuQl/7aibLMS3B0TFMMfQNo1f2FluT5vw6ukc+f/zC4wgV/Y88WIDcwbtEBQToQ
LbZMimNFctkoc2MwpHj/v9PweK+Eves4bXfI7a1UsqKBd1ruRN5MhU2JfePTB7en
YYTBaFtKzTLSGOyYD3SvRcP2qLRDS5mJfc5mVPf+kac0jKr3b512iZV7PK++nuOq
5/tBr8Y9IaVPKVIXDZTmKWh2HIzvrsw5f8eNYslNY12T+thcrWIYLEPJGuysgY4K
mXIUX75kqVS4WodU9gEY3EYDGzW4FZrVCTKrvJ/sHFMYIScE+bEsZ6NPstQYIy7Y
6Z9Drejau2q4Q/as2xSwW3jH+HwxoxhXt4gtiXL5YlQaYMoD+i+uaUpEIDImW9b4
wcjAkMRCLR8RtKq8jlFdy7Kkr9D82YWUmnXzbVx9r3DlYeClHeZr6xSjHZRKdc4Q
omOQE6qNspS/oLfJipDWw98WO19a0+F73eYpb857Pxa4P4cnOCTkllokMoSKbDxY
c+vZnnYEJNtNFM0NTCTo6dswM+zz+uSs9lT/KZtfWNCJtja3nZcrofSNkl/PoBIl
NrL+d6a9kMOsssAqDCWfUuw/H5uDEwW6RtYrpe9ktX/QWT/WZwe6EsIQlSqAw0f+
inYf4QFNKSsyTf4s0kU1CdlNwM36PtYtlfkcDYUh+LoT2b85g2SOdau8AIM4PnDB
+urznMe553CyCZbxxmUoh84fxRAczS4epO1Ps8prV0lJLjV3oo8C6soGBzOIo/FJ
DD+ACQtPi0fCUiHSjuYbLcdelF6t+eSkd7pTHtqoWXgrxWGAQO2aJPTL70YBKS2b
X73581rQ//cCMfeA6Mb85vEkNtuD2T1u/UBu+M9E32GRfcJt7GXQoPBADZj/z3O8
BAZMoU0/4wfn3q0RswI3vMA4ynnIQR/7Z5o8Cl5wW54cQfDoGTH0YTgzkKmAwoxL
pfwllEGIb4gs0FmXwmdyR+qqp4Wbn2gmdebFGo9coQwiu+J1kwldeEL/iRi7UZeO
qc3mjEQ9aF9ncNR7SASk92TCCmBa5LncCzgNsn6jk8WjS+nOTGcCBfFWK9YNHW03
NuRpJ6h1ZmWy0rt9SWPLdwOIwEtP0PxeCpxFnrH5RpdkxopWR8A7ggIB7XNIAFKT
3ZWn78gAH6lWpyxRNfZms+VVVzuKZLSx2aBh8yufvg0UcjZlnfwmCkmTNOZloebj
tJVZzWoSfHxwz5TisCjb8Ty01vgFnY7NbaSuQ3k0p4h+eEvFwWs/Gy2gwH6jWkCh
ETaEvEEtcVSTEJXkIXcryK4deezGuzT7l4KBf7tPpsrQdJpnt3do3H819uGnT7G1
r+kaMSlpBNAKn8PreUGUUzzWwX95Hxz8LUA8x/AOSHTBU2N63wrTCE++VUo1XPy5
MCdgRs9ok7NT9Dtauw0Y9Wn+ZCGCxnmN4xBwq+t39DFJluK6gFESRDaMI8vPuzwz
VQBjN+S1J3oX/TAr4UbnDmS3nwYvwpM27NBgIOjl+I5ubfS87YnSYJMSjB5d5JKg
IaoGdmzhYd0694Etl7YvX3VhPemYdJO0d6ksLBVE7hR6J/w2hc5uw4JG/l5yf8mY
URGSe6QTb5NW86VXAqpCN2aOZdJ+rHgJyP6vgYKnAgSkTMLjD9p3wA8YIWxjCSIT
pY1MXWS/rnVPxNVZ5gtbDW0BwHzGcPHVWBLwL6nbBQ7Z6+j/CXHxZbnm1zwozrn0
OLvNZ/mXCP/PlPyRmB5bsmuncTxR/w1xFwfSOwWTu6NRzlocMOWLMOcHgmDMM9mh
i4l+UGS8J6PX+l6+H56r+sQyn0i5Gf8hOXTrp3WPpiZDmK1idcsNTrtrhXhvPdG5
u2H0M3APJf3g+RM6KjUXl95yoImp5VwdXJ8gYKI94/8i3/795zEYiHmVkFymalmR
y2eZbY+mQCILpE1w3q923qCl7rJQLRE59JuQifSXIkzkRxdfCn23bIdWG7QMTrfL
Or60zzSXr2nUs82u3cjZUue8ny0Iu1xFusTpui66Eu7r4fyUrqnDibJ6ica5eHWq
xTxe9wl0Qi7onlsQrYTN5OBv7nega2dis1abNwewVc06X1ID/yrNMo8fCLbE7OmF
aVogWB5Xt6WFU8kYg9SOfBZC44Ce+BIKq0Ca6GshOhDjOzMN2mAjEaEALz2vakL8
aRQGqP+pdl8qpsEWM/LOvFdlfMsGeebkRCV613M717lDy3+YjCTMXI7eH4e5kYVp
6CJMIglQIgNfHC6sYL+BfTBMC2xUr6KqjqcLAp3P7bGM3KiSDEvgwU3R7ka1DoYb
4tEHqrUvGr2COxsOwjOMWj9LhJgyIzv7lcUhhy2Hb47n4tEuz0CpJmtsOoeJH1Qs
aGBtS+Ao3hnzaJMoF224c/1SmTSoksRjeuhHYCwZexgPiCrS/bpmmFlDtZ9xoj+V
woaO4/VKSl00YiN5MoT6N0uuGB6fVDeg3lnqxRnHJsGtCPax5itIUqI4RLmcDInH
aAJ03MZM3JKGWmkFk7UVYFlJPCqg52K05qBBFggNfA8gw+Wap7gtoZlemKFKb8n2
0CsASEaVj7gd6ic01Eji1+L4ega6yHlgtfC0AKV31d6YNVpGcjFCnQ38vwZd2EIb
3IJUdNbpSntCP95X6So/vYO55YAN9U+KvIBAoDZcXEZ3Mo4sldc79XCvnQ9UZNAs
8y39ogoveeuX7/SklFKH1VN82HWuWk6P7Ke+qHiRJKrI0MqaykfRs2DiNtqiQKZE
rEdiPP+0DpUqF9569fLDOtsnbNIyOUWcU6MhFDeXpF5d983HUqys1he/Q9ZLvmdW
hUKtc4W5I7dGKMIogO8oT9z7u4smnQ3GfSWSUO9Gw2H/98EPKpsSBdCb5Q/wXykq
59jdoHFElfAoTvkWil88+AT4+volgM6kV6NS0FtrEn55zaDHpRE85TYtqbgVH2zg
Pb0ua+f8sF/jUN81twqJY0jOn/vJeuMHUMTKbYs+s81dwt+9E0YdcuLmGQH+Si67
cC2wQzi16UGkyT9XRhBnHBohGHm8gWFrh71h8jRzR2GyfP9p4RsxRIHtKG2f6FrA
Opd48DXZUydMAAD7l25fYBH2WC6BSPtyVmD7cyq4bqbpUVrfvZDMmJwM6RHe8Njx
j2JbkWapD9zHjrxxMi5GM84O0yDXL9T1OZVGg58N9DdLbNYLWKdlBZUT9TSzFlWk
YPGmylYLY1M0vVs2ppfacoV7BfxXe+Rx/DXjhQr5DzwOksEkFyykuPyNjHImhRnq
af3MxZf0uIJ2r9fhGbpsSbm/VfugfxtS2DNiPrqjBIP1HpOXu/lxixCWGzgefbDq
y42J+mi221T3LToseQHJEApYGY8PFVs+3pA+DMWZeM2grfaFpaIoTy5Ge+NaJrUz
jH2LhcpbghL5I58j1/f2gSQecM5RYT8HtdFKpVDoTj1+ghbhzrVZ5Pop/kgsEaw4
yCyC5eTvYFNfbVEG8f7JwbW1AM/rUFaVE5FyKo7Nwp85DJ4YPH/6wfJTy8xVBsl9
jpQ3GyyGrAP5+rKBB+2N6XDUQCZ1jm2BAi4ERMWbZYi9SfPN7Xcu9/EFBooFdLh5
OdkqVr9P5CLQJ3UtlEueQxHanQAyWp+onrqIchvknayRSHgCQl7QoU1HU5EeodGD
p1ANDFO8aF+64iAP+meAJch9kUj3PKsKuABmj7oPOc1+ya/8h4sjxsoFO54yCqTy
IpZXaxtAfjgHwqaGaQeml1YLvJ8fctftrH+JjuODRaJri22mBNy0Qffj5apVbAkG
CDX3F6ENxv/lTiLwL6LvkQVoHBFSNm836yCce/YyOVCX55ydDQOyfEszWUuRN9NM
IcEe/rifbPvBJs1jyn6YqrVBOjGtx1OzvHtQMICQI+PRPbyYnGPpEwvGdGX4SLwO
8z0KvGjTd51NP4SGQXl7P8JrK8I3A6cjPW0zSQ6LY12vaqzPJrziGzfjAzhtJclR
N6NPE4D80r0RviwSpA8yNOWak2q6P08aIQEwSRWWx1djib4w+y1Ps6sF1syH4zn5
9MivUha2aJ6YvnMTCUl+fgGUud6nHqaUn/TwqcuVjR0wNZVfTtVLg0p7gJjMWvUX
loEGokrqmRxS+FnR8wxqBlTIYpyZcszf/foZdgAwP4RMAm9l1WCNk985HTDsLD7i
wjbnD9odZGbp00CAZO6dkTCyV10ephTVVuGtIrBOJ9805ALqE/ul4o9zgjME5MiW
tLALV5pscqQw3pewr0zn2akVPsgMniEh9tZ7lhqLp1T4ZPvkVI2FjZGiw2AdpmLK
uGPGP8wVXYIMoExXSMQ9sPKJNJdP43MM1jYleecTvXX0fgSIuv8PQQeZHE0rTo9c
Q+BQAEUMZNDa35yTSAQp36/WvP4hDOEvbdJ0epK6B2Iu8sD42I6Wx/QCSnpNeI8U
Jb3dx62skACC34l1OCfSCOEPVOGvMIE+D3DqthaTsHJnq1OZddoI36/P3UuMNWhr
1YqRl743KwBoh6nyITvO1lm2wqUWbLzBzNKrTl4hdUyn261nGqwYw1H0k5G4RtvX
nopKFKbb+I7HCPTYaXR+FPXSbR6IE/1cOWo56UxVMDgGw5M0KnPmX0su6qgck/jQ
PYJlvOCDXNonBFxx23h02ICf2jE6hf9QyIy25dJBHvf5h+wuI5q772p2A7SjKvpA
AEw6toHUbp7LnvKZ671wXFaV97Al45L4Lbz9a0EGd4neWubRHNR+HHPYZ4OOi2Wz
069kf27IsN6TBeR3Z7zOIt1D3SFvGiyxVLBIH157jPNtbeIJ91makiJqo4rVcQgZ
vDHieRXMpmL2HLN7AfPVzaWfYxEVGqtP/kQ5OiR/LCapESkSnbJAOAVWpQuGnht4
xolzsAD374tDqz7sjYFhNlIiAaHCVKJi+Bdj9gPTxBVNsg/HGPe5v170xspvkmCn
vkMRFEYfQripyBPGb+Nj+cAVck78Yh/UkV45a46zdHdtNK0jcn2h5sqsW5sKi6My
xRVLA3362xI4vem/ZZYyeojT/eL/r6ILA3riqB+FljXnAEcmQttw+nMGZSBza0hZ
kR3yl9BAi5c3FCwGuNFnRloOndNtPk8n8tBZSn1dtAORwMeN/WmX3KUMBgitm8nV
+0pkNGGgrUlxnj1ZZiGEnYo+y2bVx/rHGrUchoikRLAWtXIpE2aVnkEr48ibe6DP
RU0+cp7Iiyv4mG0B0BLaBRjSjxjV0jBO2yyYFttQtXUaVEG5Tz62aOiWTSDn319o
oal2r555uqqc6BhdqCesaXX4C3V1NCGyfShZHFFQxewhw5LmiY+s3dl45V3y1aMK
tiKtYLRlV3diwXkMSyIi2eGbtkUPbxepO28RC1S4MGRuI+q4q8GA2OTzaM5vhED3
xpifCxPLRu9HwYmTLXyZbf7libMTOIA+L8BCrSsv93daWWE8s5PzMa1a7z/x0+qQ
CjdJ//nSrwiJYEYnO6ZxaxzAvDypXSJRr2a67BO8C3FoqEWEE29bn5hpc+F8ZrWP
aWY0iXsswPoIA0BR83xCs6Q2EKyoCf6lrHhQez8FkNN8A7TBJzf6l9kqlW91N2MN
BIL7/1Wf7a7bhhqAfTnbMSJgiZUzCaloOrTPEPcRWKEnr3xiSuY0X5epuQoW5TyX
xo2cF8M6lCtdcHWDGvcRXDCYIAu37pR5S4FgZH6X2yICAlaOp1XckmlEt3vBweEY
auXzLX5NCurYDzLkuhInY4q/UbHCOMltotRX4g0963nVrN1+OCtOyt0l2PC560ue
fDaHpOPr0lLbvEOzYsvx8NnzPBzAIFtqyTw4lkGYWUe9IIRLhUaiXBg4rf5vlkbJ
qv9IsNMjrCbik/vM6JOeWSBzlTLbHMVjrnI1t3i5yhQbnIYV3qSyWjBCdsHPgnEm
BKwfczk+xPh3LZSxL5y9g3MIfakR+BxTS3yCRFKtH4MjK7fQALTXbniy/mEkgtwo
HiEI/0ajLEXcuM9QS0tFPo8KwZRFKphINubLILkvSyBEMkJnOPRMwQL7eEvQgz/D
LVlpfzYBGMa4Fcrmb45wvltV6ABNbqcYyZExeleOsc/88bzny/3+1T4BKUEX1LGR
S49wOVsQzrTbiZDRz1N+s7PAcI4NpWPsMb9LG8HldiYpfxNyYzSeJYNYNxZYUXCa
2uHHNTUyB3PKBJ2yxY0R9PAEEY2bdWEM5JYv06E9q1QihAXIfOA2bqkJhVSux/co
Qoy4LO5RxtMLqqI7antkwdg5uU3/Mtv+ZzZXYRIdIigi0d2z4XQeu+HzhTBjMkn9
85rhYN+oS3SCIh7SRVPc3mo5tSV89BBiJ5zd1rF1oySK5Piz3m8C1RcLA/OI3xUJ
ydg+BSAzkTWNDjh0Rv2ir2cQ2qvfkS9U+nBD9MUwrJkjBoWHLE6Q2fVRyVH5vPEN
RQBFZbZy2Z4wiRphOKE8akRI5+dG9C7i2AN53evYXJCIGliFj5z5EQ3yJ64ynsTl
3GcJsa4XiOAg8JkkihAYMIqkU0WJkPUgMGHUarNptMogtL3devfvHrcmdDwK/mIJ
eZ0VaioV881yaZ+9sChD8WCjA2onYFg6RJDza30LaG91agn2PIpd0FulAxUujsNP
bHKjB++lzEk1mIVipjrs5FJTbmYspKZ/HYD9sXI88AW374gNmUfEAJgz1wxbipnm
4PdJ9GU6GcITV8WnkFy7CCwf8ukiqhuln/MpWh7mei6TRCscNK1y9KsWUhww6fvS
Z2YXNOjUuIqRAX5xkjyTkP+D3fQkh+BWNTqczmhPLxua0apSRRrkaHoE0p14Znji
qQKbGmwuQw2BX7JQsnf1orSWGvDHM30OxInAYpyMUP9OUQR/UTAvpLkm7FfrIajP
a6jbLK1OiB8mpLPZdZOBH5Rxf7tSa4pROIJ4QI116uihmHphHH3j7xruKdTQsOgO
CbWffO9u8ZDZtVn7nbLisw96ztsGPN7ZdQAK2hyCsVb9qshdve/My4S5WGVID5vf
tbisrB1KsOQybOK/rlrsWtGmINKruBRwr5xgKqdGs28dM/bLZdBDx/mkPum4ELNp
en3Ls1pxwGjssoKtgGznpr66RXX6fJo3GfNddhioSU5zq0OTJ95iLuu4qtPu0JBY
ho0/2hbbwSi4nnZfzpRp7/LBZ24iE8LHXjuFeLDlIJVNn9cUHPu8tJxtbwd7vrxS
Hp/FiD7LQwI2hbV5ojrfnH7m0BoYCQeiuMzoPwqKm1wrz+/zDQwoQRntsgr6JLyp
N8HN5Azqi1mDWnIczOgrNI/bFFExYodf2y/dQz7IEPk321SDC8jplXidf75cpVZ3
rpbpLS+UcbypT200nqWirRlMKAObR7v4mbUQ9VFvsel/Xuoho9ce4arpC1HdxCsc
j99mO92LVAaGvP2P5dEhnS5vjSGeq8V2xAuSOfk37OkivkjYnwO3HglxkUcu9rO+
fYVqw3eTdKbX0Dw1lwTCNqmbGwpIGUAI8o01JiKreiSRq6Bs0yEaIDMALFuja8fx
YiRYDhzJxc0jbJx/02AXuIa8thCjFpr8ZF91Us0vWgb6p38ICYL09AslSmfxat3e
6nQ0QSD+6LcGqVxG/WIl73hCXxclCrYJ5i2tddn1gJskQwaiB8X31C5AFaCpTWXb
hwNpfMf86So4TXJaF8PC2xOufX0Q7e1fu57kfTAF+2HMs0Zm5RP37az5oLDfL3GE
SwUrN46dMqJ2aJj4c7X3x4GfI+ZDwVCuRViBtqaPYi4PUvPhwKZtig7xi50Ci7JE
obkdMRIBWUy63raFvgfy18GQP6IvmviK9Syw4yr2PHUowr763/nJ5EkeUel8b+jw
iynIitFa3G9zyChk5Jfav3NN3hUFXVC31pt/eMuJ1pLTKMuZJODaVHseuNNJHPoi
CjdVmRmOdkDsZuQ1YAtrM5ZDecHQyIvwkahxIqaEklHfcU+n3kg22VXmJokdscnG
5aGemgLRvfyUwv41SN7AGKJdkdXTt1sqwAoWBj0tQIiEyRt3Lx8qIvizMG7wkzNH
zcylRLc7YKInlDsSfHRZ90bjbcnYQb53DIxqhdPCK35vADOA6BdEwBXXwYlzjQHL
hxw9NPEr/bFy9TpmFX/PDrAkBYhftbeG2b1kZut4DI0mo09IBI1+S/Q8/dezF6qC
nIS/7ctZ/vZJLud+Uavm+GPvh+djqw5ergEEOnGnNjV9+pR2Mb3H7V/uYxftzmbR
RPvbNYooEqJMg5ybMtYCuKHVtnPsTTX5n2erqq592s2UVeYpdEOmpopvqidARgNO
/kcdbMuuMizItHeynqvNuRWfaUcJYCNo6r8dQW6IcaiIe3CGLPv+j/qGYH+kqEgG
0Q0os/EaQ70P3jZ/jLcNdnLS879YglKWL801vn9C5qj34JzKtyQT2FBl9fScUnKP
zBsD5Tm+lbALj3ADXJ5cTKfpApk8lqG9R7XZuGMJI/6Wtgfe9rk8mnc1fktqoJDV
LMd+SE4KOx2PJevAXP7DLOvh4oot76POJkcRadcWHEAbU3j0Zmqor4dpkEHYtFHq
8f9UDM8QDqjdia02D7PZ67I/YZvBJnMJvcAhoVekmGQZW+9xFjXU52zD0srHvyFg
1IrJYJMaHadeP7e6awtC3fR1pqdP2IEJ/Gg67PRNSe47q4VHd9b5dk5t0MgYfPzz
LFjoX5hbeeo8nRloS7BZPLaamAMDln93WiZ9rbMf4MucE0vfFIvjtkkWIz8UYV+2
4GxeIGjmdY9Z3VDysStga8kZvBbEHBOTz4fEFFiLiBSDkrCz8Zcw3cvSavD7L9bK
epRQ7SE+Inj1Q2Vy3SeG6K/IaJj5nWgmdymdUzKQEjkWTt/Ew/SQSZjD+i2e+n/Q
JS/MPokdezDtpHVrukIYEFlo6mTod6ne9tpRNEdtkqO9h+4pYtcFtkkOLKuAwNhc
teddYiP4t3YAe70I5ok8F4w7pXPNqeWaLo87d5tDyg6tfsgyhE3w7KpDXMrkBtCn
meOi77X02M3tkTWCja8+VEVpILFPbLF4M+04mMyPeQrRokqB3/1roGBiDzBtjJ7P
3e4j5pgjKlrqLFezSkLm1TNWPP0GLrmxrM5Xs+TbkJwdpI7LO1MZUJDexdQJA9Pf
LOUO0PUFdKp0xGtD/IxjdTMhy8hal86jBv34NtLASO1xfjoj5XJU6g2fot3hqthP
3kqq6u8gGoYTLFim3MWyijSF5Uvw5aaBn6jGZ4Z3RgEiUlQsxQWjgjAuPXIEVogQ
biuV1/opvOItR3rNyVKLNRhvPGXy6b4AtEL+w5Mk/X1fMTFuWMvVqAPp+ts8FnZ/
JC2AP4CsxbOopjycOGZJKrHMt9a8ayYvb9kdmG1qiU/qRg5Vv5NIZi1dLTgH9R5J
60HA6MLINNC0sDlJJ/k8R88eRN2ZLc7UFiprIvGR0JDb3mFUrRwXsj6b2H6GOS29
dLbXnq4qyVebEJtPkrcPiLKirRh1qNUaoi4y2/Gxm37Yxn8igNneeX/4G/X7a8dq
WMd2u3+3c3APiTIDUzQhSc0ilzlsIaau0rxEY3R9044Xe8xPo0zIQtQvFrrRiqXc
C+07zNvdGYXVDvsbei+9DCQbZmFQ0FpW8CLq71lMZMYYEocXuACH+a9bX5rB/cXd
BOqRgHhgZW8V4ed0r44/HGXCiqidciBefgu1Dq5XZWieNWIioNk9b9LxStdEbHSE
1rg5RXhJzcaAb7EHBANhFF3G9CUpghQRnC/77XiRNIn4HlgxFtPLC8wWEEZA+4DS
H40fLxLjHs90Cn0Wj/YvJY8V/L+qWv3M27lcDa+PhSU/qzKKp6Y6W1MD0z45HYnd
vdXsdfW8Wibuud5S/4Kxw7PP/AvWQIJ83tmRDaVpaFQIfhRB1dRvmhGoqZDy0Zrj
tMYDfyo5hP809RsJQg10ng15JPs/0kDmJqXtsNlgIwFMaXCpe7TXw6MsJh1hRSMm
Po0IuXIP6rMfz46Sgh35pyoS6bAFz5AJv8XQ8bGLWD3bkCUW/UIIz8ORQz/9bhC6
dLKE6ZA8tZRBWhtqLjNwaRTe6LPNnWbbW2KYTuwYo7ye62XDK1tPXHXBAHqUa1k2
1j+4ZeoOtCoulHqYQ8yABSeOeb9StcEG1nx8iJDTCLZ7XDhmWGiUA0R3bMJA2tlC
uRb9xeBYTSEFFlAZXxuguuMcZ6L82hQ/uAfZIh85W2kmVE5gOmqpERDNwG0LjCY6
5muqU56elsbKVuPOk3tLgMIiurGZC+QSjD6bXG3PcYK4EqGrp+5ZuuEm3gMDZMm9
rzmmqU4Z8Z5QZZjBYIoGKwciqpJVB+tBzi/Tf3LZ+pHgOsRQvcaXB+GCYLQwvoDv
w/DTD6CnkveuP8Q1jaQiEOg2Ir6nQC/zuqRo9i6v2fkGzyo4+cxWIyEAk2F+BHzp
7Y1k9a26XHrmDY6FnT0ifWkIerYd2kIU6GGqVo31hTEp2Ivq6VWiQ7I6Y0A/BUhW
WG9ATW27Lj5w5StwBFaG+5IjENZo6IIS2iYGKWHCZJANAW8wW/BVdBDGg89SrJoA
E8c2VRirwkLP+GRt8VXpWIhBOUZxaYHCnLk4OTMl9mLsXOR0Gry0gaW7kz8+l1Of
j0b/CC0tn4cM0Hx5Y1Q0OnNyj2S8QaVy3g/GdSxjKd5sCqYQMghnyr6nQjsh+2do
bAYcfY7I+YLNU0OT0vp2nvIYTqozPSl936G3FcIluCNzd8Qj/VKa3N5YWOcx/2iN
JSfYiZNnnoinoTjVjGeFE9oNDRqFncr+dJm4Av/W3I49ycJ6knUJvsON/dHMAXr7
SPtm9vsWNApoRmTTZAPyOA4alQuK1X4Qzc/5shEvbefuAiX2esYRNMqvfrVrydyT
0WhYWIz8exIbWk94Xy8KLil6wkZE56VepseBIDtNZ/Cs9nBp/JWQ2NYJkM2ta4sx
hBIe8lo9EbDG9o9SiTlrh0lz/jHeURN0qWDtAllkQX9pv1VR3vyL5vwR40gB+CdM
XI46x2tchfm1yAzsT/hJ8MQTJppn0jzyjO6/fCE7hxfjmKGzISMJPwAtCzZopQbr
1p3EGk1kz8OZMeWOX2TNPQplIx4bWRaRkcvapZFfNcNgMzMTYs4LLsQg0iDL7zFx
GGdLH5Yk92hhiNAt/CkDOYAU1U7GpffNv2uqaOBKOW3wxaY936sQUIa7Uf/2SF10
FTm0q5c/0VlgbgeMrQ4Aalwu4D9lqGzlmmbe0OSc/iaV+Dx4DULHzAFtlNspVRj1
2BdW2bzJjsfa6DDSA5Ad85lFCY1cQaC2TFYqrRVkYjVyKZYNKeFII6qgINlVC9EG
nQ9fyMUZRIubdbG2Y9v/t7glnI8XTYYTsrJHCBNQedNT/5Ave0TzAkKdKTnF8Xbc
98J7AUPWdaT0roXygN43b48XGleZsjufd/n9m2E2Q9W1xdesvu//7D3FhIfgOEtW
qOVlIzGyva8rM3lNz7ABryFCrj+/t/jMIN5Pb0DCB7dDjSIn32vjT0f/K01fp7Rc
VCTmYqWhKtOAL0NeXQTSUnYXI5Rg1RN7WWVCVUal7z1meeJl1+nVjVCrKM6F0X22
1YpEUhyiP35ACi1+hhhVJW1tsM4WVHSzODXTC4YMCoC9DclDge3lvEweTrM69J/f
zThW2WFG9piwLhWQ+a5SHXrFCJXC2j1BNoTIqckhDS+jCuZ3UXJpt0grG3daq3Ok
WAlKoVdb6mA5dseAS53ZY4tvA/dRcvefmoY2xV7h06eem+IwyM+SAwDHrpXx9HiF
h5N5GAMdddT2d74JqQ6hNwC6VAKSvIEq359pWvcKw110WMXCld+j1Srd/FhDS67D
/7tj7Mlb2jY/xg7ji5Yr/t3kNtzyVo7LFM4V7qaN6hYo6U3TdNFeGWoe36eJIsX3
NmwJQqRE4VKfhB2//ASqCVL9ZAXrivzr9LKAOM3AXNDIZw0bzWq5gE1tJIcIzNBn
hiWATcEXHYSV+6Zn0qQEQw==
`pragma protect end_protected
