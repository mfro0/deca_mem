// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
OhbZWQvmah0ViivTFesSHSTzMaEDwBorzofIkRUkfzCwaz5dwf2M14zd4WkUwaZy51sGJChm56fn
ZDMMaqoYdC4GG6OxkwNOL/UgHs3C+ogyzzWNp2FsDQOUF8MC0gpgow3FufK/CDPh7vTpvhXUT5Dl
WvDLI57nVLcSPANKp8EDXyR/G8PtRY5hxvqqnrUa6dKftRjjLsMKeX3HO/KFeAoAXmGLMpBviD+t
avW3WOp6Tc4Fderwr0b5vdwr+Pqn2jOhW27xHJFfnin6/fNDvqJW3SnOWQDe2ue8CW8GBYWDLGYq
og6Y9g6PVIpMnlWdHm+CNPgWNJ7xw1ZQtzpnpA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16896)
wdRfME5ExbNdxg28Dr/sCv3ZiAvC5Lq4Un3ytlSxOlIzL4cn/ei7kl8uvP7MpI+aE7AezfDScs9k
JQ2u6E8b8LdVrDJ9O7V4EP3roUHMrxg89jEvBgTLoH+pyFPf1EaqCqQBMq7vxPBLzB/zfS6hSuPX
jJ683r6hXRPeMXanXqdLSU0OI+hZPiPrcb0F8jNJccjRLMiVL6cRPtBRBcH9keQvpwV4Rq3wEfDY
bfZS5lXVgkPHZ4x8/FbXdOpIOvBCAUPJmB8OsU5PsvEB7SV1K5z6C1Z68RSa26HZTXl9pbgJTPnW
nF2ZrCxbuOCqO/jNw3LvKsLg8FqKw9btLRFxWK/0x2UTaCBZcbDiTbIywHR7yXoQ0niBUkZHdlTr
e/yP4bQG0GCQ88+IhuG5JknbgZKKqT9e2snyCRLUFtFdi2t/szX08w/Uvt6Mbgct/xIhHfEAF9tR
zzDf266MfuECwDq1zKI02+40aWkxQ+buj+Gi9xjfhd3/RL0PYJppb96R+nsa8V3bnc/uHZsrwXeQ
IPBfEW4RAO+Zot+xWpqIT730OCmVVY4gR6UQlQimZd0c+rccYrppdSzgzgTqmSFS9nALlXZBaoB/
z7nxXH4emeXfnT2DGy2/V1dtN7usDjDYjj8MzDaLQVibvd8RSu4iCKDxJ/lLK/5qKLSk1ZjiFCuZ
wgokxi0bPo7U0paNDHtrHBpFEHo5n+Ee30+S5fJH+5s1lz4fjeJz9YCxlKOVXkG+uAy2Ke/HgDdV
YfE3eYrpN3X/l1vQh0H290lD5uBiA0nCclDWG6LZl2FfHpBZLsshJuJF6TIgHw+sdYdDmbN/83XP
Ov+MuEm3ecUZBiP53dKZGtMAn2cZem2XiDOvyhoN5ckd+NjdTkg+uKdZsoWazQfcJ+xMwPQpfu4E
Ol5TcrCK84lMQu72cDRDalgvRbNGj7VExawNu/gWaGuIjM8lyjOgjhxmemepcHd6pbnXhoOAUOX+
Ijh1uofvuUOOOu/YeL3O6svVu2VZxwcty3yMvoDfcnEkEGiywfalJaZE7XfrLvk00gMEteFn+t5r
52I0JAiNTNdeBNmRdv2DD/SZw3E3hOwxYDuL/gwR/hecENe8LStoWELN2UFg64dFbaHk2yXg8gF2
bxQvU5AgYplReRJZEg25HjuG44DGHsRxcsXWfLhuEVRTY5H2+Rx4pj7lLgaLQ/4zqr6dxSGdOpO5
/QVwenlb7oR8QZ3JkTLcX9JiKAHYoYxRMOQgoDHazBthTmtML2N5trgHtpLy3CL29uYX4Ff4Ms2n
qK8kterjAYmH5hOXyEtKBHsyzJ3EuSvjcWyW3zNcKo4JD0n49KVg/V2gbeDEQ9pZwpC97h1tfgRm
7ZvnoFcw0TLiiohbp6gSoiK65yE5wSbwE1x/2J0/zqwlz4H+Hh/vxzVht1apRibNN5mYbgHFtJEx
ahmg6L/cdS6d90HyUMpQUrl8BLp3lM6148WOCxAQA6tgkXXbGxZ5sgflCz5sgx9MU2TMgKF3geqy
8rmi/LyuLzTVKQUcOqh41hYCCSUtQ+rRBHLywaqi0kMI2Xz7LlDdoa5/Z9pqDtY3LLajPN3r5dPr
3rC1eE0uXUehKHzLoYjSrrv4kTpJkDUAhtwFkV8bh98pNQC9QJ1y6bGV9uc9e+IDA181lnAR9psL
uQgTU5lHNm1Vw8nBs9NYWFIeyRfZBxAodF+JRCZRMxsN2W/OQAKdQCiHIusWuL4Ks+y5Se7Yh6pL
3MHHg879VpmJqFXaUrp72LgUQMvLasz5VTOx0//i4/zbanwr1b2st91WIsWHjv8+Jv0/SkhoPG8k
vsKxe9jBPPcVEAX56h52vFmG9sa8vFsjOtGlrCLxckDlhTcf2hUjPC907eRF1p/JOz3OCLvXHcTo
0dMyITUz9QbqUT/ztPm6X6QGTaIV+SDs9gZbqYv3GMFQPcjsywxr3oOQK2HbygW29QY+51mJ281s
7k7TT7IadqSyrLoos5LAd8KH5a4oLGs9nQ3Jra4yL1zUVE9MZiGtOG7/ixKUxSixlmSaScojiemo
IFsK/UrUGtbSW6HO2WTyupdPpLD1lX4L1lSxTNL/u3DhjeAHleGa66gYagBBhLvytv2Fj8gSTZVa
R8EmE+iIUxuPLFQrwmD1UXMtCkh4GAL6dpvIfab8RJShrmOPYbCyKQzII9eFANlGxr1vA0mIRdza
pIZoLkksrdQjdmd7897iCelMFFiUOiYF7aagqevVSIQPbEQwsD2ruDJIYiHm+Wu2dqqHqDpBsNKZ
qU0gQ17q/jcNelbHFCwXLYjZkMkpxXRTtzVXklolEn4++xeR6D1KZrhzTyE6+siAWF5kXnnQpuKi
wp1otqxBE9x577LwJWFKzTIxvy87Xyfll+rBC3sTPad64mSlIWjNrmvCDIEd1TJtyQvMtoyFcqjk
eePSulU5SAXbsPieNP94qY9gwAlYyB0wM/RBVjuoj1t5AwHs3fS7/X49LpeNKQ9p2puruQdS5+lT
06rsXXuL5b7iUDoG4ZWucjx7epindDnVoUB/107dW1eJideo9WzHjTsawxObr1ejQHau79NRA0TM
o6ZqwhQTPkcZqZkIMe0hH/bbar8/uizcdbBA79a0DVFV2TAw48YqtZArfvyz43YdkYkRk8pjlHeL
sI7bWQsHqCoNvuwMMsT9ta8LDHqHVhR29IyluMo0BkS4J7aEni2P6ieBINSEx8nQu9W3ur55DeG/
GiwSYkVLcR9ghoGDIgN5oILXGHgzCq8njElNSUcuXEVKNKbg+U+3Ua1V7xeCel33gDFWEPpuO8Gr
yHiFwEcMjR00kYCIsolAej/2lDvlVNDKTVc14jCWu9/+6j8RRSteAs9TzO9MWKxF6+Xr7KU897to
APUuIKzbpDE6JF1JYq7K/wsRRMoyqY3hBbVL3pNVtJiBP1364fT/s8oRzBW9tQZigqL3WjYc2Mxj
KESSwLoSOv2TEBr39lCOeUloP7iYD/x96v18d6hbePWnn5Yx5DwNzpJjCOtGYrbHzWWGcsdiImsD
vwCuE2m5iLE42X3i/zuHHuMJWsFbzKWviD9S1W3jsQyyIraiUYPYclhmFlMyLtsIWm/66XzC/tEv
yxjhU4c0RT2RKzrUWtkgf76vrad4YVsvPlscYxhNKtQ8xsRXnxmW8wru2zcZdS/7HJ1h0+PjaFkh
8Xv1dR1gbXrXOWfiuageIBYZlPFmg22Jj9RVfpkgNki6W5fpiPIXhLGY7bzu7jiQHB3K9vB7/510
pFh/0RcwHeCYR5sIRKAWmLRTcZODWq3bO0pIKDZ//SwP20oBMI8Py6W5iMQgyhv+ytrYASedXxen
I+kAMLEUPnFHr9yeAe5//huCE9HspKmV/6I9LeeS+yFxPlNgcr+lWqoWuweSFPXlmSFIxF1LFzRP
fLh1NfLykceUX9rBLWy+ulG9bZ7M75p1rj1mNEAYlqiqzWeQ8VIMyatUN6/V0o8dw3Z4V6onDgPs
kVsBXMjfxkJqjmzRfbGxCOybp4J+TdwGFAzuJwhoz3cKcKMAXb1KIJi6Jusp0h8IdeFuQ8EhOOeb
4FR8vW67k6aLHkwWrlT/RoeEJC4vISIe/EdvVjwGKw75CBoBKOVV7V8AfmuX0mZjy/w4edS1qDQg
0t7NGDuuDDkKi+gRMas74Um8dpS2NWW5kCUiqIEuQr7IP84UNiRyz5DpmLSb0M19I0o7TXTkrnbo
LhjRlmOLthkxNZTaw7WirH6ePKGjHBDCsWrDTOdn5kY03A3OnW16D3IqdZ8hjlEJUyvG/7l/lPQh
/MYZANPxuRO/hlqbdZSjYm3eLyYSarEjRNBd29kHMyONU/LsEwNwOIhgnVsIihtFyatapYqfTJba
uhRbJA6//g1dFqwYeX7QBCohv6p9rTPhoObqF+YKjoF4+k2Cqv706M7TcfrshDxUqcaQD6hYOzg0
0NxGSQJ6Vl08zC6SgRRWPXT2+kL1w1/Gum8YKatrtIRjgJDURCirBfZbeXbgl37Qyx/nTfaxPkMu
30+zllWZTrwTWnVTo3GEsnGy2382fOSvYPKiubyKZZpr/0YLpC7Y2IfKJMX06CF6Yr1oeY3tvmY3
JhmWvpWSdFuFCFH7TEYrpO7DkBmWJUQnVu1VXfAORi9aGYwXQWhYrgA9mGsPOVogsmhYC8uzIs7q
zKPWERDCbv0JmNg2Sn/iLMA5mDyMifxV/4+DoHOAJXen5NwQln35fbqiePZIoU8aks1xrQqQIfrV
gF3cz/tUR4eC5xCeP7w/8tJT3BXZfcS17ej5fF1VIPTnSIwzkJo14/Q0Il8paX2yIM2qlgkqG69b
sMdqp0DxpMF899emQ47qBkwdeurkhVPF7ryJDeZecU1JHtySh8oTBYDz//AvqI0l8K8jzqobWM0W
w6ajeKgdmiKmU0XexUFdtwKbBDWe1bkIYiEwHuMV/kclULlChrkUpQjHVzCfZmwhctPbWJN1WxgI
wR8P0D0Lq9tEHNy3jeOzKIi0sR2IZHEn6rfCP5KnvO0W8GblVqnssnnsTUhp9jFUVMPRWVs0Y/nJ
5DsywrZZHgGUPQNpq5RZ4Nkl7kVvc4e2gUgKOMUJDRIYaoBCPK0dY+RmyUNoe4Em0SeeBOj4HNnW
wC5fBscXiyy+N1EY+FnFaCusA1YMHEHl8SYVL5G2SjyLmczQk/WJ2YG7YUkFAvztQ5LGqPd1zw/N
ErhF8JBkiSFVtkJrp02oRyixeQdWeidVpGIQ6iYa6npBK89aqj27X2HbK3JL7rwO3iyZ0fpa7QET
Bsjg7OIaeP5ApdRH/qNLpbddyp3XMn5i7bGTJaC1kT8bhH7YcMDHEBijTlAAeLzQDuo8YaH/UpkP
q6isXb8gmeO3TTOB+/fBCpA0X7O61Vy6+1Xa43NDchd1yt93YcdgcGuVSzYzgcSbop6UAXD2w1sh
p0nF6Nf6prgvqWIgMlX2qecMBI3eTJLo0wPWZZwSTHn5jmXlxqAh94gjA6XMydkIXlAp7LQiJYQi
WmMdJ0VfXtK6mNhPXO0vLTY8Msh5zkZiCV0Hu/TSEr+afbcHNNQybZ6HCjykUIx59BU2L1eLn/tR
KSeu9GSxemR3YpPTj4sMHOhv+Vm985r52GQFf82z5P/xuBdIE3ExcrAwazXHJcUb2M18LaSQ5ntR
0e5B4O+qV1+Cy0yjbBpjz+JNwt4+1BC8V+s4bGvKnVbChaxShNTQM7HNNtbKsQ7w2h/OmIdLHAZJ
8MjeyxCzKZNB6tinhnomRBfr2jHgIPY8kE+ogUsEJNJtvXgvr4/pG69RlOQTmDB+9FKktD028VbC
UF5rB8mXocKm5JshDTzj1FTZcdZCl+bTihZ86jW+isqX0bssCt5wukXEBUM/yUATo39psxOc16/M
+/kqWtWJnBQ2rsmHWp/hmyq9LgJN3ZakMi5Q87lMnMFovkrQuyYqVZcJOhg2Dp+opC8BFSycsPIO
Qe3NWpu735Wj41xmA97zaGKicvjtT8+QgHkp3KyAejpoXHHUjDSXaRdDs0Oi653X+IE9x/BSKNi+
BUXqpSb9lnIqcyEnTyOrXHIBIeJy14Vgop4rVTQyXecZPCfQMCl9mDkzT9YAKUAgAPyAeSrEyBI5
mInjX2+KibVbK8jL6LRurNLW+4lcqkPq6GWxuM+DazCbfJ4zhsScD4PS/ygpcNpWBVgy0MhycR3/
i4za+Iyfj9WVnA+Osp/BPNYH2gM4SrLoGZbXKiwvXeb2jedDKnAbczs0xPOVDtGbhahsvZw/873/
VxC/BDFZtUp2kuBpFMauaJEsOmRoOpZvZtoNT9G6+UHldk9PTYPjsbHpAy38zYCmKXGT1qD4pTAy
JIboB1pUT9rXEuFKJf9F1GOvN9BoR3SzVL/c13chidAPKjaByVHhWyTxz4xn3ZGbycKlHnV5KDgq
wjzmutUaIax1CDggOh2UFiCW6tgDQ/96dzxlceGTHcoouw/OOqagKAeNJwgJ2I+jhvfE1R+qqVPZ
YLaUA3p3CJuYn2H0GqI835QIYoGb3VAegFrr/o+gF745rce4ydiGmE50ApCIkfGG8duASKs7x2vQ
XoXfmFiZ6ow0YpGUWbYRHKSpe4phTdTIfrH9U2Vv9MHgf1u6vwMSfGdCUv5qlzUbz+GyNDb7t4S4
743i9cNHMSE+Bs2lf+8/9F3WVEU/D70OngKTqHN0je0VlLt2CV9yA9sWK/ZE59ky/TlNyDuMQ5BA
scsp+COlKJs3xFPfCLqRPpiZWxHHvNBtGlq7VY2qDkzDqLeq7wzWuhXzrFVZTrtVQr2ZAhddpuRK
gUj9+kVV69KCzqmnEBimgBgMlf+7mHqv459H0mP1y1WNwqb/TyXgmJWrac4f30InfMKD1h8/RJ7a
Os5KJhu+rB/vrTLE+erZj/5EbcBYRPz+vPDzofTWc5N72t1yq8XWvVolL/RIGiTj/5Hdp6LCv8Cm
3cPLMBSV2FnXFTUlgXyaHNeOTELpMXpj5DZ5+MaKXt+SwgAnNiebBtqZ24J0dZ6aKMwBzxsznhpt
9KnzGHXstprrBQfvcabQEN3VI5/BGrNHGwfz7f9nAHX4gDdj5qfMzMD8+X9LPRtAW9gZ9tUpYcRK
IvaSTlbh8zLyWWluWsfKPaLAS3LA7g9tKdk0Pj8RVR4J6GZqF2f/tPtJRJbfyP+bShlHS25QKoHV
Xn3s18vq3hqblKhJwAgf2kN4gSVKSXs2ZuAKhW4su3mSc/Ey0+Dp0D6WhrlKocls/Vk6ylqnzxNt
nDc9wcPd8OnhbVZ6RA5Eevkm/kFZ6ZsQ5hdEFOS2Gfo1WQAQLCmvv4b5Ug2edANdZ4G28cfY9iZ8
F44BRWtmdCyxty0mJIzDEZjzId5ljEd0GofFrk96dkySIfwOgMZ80Was6+5Va/bwT7pFvBmnUoKb
HNpmwUOoUKvJhocwKi641qyb9cFKHkY/dhi24cCGa6gZIB1xrvXlwwafAFHqvp3WZKF3STUpKH0P
ChGQM0nf1Rz+ZAM/bxT5ByHLGYDEQZXPkyJNpt7rDF2wtI4M4ehDvyq2w+PH6SpI0HIF/cMp7S2g
4K8We1n/f3I0X2XwDjbf0XcthWHcIc60qitDI3FoHw4VkZHsBBjBBFDiBMgANKttAD2q2qtGZ0oP
tXV24tqTfr0LwTAPRgbpd1/f3cUU83CGRBR3PkOSTonSzwLWqp8+7ZM64KndU1epT5EyxmsnNomV
fyza5k7bV6In2MU2/9JgMH2MdXN5TuYFhdIrdR6IxwsImqlonZj9JtDnTJe7lFGtq+4NtAOfTvmO
hQ7EFgUfp6HL1SRz4bErJF6Je6egU9XuH8JeS9N9E7iVOCYpub+0d1HNfopwjpabX67oil42cuNV
FTLE22cukABHPp4SpNQE0Mby8RoWJBURHIfBV2rxSymqE1dHb367737M4HGhWsfcEAbgshTb2IJU
drRefWN8Q32asR6EzM1gIJDg8rDn15h4MjRsex9yRy7qkA3QeuCVPZj0WDSeMnUs4dVUJ++mq/ri
Q5H7GaD6jDcqJ7Lk6C3J5JkXP9NaSoEDx8ukG6sVaaR83AbckSDY6b2xqFMwlZWSBBOLTq0f/UQr
einU3cKpxwt2rei+89QFDlZPZ5TD+dl1Uh6IjqOaiw1dZsy9AMolETe+gHDPAsF81Li4o83zk9SU
xXGQLVq2rMpKVgMwtgVkwKNUALNEa5DmEJ3ibZZuAk+K1ZwMbykgQilhms5cfwXW9pmUKa+etzN6
6PDKuhRcRo+AkSXblYsrSAP3jg54F3bmByhqNFDwcv+G2XAaJMuMSbzqAFQRmi6QWeo3rJow/bpE
Io2CNInq2Few0jOYzmuZRkSIfiUkj8KQzdw/9ldch8tueKnFd+sAlemTkBGnyRzISImFWyFIkmZX
If9rCe7zFnCJGuOLQTfar4tWq8bnov4xuGwyFKff1qeFfVdTCXMCqqSkQqPZcB6HqydHNKkveV3D
sucXiJcyuVYo3UJDSH9WIm0HoqTAi2mX+ABl8TPBC9dTlGnAfEtY/gMJscw7oMANrHFhRtz1VGWU
DPYEFeQ83cPjaTqNkxTGwOPpuoAj4FdeVKh69w4HOhKPB/83VUxku4hiGNAng9wPtXp+R9tuXuQ6
TeEzdj9CzUSGvjXWpnMExJXeqXte8FD2fxPiBBIvfwAoRofZeZivC8ZDBXCkBV24TRDCpQctsi0n
8G2Si22cdO8AICbs6XmTd4L2PiwRlgHXRh0ZyNbaIr9/d0vBxzGn6T9kGdi7k9ZVkNQIt1AUB25n
uGryTe2oP/yCMFCcpXrx0TXNTngOILfCVGB0N5YpeiSkf383GZld8q6xykhquKmj7F+V3wtGIVUE
ROvpvxR4OCjHq4ecq+BATMy0QcG3pCJ9Hwp4j9cQegQt/U/PgUBhZT/BZBvWj9JOKxcgRXKdtiJh
7BSowuruuGMsy3wjAoWHd2m2aqEfStuYkFKwnjRBK/wGGEnlgSPG73AQq0e7+om/d1cxUvIv5Y9l
gJIaMfq20CbWa1XOigekTNUM6Pu+dZrOvzLmgVg1p34M/0zcl97fFLudMmj0ipyTLxLff8N95uF7
gphfWQEKsxGR7rFK8sAK0sP7NW6D1A3hijWIfM0+zuvDKhqKMSdf3WqF9t1LNjuc5S3vW+vEPKG/
qdJXvEdHKOHbVfVszmtXSGbGHasglHZ1OuZXebp9zkBscmtJOlawyLC4YP9Pq2rSWwR+05hF59SO
fDtB5cSmIN5598zrNf0h7VgSXyEEzNnzmff6sgelnei7ccR0L0f87u2jIrtn617A8g8TDjq8Qoyw
24oSpDr4n6MycFpMaHQaVkL0vGGOi22R7txMNLQaeqE0JHTJkZeYdoOP1+FAwXx7WDcbd2mAM+L1
s9pYguWvQw1+Csz2MTZtoNJ+F9ITcuIGPN5yR+NWsQaV+ydgUkPlw/edKZxoF0k/Y5d+d1floNXM
4tXxDMwc8l+9Dkd/wHBuzkEIWOsrwqCFTnHcLmp3IcHFKAYbIpFufJ95Mw9Noyv+bL2WMAkCmTBO
gIKg4bXmKC0IYY0ziM0eGbx8zuPlL1cvz0C/quttnptIlUckJrXec139pouwIDEyqfGFHJoVAXsK
7LF9/4aCs1Qq2vUMInMbsiIlvlAsSN8qrB/moYF11kh0JnMZLWXgIBOCkKPJWXOgKBOaEghAjVwS
el86uDvUf8mZ6UYyqNl5aOBDarFfSOfqlhc95gxvBexAjMLoUXMCx8F0lS4C4cXmrDGyYCYdahv/
A1oJH/B2uAAN8/ufbrp7UoKUtRAgYI63/Qnd5C4KDrWinzjEuLc3IaqR9IQGvgZQW8hKZSOYsGBm
5M0OPoTcV0qDQrjBPeWFbPeVTlTgnJ8anInkKUlDc7A5jjDUebemn2WaLPcn70OFBilyDM8XzCQ/
BULjRJM2q/S1edIQSy7UcTYEEug6lzRzzPEOTOuCctBRNVqZbk+lzC73Iu7Jme/yO3DgjjkeoShW
74Q+Z8g+HH22bUHm1kbC6a9HZhJIylDKwjGRturpBXiQiY2Lb4HO8Tvx6GmoGY+tkUpOn0+kHNpI
lqawCSgxqBJ5OA7cBFdq2XgDL12D8tVYwSCmYKxhWZJ5hsRYQ0E5+xIG+lXfoVAxQ1jWBTp23rZ4
BXM2T0ziUTgEXviA7tXiHNVsnHCIFVgnPSD5B3nnsM7hMV03cTdldKjqUxlBHYnKOrZmPxe3rizz
ngwbL5N7GmtCzHfH6mg8fQksuvFrQYlf4vjWdCwEOsmDTbV+r3nzetRah+hY7/FZCfgGQ+/eRccU
qVo+z+r5eZn3tYGu2Pc/FG7sSLs4VCLj2Lr1xUfKkiWfmH47YcXyrmGKifDseZdCgNQGY8ypoc6d
tUUfNXvaQp5Qymq9PUED7AmxFd/P7G+SUkfYkH8ZIj9JsG9ObiFtFRuqy+4l43FBYSnXKl3VozD1
/fQn+Oo54m+1JvCkxVg3bIvZvV4gCnbZdbq7rwLollXUYD/MkllBckYlLbG2X45O9OSeph7X8f/W
FdZMgtFlaZ0Y4c5IMEjvlU7HOA2z/QkHtBW2mYOXVZYL4wuclTay7nSP0le0z5vJilsPXKGow8C5
mQf44T1qRhf+H/anr6qyt5yjxMY/bfcnUuLiQIBVzS/HOfRGN/okCp04VxemdtGWI78F4YWkaCGT
3fxH/izh3h3isB1qawdj0jtJABHXo0Ej4XjLwa61ukvk4PXdrbBE2nYoy3cFqFA+jCqUwtrxPaSZ
5I3yml/W8A/6KCc9ppsOvXoCuSJEzWnHcwzvMOspxgNY5Gde9tHE5khC36P7imkcD1nMxDsnN8WD
/q2oejBi0vh/RD3/U9VwrUeJKQfk5s3nDDyfJZrmSVFM8CMGUMTZ/yoActeqOaNEYLXbzvVCyRSn
9mw+sawb8ss+uAGD2EIxc3SOOEdLq0dOvQB/FOQC+xn2P2FSs2ECVLLPZMJo+QhGIWahfT56T3wU
6KpsxSf8+Kx03XgwYvS/ZBjiJWSN3HAIL29F/jOoHsP0PCatGoiViGIxT8zCJ0TocT2yqpk34pS3
M8ykntvmbl3uXaVZ00nePV1T+vbWluIi3OjM17p2FxybcUAAunEXF2voP0EOIpEhBUYcYTF5Ddhl
G2xcn/BmutaaOV3paLT8zP/Mm7rIXR6t7vpnRovva+MtSJNMsSkTajrWCTNJa+22BtA14h0BRNVB
3rmv/tmHQuBycjgJUh/q7AVIA57u8RfBZraD4QfeaSOwuk1Sm0qYE1kJONRuT5HxEBZZFVLBcI1o
lzBttp7fDQrZsb7Ji1FkMm/ugepiEbhtAqsEV3Cf/uMcPJhxem3b+zGh2IHLl8Poml8e4bArREdX
ixrj36FGal6en3f9JXX5xbGbODE3r3hFk3OG6mjU3t3Ts5cDsBuxe25aTLTXcsP3uh6RX2bg0u+p
EwTwANcJKa2VdA9der39gm39yqbKF64BIz8qty49YehaCP87l8ydsP4C16LB8FEuAlsVPgqaoK7P
K05VPZRLp06sA1Zb7TTq3f/fqZOKmItjOgM7zb+p/0ewBEHzRKaKw4INLhC8kMbYCzdOBfCnaNv2
SDY1cXFtb6IUfQlvqo62qsc1wHaZl2nZzr301zc3UQ8k0Ctowu4bskNoo5Oemh457Pg/5REnzAjf
TSv7a2NXmhsh4T+CY+TnJV9x8sgIGs+pI7PEZjQJFZ/sljHFeJBBif8bRzfLTnnKc0Devkn+YCjM
9GysQn9AM6SWZThrlB7LeMTmBjT18DvFvD12rA6ozXeex6GzXseeS0qAR+Se/PVwdU2flrVhm6T6
NuMJkkJ8lDCuU6VD/TnSRVxPEK48iEZtAUIesW1dxDCocsEBD0waalS62M7GY1LRCQoBl+dKpvaE
mMKxa8EPm8r3trn7DGx3eVLNcOZapJCohMT1EVSHNB4AacIWxQtEQ8v/M+aZyajW58gULJn5w+yk
gOxdNqUUhAGufPvlbQtHgoOCkJjNxc4v8dqh4Q1M0Fd477ANa9LyYpFYR1PvtsPT6+Im8pET0veS
pJyD4poKPmXFUTaTuqVLGsb5+pR7fPwLL+KwIK+aLK12NQAAtwWGftqk1enJfDej9DthMtZTTl5P
rA4zL0g4Fuv2H/TvzqeRi95SUG18jBQI22/qmoi6eS7KvrWEAdey2vIdf5I+BfDvsW6YJp75UO3k
wN/g0Q/ozgoXBCg7iNgWpKjFtdXPjAst/hjdNRnRhme8+yiJGX2Q5fXMWQnC2G8Elkxp2/9ki0/8
pNHAUsbrprxNeIBZf5yvcGll9OaVn6zu2nyXi9sSnELxD4Rl8dfmYqZ5Tdiry2qJqJUOZ0+KI2gw
3VZN3KzOkPk5BjkWnAYAEH/sBJ724iG3LGrGOE5q6ccZSxKiA0XGPafxtF5zaRh7lmmH8VhQ7Keq
wg/Ea9eYdI4Arf+Bx8jEEapDfxnwCEegOVCwPGL9+iik3s7lGIpASSMS8HPWZS8sfFgwW4pKghcI
2guZ1AioJ7Lbl1T3kprVOjIPM5c0IH+uC00jfLShART+B/iFii+9icEDNhLxE5C726wqyykonLWX
tISwSYvaXt6Y/Hli6GV5TxhzaYrRYviVFB4PUMCwR2hUq9zRz3Qh3lCTOkaGQjzAwXvxABTyhLsn
Peow1p8/GzKrEil6K/DsIHViUlfoLbW4veHSFIrwdmmLg2t8QSwJR2ipLr2esntQdWdmx6OhIYlK
aZLjaYLaWH0T+OXKdB2Er1C5u5uLtbgyaZc2DziytMA+gYzQ8sDot0HMnJKGQP8Gpvwh16ObYPoC
tOxfilp3YRi/B0he5hv49EpFzgzJ7t/btmrwipL2osCxpGAI2XqFLWUgQFsWNjQcP9PycMJubP39
kkwrs9pEWQZivIUJogr7Y9NRmQZ6G72rI2xhcfdg+/XFwnEJVLJEhdFM/lOTNeLoiFtyoMmqfw/M
ngxvYbkrjiPDa/+ERFV5gkZDP0oUWk/O0ywbzQFf4RUIu1uUWlGwrEZxAr4A0ONXRhrGWKTytoVG
8ZCWWVlankGjMxBN9mrFqxfa3d/CjpUwChPQ8F80/xiliGP6OoR6nMNC7AIdcMYE2+a8yXWRQHoz
FBfU8AU8v5ExvGSjhQ+wLjNUV2Fkb/IfyCo8G3MN1+Eq/DMwkCU5wzzzcBIRiApiA05s7xhLq9Sd
87Ryhunz5Cdczt0iC/QTlnXn+aXHrJsh0dVWiBhUdsczG72SLrg9fWTftoaBSH0+6Uis+Lk+rAHo
GvT8L5jn08PTTv+dtwNyQiIz9pPwEuoXw2aAlf+HFpNiLz+mbjdnzutWRWTeCwJqthTYFgJOjJ/c
KCulLmCiUCu5+hdMdub0F4gY1u0juOZw9KI1lLlYeJd8yqXslCdEYqOZ97xpuclzbiv9eGm3LQbz
G1bbmNC6PaGMFEyj1D/uTzu13NR1ABHBRhNpsbKm+n7PFqUQSJHveWhQRX60AivR/awCj9MoD/Kf
iD+drSY5n3ga1kfKPlF+oDhLSjDlezxdBUDcOuc++4ufbvOGkGtrmEMn7yWhKRr5WUrEW3sLLTs8
Pce5waeJFeklW4opYJxcYIdgYAA2UCaT5Kph8m5io+FQV77kwEQW+7MjXBuz/ZGuXOdjHSeD2JML
8zO4oB0xZITbqiRJqxxd7kPtypmp5wJdRi3g+tpxS9ktBRMpv2aVyEhpYmFzoQKZQ52TXtOsB+Mk
I151yuKF8YPgZ/FZSFoIQmD0WRDxJpFr9ir+T2BgAkajAlsbDt0oji276lpevB99yd9+f/jgT8aK
HtNEIyfHbl6ytyzEabSbxjM2EsGf9I/9q5KkszpTzptiresCqp1yJ8KXh6ujB/BvTtfSfBB9Yb6J
OroDjIeLRhZ9hM8MbaR4DZlRZRt5EPnU5I6Pb87PlSzccpM7kovXICGeFTu54DI0vjh99vCbCG90
v72vssRkWOPByc8lgRZ3gy2Rd0so4E5g9lhYezvCm8WGHHi0RZApPfFxHWaj9NTnh9N0+nPSPzMx
3snUeqnL/q3pMqp7KsmE2ExrnSl6feCyBWZXTEUZNIPVUSLHr1ekDC8Qpz4E/BGl65/jY+1+WXW6
oOapnFuZhEZvlI5j48yRUsoZKWZM8G6CPEB1rkGHtpAeJlrsQz3GX/wcqQS8Hko6N9VFkhWkD1VY
GXYwGDle+RvR3yScASEW7amUC/AzwYWKqlOf82pk5o4mbT1rscoZNoop/VHADVgLRpHuebELX6gk
MzgHEoWb2DcQxqgGkoFKrNXnihFyTMlrQZRlw5mmP/uzQIe4cmGzaPcihvv2ANC2UBjRDuQWR6lg
noufTNxKJMR+u6ZCdyZX8QeUmTzzD3KYOuyIt2VH4SwD38hrEV2UDdcNAN2P+kkRvu/YiYBj0WvX
EadeugQ+vR77waawfpRlaBe832jD3yJJMppIQpeivBoA99fnrbfbR/4e6vKkj0j9ckA6b7yFFhbt
5QfSSRkB22nJSGDAbzfQ++b5RQgGYqfQP07zgSkYH/Nyq/WBcp+GnmeD9nmMFJiPKLIEuwyPhZLd
1djc4J8VAqE0uoqK3DrsN0P32U5NZ3id7bgYYS5Mr5IDGMFlKY215miENAER1T/gXsTL5miFephE
cHAldK8Xacr5WNDC+VGDhXRMqGp5UnVh9PpqmasmnZhz5RJMBOLB79tj7NjloMf7cGDL5BuIF14s
QCQlf++frBms9yeetzTacnoM8f245rtjfF1tnWiNrT9wl9Fa8cH/WEmiMgCJ2IFLR/r8KvoqBYo5
A/78eo5qt+6JrpUmx2ovWWpvAWAZ6d8qc/1JS9E/bmeYsmPO6mDHIYICv7GHzb8h/YLcMgcjRPcn
jCur2a1XAFR5vFXy+qv6FbH8rDBLUdRCQksjQXyg+rhb0zxjB5OaxfB9ZKDRbMKxi8ZtfvHoEGAf
OgYdm0GHTTpVck2lUNinHzMXJpx9PStuL8is9zuyRL34tkYS9ZUFnMJ2l1QDZbFfK30wHGPtWXfv
6Qa3y3y7VZHnHrZMT8VJyilPyrtTqLvrPysfE5gcFnm1ms0VAamkDALkf6RtnSZOPBQ8vvaKYHpO
9UmNWKaPnLbz0mPQy+jXvr92VCu6+7rLL2hVOAXzqa3eZReZbFIwwyOK7/TTRQj9bOF+kCcpaxl5
im2no8A7T68vJUxxKbBt+IGkVRJeos3k476hYDn5R2fGxPoMF1bpqEf+cYz7pXJtP2RJQ3f+E8ug
CjFDeO6qbL8dpvWPQxLQpDdlLKjkxs1g+ictsmGbdEVhOoTYzb9r1PQalczcFqBphMxsb1bPGuG3
8BMxw63tUHcyd6MXvIp/88HX7gKy1fAfJB+bilUX/FlyUxMKl0EqBoXK8wXRDqqXxv1rIbgQWhuN
vEfTMkSEosshK2KZgzZLKnyu4OhB8+KJs3eC5QZgvk2z7FCNHEPYuNPUrpCwWpO5yJjIxynuyjqy
uV7WTuUO6+wX2MUARme6+NnDvPJYqZsLmyxRaP4hZg7wuwH/KO1LkaBYrT739pfNO3ZDqMyvIic1
lQnrGmEExBiAFAbJQUGdjudO1GYS9Iv9biSmruDInJFVcI3s83qnvXGCTDo4/F3qhrNCK5BlHgdI
HdO1mSsDQqvOlLqUxfUOTcb5frsiNaAHeGDhA01qlNmFO0xOFJaqWsp2YlxMsT1odAFygQezDPmE
LcM37rK+BNn0umP6ebPJh2axKxm8xmKJ4W4i1zJ3e/hkDyDIwQ3mZ6WrVCijZdQ3mXPm49/RP2uc
5ygxdbcYVvQay2O2e/IVnjsCjqCFm8fLHQ0MHlXw0FVaTq3owHN/ngJL1qs9ZLwyU6sAASnrDUVB
eHcOMm1AQfKtPQjn7tt1ttU/QACl40PALjPv455KsMjSZ82Tt+/VOOP78xKnBf1REhk2jqZHhB7f
NhrRDuwAmXXUds9H0Bq+qxoLfbjFdGd0Z+6NxKH6Ay/cJsGV96iP8ylRIV2PIWJVBKROclRcDBh2
86HGX+DydrCfzpwtVnu9Trm/SS/c0vtT+eUqVuHMKHrCsUcC4gyuoLsoYLxv9IIYaY81Qwe/6JNf
S6q4+8EaSLVVptJ72gxlTxE8BibVPhtgJ6vlgJCapIef3GB7oBMjKWsQ3D3rsP3kj2bMgRYFiiLe
JqHjfnxl0eAUXy6bG0HKW7qTSVfoycIGwWaPvv+/qcPCmrLMCWIBEKXxOfb+ukKvSZtx/+sGEPo1
RMD9lGxJgh9frjxOx6v0JujGUeQy8XkT5GazKKH5led7l0Z6vPW6vsVtpyvEuV726BMm9tajom15
KarmBtj++4pxEwK1ZnaO3U9wtHQ5kv02+C912FoCg4YqMmey3sSUF3ME8WDvKtFmKVk1sE+x5K9A
qMx6RaWO0ZZ9qqBhws7vN+zfQJLupCCTX6AbqaFlWe6EOr4fm51VUIt+QLNGglj3Q7aGMahgSJBy
ou/3hEkjDD7LZAnXmrvBXFOQwjH3YpRRAqfBWHKr5+6MkvrAjkR2OWFJr7DD3Hc14WT3WGteGmHU
2xpFcRRHKXJtXEvRZVvg6/4TsdJulSEjnHuSEiYtJJJbCSvgZetPJ9gGddcgACORGlEfOpefWuzo
udZzXOlFim9Jfp7bm/gqq2XtUaoL6KVs4s0627Y5KrWp6sC4UU+EUqBmdzO1qesN2QVcFDDwJlhw
qX8T9qQ0uX3wMjwz6NpEIyWGNTjFkSTm+igf+ZVmhfXNP0PcmI48qeBel5R0mnGuU8IcwRMfIOFw
dJxPd6w8oENoMoWjlGItzoCQSW+UWBxB8bMIxcliGOaJO9fXvK6xDDK07MbsIWDE7gfIym4RiQjg
lRz35Pvq6VzYSDBN2TJx1v11FqAyE5sXKyGWhO6WgyQyxrGJoA9XjXDHO00cO678ksDTfSUH1Ysi
ih2ITqD2DnSHbNVn75oWme4tyR9qqFDotsd4voxs1DyzqC+gGisfrikwHn26JBje9BqCZEFqjVhc
tIGxxzk+qadCahekSJPoB9TxUZl9+ASDWcOoSb0ASMwZgrN0+5vknQBGpcEgK7m9GcDSWYcKyWb7
W6JCFt/aeSrUPsbyutSUKiB8VQ56ccZL7x5ROPMGDzvC4iifM0fSYdTWlY5D1Vi0+6/J6yW/rFIa
8n4or7c1h1c9r1GrnXcHTcD5/IYR9EozgjCk0Y4ahBn6TAHuCjpJP/UGAyFt1rOuL7/mT2rCo9R3
6FLPo66Kj403b+W+CCUTc/Qv+b7Ow8aV9BfIHLe29bCix6hkLTuiK2FgG2OMvdhrdxVTnTrX5z6A
a5pA3ku/cyQ9HP4TrBLzi8mAMoGmBnWfsb0+TgpWNUYPGV6dac2zZxBeGQ67YW4n5K3NjzwC1q1S
fAPwktrcVusbx36CdZmGj4b5XURMA+9uKo3zzj1kQ72goNsmXgRv3oOziZmgTCP6PEhJr+XOl2h7
PRsY9H84F1QAxoiRstiObJxB3gKnEBzfz2e413T5udwWyGnU7a5ew0sZlNOl/YD+iB6yg1wh+wDu
iuh2l8HrB4MaqD2HCgFaJ8up5Jx07nNLrLN0PglbKTTt/Mg5kYVoGGW+bkAyb1zr69I2QjFB19Cc
pdjiKHwMtEGsxImMyZc0lXtuVMdOCAYkkRx4cy0zIPX3dsBkZXmIkU5gLPxjAcBukf5x3+shdr9B
JRpYS22LQfnbkvdpf45Y0+w0ILQQ2tanZTM04ZHc/7Uf/IbGZiMQ9Aaj1OVg2ID+d2x9qlPYEakb
AK+bqBfy+/GZzUW68lDSIOiwF6VgWRNtI/NQLS+4qWsgWcpeMemAf0m9tLJYmuoUjO8mpJ5ZvR60
23FyuBkSjnkXpkVToYV//4nFItA75EEaE1B9l1kwCwAds6H4INF4icJf4A92JcxmKu8+qerRlA4n
M/CqR4pySNsP+JEb4Q1hGu/cMvoxzYCL6lZKkhFIcWzGh9l1PbKeGZmC9RGXPfs1G9JUnvfEEFQf
CfReQz2DQZsx4GFRqCeTTUpqeIiz/MOK9MojMlEiyqKeRLmjVKxP3OSgTimBJu5Xq0r025VQm0hW
7cCtPcXwUssJqSxhlQpuUtLtMhTqYt7F2sfB7z349Xh451Ux/0CWHNvN/K0o4GPB4+7s/ez8hgWX
lIpz9kNzFtw8FgNFEE+Jzevpw8iFXUehXycajsDGGdNLxCe/j7+WtnSWd1cvAQZYOcYlIvXkFFiW
VRBc/5ibqsJ0GVJeVBHEL59QmKRIKo8ySQjk1kiWNX/nXKKGPcXdbGZHgAWz9KMhtXYWw42h4D4P
aHQm3NOngNaggLR2erWDK3PwGJgA6faVR2n0rQ0+UMBk7BhfDpx/W4kAibIwLsMuzOQawWbbmV7V
v3vwZobnmkrA67tR1D/Ntom1jp9r0Lgpuh8fkN8NlKv99azNFiLVzyZsti6LY9IlrDB6pDI6Ldsz
26jtXdWR61rVVoQmbD6XOg3duoL065LLxmuQuU995L/beqqI6vA7Nnr5GVW77oaE1zqhXmnu07la
vkOxLJoJXK/jRRoWupDXWa1IIuNsQjTrkApycGr/E0n7BYRoVogo6UoAMIr2DGYehSEpgddHgoZW
3u9ImXlOFccCq8inFR1dmooJz8Q3AoRogg1hXyP4bbPc37vP67kLUepL+pZoIkTZuSecsUdFjt9t
k7RRiQG7GdQQmdBamEDCmmlveXa+1nt6nbecaVn+2+HzHF2korzMbapIXSTWzRyNqMs4U0BvvoCZ
ZDA6XzB7gjamrMueAvoVV3I/3r/NkuLPQKNmHglzoiu7h90Xhtgl4dumpXdhBdL4ucrpMGHHMKPX
pNaqSrEItwJ9Y6ykNmoiBOO20konFh3v1RaeEAkQU+KEVba3xaf7pxE7IYmrYhipOlSKMzJRaD/4
I3spLmSClwNXEvkDDLcc8yeFc6OHX5D4R43td9qeTWwJGZPHDmahKlxkRNHveG/GiLi+yJV843b6
zncQ8PQ0O8+gzX2cn+BNEqDA+CPojnlRcUCy0BzuPywgcx7NF5MVaFUp9znaiPGdno5i3OksngVM
Asi8dx5fb9BponaP6qH0/z7vMXnKgBQJEje/j6hvMErJGwUWxtGf76EOJOjVy8/Nutpr11/87C9/
xrvVXBiqSKDLQwEJmjxWWz15r6fqxXP/sOTMqjrtdmEOiEAIYrNyhm2vZbf8n5FlwD47y19PDLEg
KI0tXD7S80dV/oo+yJyKeSKcvClwhmWVOZDmNnJeZ4nYDlYPRprHL+FLERrJ02Hl0QQtJMM+Spmo
mAvEQdU+mNA9GogOgjLoww3BfJVu3vKZ9bhN5KM+UFwivMB/oY/DlITgxoBv5tFJsLhs5KEPz7JF
F5KfSsJx79+cXoijwCkooXg8LQ4m16FTgYwf6/dzvhRBZPNK0BDyztvjIjsOZYo4kNNaGeZhrHgw
riwlQL2OxUtSx4Rg7B54n9w7R010hFw+CznsW6j9gJvOcH1zIf4DGzXV4CQ9R6FcAbSV2clEOBuz
YZWuRFT7ZBkyPJVE6yiyM2kAyM/RLzcPEHKdmVjlZxs6R2OIKyF6OaNBL29eMrM/uq2c2nyOEmyk
A83+tXeflwezum2BjQv1ayMvMsg+zvoxw7cxtVLt5pAtoRP25FQpAsKvNmvtcisuWzUK3TWQa4wO
DT12ftBy0rxFX1krfGyN+2PNKmLJIelb89BuXhKB51c31Ija7S7dprwLLT8FyhTk/Z6Q0Lt2nq9H
6yY+WlROzE94PIeRhs25JoFynkYaxIKnublGgW3bUXgwZGtxBZm4rdIkV5s+0d/e139OoUPVndmg
qdaURkFivhNjhY7saEtIEviRjJpUdxXTPeJycqQJicYeNNmgKbxsKpX6qQmUkSPsXw8tSoKk3g6m
0rZXBiKBMwXKfTumfYzxxsvaQ/p9cuiuzetDF5DqtmkDZWOYqBs95GsvTT7Afyx78JU8PLz7uPKE
4V7S+IbKyI4CiuCqz3mUkz9CYWnEknI3p7a82mO1LaRUqjbwcy0MNJdvvnyIqhV44uJ1T0GDq7if
42fWya2ZA0sDxGRvOTlFdZCAsLIUNNNsgK6y+vazCAen+6JPawaaVcbXqClxXgDmCMZ5dod5PPJZ
tsD9mTeP/aQlfMfR330+enr4vmXV5VSzvuPp5mjwM2gfXNo0FG73CVpWhBeqzNeQDD4LPV1GlukR
23NZt9m57Lzdd4csp0jLqGigvmunZz8263cIm1qJitlIvpmZudTB0vXyZf9aGXI/4VXlgdcqw2xG
0ijqR3cHlJ+sJCydOdUqA7y44jmNCDbRFgcWtb0praAezV/2rj5g2NBRWvW2jy0sxV8/aUMJXeJR
EhvCjMBsM2JAl/fnhDmKTJQDzbPm6r4C3YheYGTO8cZD3fY9IZsJH9bVVScWhfBrMmkS58RN+12t
EwdmHgnLe9mawdwoPX0vK8i+uqQ/BjpvAzqNsNCl9Arcmcopzo6wV4UrUmhssz+cf6mjmYWii1vs
ideFkE45H3M0hzQaHpe+Y/REUABCLn/3rMAYLfQY8CblQ1tTN/bLYIEo0yeGZBZ9OuIBc90pCuQ3
xnMxRy8hgXuP/ZSvbbsudCFsvzeojRvR7hdnYb+LdgAfM3jLp027R/xwrvJ8mkjYwtB0SPWovH/P
T0NSUqzRsn58E1IxsUd06wObKQAmN9nVWht/P6557lUQyjEzyK1W56xW16bTK1MSjma2LW8tAROz
RaZUcCYKDRq5EMrsmBOf05wsz6YAqATiLsGfJ/sUflvo9aTdeoKXjpVsv6CCiJF81eRzvk3eE6bO
HVPr/qal4k+aOSokTJBVisAtepdIRkghVm/npl4nLCM+PKsYV3xQJfICXe8QAvmvjZqF/kXpIJ/8
dTYWMo+XWhVLZzy2RsHn1kZCZ79l29KSf/fNW4j+qEX+jLVtm7DB8JVA+UitEzQSTPpdIw3xq5Aq
IN/THM4bbluK14BoYDiyC7hNy3bVRltkjtj756M7+4+mzoz4svr/655zT6Gc3xy8UPAfU6XLQjL2
d5cqiUCM1WMZO3Hw6O4UpbDy8C3N/NT0UXmrybUwLLUd753BWfReJK7tST0NWx4f1HJR0DXkol7i
TMVNyHvAcGKMGdr3fuzOWRPof98IpFz+Y1bKEjPYTp3Hc33VbVv3oWXC6jXZwENh76ne71X1tPEh
N8ssqOvgi5iXQAta/MZjfeo7nIkGQgezUk+DKSzvPUn2a8OvktD413huyV7xN8HqYiOwyDJYBBB8
BhcYEakLOY8gTiwhyAAiYtr7SKf7t67n6KYkqcfirHtk8skivOkjYUVt+Kp8C1t4Qpg2ybe2lWDV
SoxgeoP4kQ8FO3w0BYo9O9i/6qGNj/QQOTgIR9sj9MdkLqw9Ljr2yBbrLxjGZOpXULiVJgTE4i3K
xkwjytKCErr0hm19dqWG8tZPJEEDqCVRZ2jAGT4eEEK0q4F6FbzzkMD8MkPon+jXHJ6GmmSgoHFy
jhjT41gwJBKEF1zE3V/sxjM7SgWpW0qrxrWRW5R4HPTyKbqzUlA6vlzH8YBHnMnZ7ucYjtOi33el
1rFwNBc/DCujdJM0sVMEUiAeHOYmeE6sqsy9RW39uJBU/p2/ciq0GElTOiRCsSvoQGKMKSCCKUXF
E3l77XMPQ75KpFPD5o6Cgs47I9LxDtqz26WbTp2dPssQRU9/CtuLwgkY0o2xAoVeznlI1/5N4Fko
SHmOlC7AKvzyQdmqoke6rEpY1Nj/ECv5ZLf+e3VP/LuOSyKkoypw6u3i8OiLk1GCBvauH6D4i+xd
mri7/n9oFXHCNyrjD8qkW7UsxoHAiC6QCvbOhZq3vatsASCcC5yqzr27SmgAz03CIyAeCZrvB8eH
j8xG+4nsBx4gmH6xP6xODLouIhRbsdZDZgq+g1FyANU+83v+J/mL5G9RoFGLE5BxdqMO2/1MM8RF
mcEX92mCKpAmhuywNytNJGKroYCmi7hMr+bfu6nLTYZWh5Bnd7haonFTUw/fKE+O+jbDTPnOdC90
B4HjD78vMSRWO9QG49Hjeb0P5BFuxFlMRcii4DJCz4zuJtpCRnckGdeE6EifyDAWFg8FvyD2+XSo
x12JAto5G00P1CYggo5lvGaRBiKw8V+Na6aM7b/la6E7iM9cxZG5Ip4zFaszxZzyZn6nhO75cPTh
evJ2o+CBqXyPOWQ8Th6vE8bFuz31Ms/uPm+uiExplB+mQ4L0IyeqDRP/74oGouKgU3TSge3sjl+F
22qGc4mDbnSVPTeWxPN2w7XTh0pFUg/ucC/QNTUYAL5d/lqfdDToX9ub1RDXzMvic3G/hvH62dTs
FDe7G6FbtT8tVvFdcdInupYOoGB/6A3SOVSZG3kdU29q2eDKsb8r2FvMzrpvSaty3v7FVfupBi4L
HbxjfcmhKRQmP5WHLkFhh0Ju6eqdZysDUQcPQXXUcK1n1P7zCtoDnz4E+diGERFCgGMhusVsXWKu
hJUQTPsfrkQlocinOw9a5YLPCsB9YOUFsAi4DJ7Qq8h+smi0ffC1FHZsHtzp5ed9VWFMLHSaDUgl
3qWN6URvfTdj/tVdWvZ4C5bJ7YAx4vKrbUR9ZfIKOK5lPWFWvaiEiwpxcwdebr7fPeTGn6M5gSWz
oKr3McS3wscjfZhjhLfq6BdP/a4ZpBMkiK9bMuttNFUUPdnvk4nknRw27PTBhJzw3rhydY2xE+aC
HuhbQcc8QPjuqMWbY2jWRpillU7Fgnqv54IWWTvrlTtjUaU7NoONKeY4o/Uxx/VWP/Mo5wl+n5wQ
RvgjgAU/fuDrkete5Yl7D38PoWbQl/wYe3cr9zrUVOl2KL3OKw6eKfM0uXlT3W9tH/mbUlv5G/jF
w2fBgkXJEw9K3jRk4/H4e3JvfX0L0vFhq6iy7v0u/oUlYQkDXHz3HzsG9WSFXXBDPyTOjITXI6dN
CU/pej1YGnsz9tQ0Pi1T+ZelQiaJq9RrwCJchlYlGp1qI4I+pgqBs01heLuQxokQQCvw/xQyXNMG
lFf3vEx5yGgu+ACgJwbnj6PWbfEByq1P
`pragma protect end_protected
