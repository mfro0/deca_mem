// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:50 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TUgeGgXnSf+G0u0Ho3K7+CIbBpbRwF4/TFJIvTbbDKY3VgmawKkzf3sI5ReWYLYR
xWe2D2GjxJ6W4opiqcSOF5Y3/iPTq7clx7z4vb3EjOKL81jgJk0layzWTkgeRxBw
Yw3zfGiH/3JY0fNzFkXq0yKmgbUnvuahqWsb7r/eHyM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3456)
WrGisCQWPd+unDx/VpL+5XpMTKJMz6cvr+NYG66NE3AAZnPnaVuiU5O3UgbBDNoU
fqYJ5x8fV1Xg48/wGyVgNyffojS5ZIpxubyXYdVlC5ZDu2Xat/4p+WGKqu7PpqAU
dU/w962tSbm7m04l/bZ0piPnXxQ1LSkm+PAyB9Pm90YMOfEjOcZO0QewOXDNDDnV
Li9nfbFVTlFnLWQiXyPyurTOlc/NguB2han0iaixZ+5AnJqwjp2rp7A2lMxBLF6f
R0zavDvOC2K+YTgAIGxTHQJ0lKcMvnwUG9XPLzuztrrknugjKafBohxUnB844kMa
x6CKevtN97yhKAN4TeK9cHLpuF9y12A1PGybW6C+3pg4x9tJkRrqYNDOXKbc0F8i
WNRxQbnpMxl/9gu4D1GWKZ0lQkmWZrDbQb1sxQkf9a9v7sLcU0QgfhQm2pMIticA
JhrK/t2sf3me7dCbFheu+QDXpljrUGisQC5c1Pv2Qa/UhQlTL7bP/rMDLgrTaVuT
5vOZm1xvC4YKOyouaEdYXbOwxoQ7LoNdINPsk4KdAs82mX4pPn0Gno4DuTGBlBFI
smeAs0HQXUf02vh+J+3/iM/8Qeq5ZegujgwEmD767EMPWRk3jqaG1qjd1mzzW9mO
rXcBrR+BQQjZdQ+4Rblj3cqrKvH20BLr033Gkg0MAQwyfoZOvnKUVFOH22jIjPMK
o9nW4M2Iy0+hWMhudyIlfGYK8OgunPn9yk890ZylfX9yYQl8Uwm+tmWeC03PRGos
erafTmlqmjB+DOokOnqXOZZP3mDe3g3Xt+mrsL08RwVSyHXa0Qey8DrhnKXEKzRU
q2OaP8x1eEWng8z3rHA3R9O25hFyywbF0FlcE9nddeEqvwDLitPJvQYmA1XR5Qrq
Az44hUtp661mse2pR+AqndqtOqcHmW+1Np+uII8hxN3rh4G/s+ydJnBf1oGAfNBK
WImx78YLSH2X+JV7OKkmjG4b7oay5dM8H+NlvFHKldFgOE8+z5szKKH4L7xOdHkg
iQmOGVgCg/Ulon2LYivmQApGMzAxfIVj6DwJo7C44vDeZ/YlUNKGMN4XmPNUGLn7
xhXKv8OSqq57XABkk0lZnTWzUE6WXwGl5NE2/03MyRZjXtey6UnA4bRXLWEsovQ2
obmAEzZy++Tvb1hKWqltfpXZrRhrFU3GSHbShuzTgswL1IN3Rd9NqIvTBELwiTNH
fPrS3IyUnwAPfcjHcPev8tgSNQHJWTIEEAW3DT3B+ERSVWg1qIhQlAjzhXFyW0cP
WpFrosXR4643ww0l8PqyUT7AsCyQozn4P25KsonO1l8fVWiLCdYJVku7cIV1Vold
cb/s0LT6+gZMLbEb5JEuqHzvF4ATshEGT8uRM0umEIG4aYyvXO8n17ZWc5zFOwm2
flOwljKNt4LYjoyCBqpzwxJ1agXtnH8EPXrD3HjriFIGKw+GXvHqzYjddZoHj1jL
RLk9yvQShkdsNQFChiQ0dh2gNLbCvIliabA1ItGNnmYT5zgz4u4z3B7qJSwYXIWM
znYvzPBAipZjrZOUtb//xaFNOtyK1KrrrXj2vJUUXVAPjFf2/wwkry/un19c3s85
XlwfWMHQF9zH1hzHdsUSHOt63hmyDL7TbfqM+9BSLe9V84g5YKm+hf506mX0ndIa
LertCiw+ktZSV+IG7j2iBM3brT2joTuVQhpCJ6fl6Bt8/vnjFz2NT8YNneafDOmh
FDPhwjOGxiUZUSDbDAOLhSEGRh5iXE/io0H4HRCGP0HHIQu0F8Vr26zBQbOB0xi8
TALGd7g9pzO0qM5gEyI1BdKIjL+3LulneTr7h+zLR8tY7IphuH2R+4pdr6Di347h
yYztJjm9eSOgiOF5OeUZgNYtmmaTAqXZ4IydGCJqlnb4MxLYBX97f+LmeDpYiWA5
zXD0pQF9JxL7l7U3izmfYolkfEPq64Rhkmv9uvIL9WpVNLqtaQ7HtgtALDTgOHhd
G8KYi/iGeMUVM6dDDWwu0Yk1gYWh79PwTAjaD6oVXGbuF9Ektb1gNpsdp6FRijfi
Wufcc241WE5tAdXP/BOgNwcMKVY77HqSTLZYZDXijXLU6m/dlZ0F74/v+FowDMyz
fo1lemYNXxj0JbLFz6hS1hQN6cMnvA/V0pyON1oGlMEkuaQ+5B3ptFCou5Ue+GmW
B20u4FKiFrZpMAdr+tLirQ3LX+iGAYtDgi6jfnJQm6D4fhjnxjoFszpzcGADSrX3
onuQs1mtSmpJL9uz7aBU41u0Gxm/MkxXrnvYIyhfGzZXA53frYR8z2pq7Y5aYf9T
zKEykMrtRrkf7o5JII447CGkA0tJtELklOtunN8AcNp+Ymmb8IhkTWAiBzG1GSC/
4L2XXKzcStA5rj/T7QRi7GTp7EOsTl9lgwR8ZFjFCI9v3kN1oy/9GoIN4uG4O7Pz
YbNhlqW9ELGVmD4+NtOSpSDuCyJ2aEMSUub1JmuqEYwtzXBYE3VegulOeVK/ITA1
EA25RhKpwl3Md4Ycp6c53gnYkyvHkPMUPErTEPmRddAuYXqfGBXMRru343WnDixz
/wu3B/fv8pXsFVvZU+JNVC/DaEvvntCeV6LDfq92Yz7VP94By6txkupUhWpra/Go
1H84FQgo59/yo85h5gvq4dqcW3FcSzoZQ0FFoa4+/LYUcqukfjV+2lLafZp/o+mU
2+FcTGD72mYDaNDw7ccWouh68sX3FIWCeaPqwCAgizGpJI+off+E2FVzsXC1mgAv
2TmbkoKKGJvie2K7WLcB+1oLdQLJXTbAea+V6esAm0eR28joBRYz3X0uT07HBghv
pvkGg0SMB10vv0PmWjZcJlz2lhfOXoffqxbMN0iJjHjFgcoU99TvXr8rDi4E3VhH
Nn2+u1nrPOcbk6F6X86DgH/Y8o5EwDX8+p/BBRgXR3GyzsULUT9rgjTh8PZohaaI
sA3Py3p9MpGLwm7iGTdKs/CYWxIpIRxz+Q6cbhiEQojmYhuxfTN27QA6lmLc4zMj
MXQiTmvYrdel5VI4zeg0BUz0GOqQvuRaV8oEwJfXphspKRPKcLgGxm8Bd+KNUrzU
fsMZBxM2YSD5lNLCfMgnAHOz8LTFIdQ2JxiM8jG18EJnkA7wBCNt2hpS+EL1DKND
sr2Ifqvbv3M2F8LmHxT5NreOA51wkuEOV9eivUx5kfWCRby/jPGE5aoR0BSC93G6
to87nQ3p0e9OsqqPhXqZ/S4h6tAQzuSDXbEgqL6KDow0EqtymwvRODKoxeW3jQQH
ipr7aQUnOae8qbD5dr+bgesY3BlTJHpwJVIS070/K9WW3S92H+tb3JBQ/qdUSdGK
bRQQwtsghZhS9EqsfrVpyPtyJnD3D6RBTY38MVqrYwp59xXfWou/uJTFOPrm/EXi
cJtYmhLPRn8gbNsg7gfUBdTcmMa+kXgtyroRhl3VYSc2MkFLFFJyXNzd7yt3Pe4/
HlRCaOT4927K2Ggi44nXpQV6BWXbY3kmP3uMj0etXTT4kInXllkA8bCm72e0yT/H
LgcHn928ZNdRxnzsr5uF4Lpv+vIyLxLcMxhWJVlL5szN+sbKdND8+wrB/fpK4CY2
kFZ0wiTl4a605Anq0v4zum1BLtut672n9I836CBhJlFoL+98MOHIG5Qc5s+Aob8D
F8XUXxa1Eo5I8klW8Ihl98oiDVdRewc0Pdjdo3uKlXpbPYMWbmfcEADbLSnvm41H
d67Y3W74Xgl7no2oPN84APXNwGRx5zBOvAQDX6SWN5x0ZdCzys6qgy9rNmXLg4BL
l0J8THxqA1xvb8n6Xn/fe3qe3rm9VISc1DT1LbHycPk2ZjazG7u3ulX9/lpdkxGD
0o7Lvj1y6TZEKlg3hMBGga/+S4yO0IoNh1BOc1wV8vUX9VUbG8vDukzCM55CmnG7
UIzM1v+4OHl/h8cQy2jRYfHOaDyufaUO7UhhQfp2yG6ngj4ms65UeffAtEqhvR3r
UVm999G7SK+Lsl6HqHwLDN7/v+9Fhv1eCdE9PV2/IAytZBKl0OfbgLmSsDEltCtD
9eCLiC0/KfNqV37gSB19Aa/XJI3qXX5PxxkXcrzPzJZAqslNHdZdLWfSosxMS8iq
Qt6N7MXzXU0nv8LczGoRs+i4MD+PYLYIAsVEMh9JNJfKKu4hIRi24zOovzXKwryc
zck8NssMU7L48X3S+B191mvR091pNpLJaYbwglO28HAqQtKIVO/OIKNTIdugUYGM
CwaiFII+za7Ayj6P9Zm1vXgLn2HW7r+/olAgtf3UXWSr/vYEHPbRTDOEkj4hZpG+
KvIDxXA2BueauCZuaBleb8tTNXvsIBjoI1qObwGPOkaH31CSBVd2AcP2oLs0Df2o
MrtyAVsmCyLKslkPggxuj7pRiHP7JuMmRipNhUZ7N/DA+yKs+vZEoadWLk1aBIqX
f+8iKGq9nk+YFiGJNFHvL2Rp3qKkeedgt6R2EMukza5VIS/+m7MLUQgmJ8QmR6zO
XsyRntDalgsZ3diyeEFDwIgAjSgPLNYDleyEYFEPWrkamvKXcJa0b3EDZNBXS/2i
2YX9vbqbevkxmoPLxpS0JvGKvvoLqWnNuVQ1BRF35g/Su/1uJHEkdeY50OJJczq6
`pragma protect end_protected
