// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:13 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QcRfd9P2x5X0wo/vuPsQRdXo824M4q/RfBzyQcecoOJC/d0FWzCL5EYYju70IpYn
8gKYlV5NYmqtuL5X+9yiwaLOZw3Xn82sTVmwKD4L8ki5pvHauB/k9Ybl1n16yTsU
JgKbQH8Mw41ZerMQ0xcWyMPwfczWkE0OKtTC/f2IC00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16976)
eqNHYdApmj87XFiBB63vPPIXhwGNeg3rkMD/7zGcz+Rv2qiB8i4v76uT+Jmv2D+a
v+gTOu3QsQomZpQT1otUanBbjJdOsgWtYMJO/eEO+BqXwhv7d9Qqp5kt079bz9JL
AlO0lvOByMB03KQDuzzpveMF1lkBllHK4CPO7FY3fEbEd81ZhuCEMIjRE2+58ELO
+mKWJ2H+M4rZL+wJ6dz3Ak7O7hWiXraxDH17Nzix50fBVkQHol8tnuS73CsNaaDZ
ScCAdsAadotynOrzcyoGufDzykwLqVgqTRRJozJfm8fIbgZSDg31Zu/cBgqYQscb
RTQO/eIml2UHeLQHjxXxtTgRmj4pe/zWDb3MHV95wTZauMykj7pENsLCDXiA7mad
fUrz90p8T2qEg8zUOwaT9FpRFJM/JPulQfufYG7I7ZJMavwg2icwkdNCmsuToLuO
gGAdcaXWneGKwmTwrjKsCRwT+amAJgSn/z/xpUvdayVRkISEk0FK7pijm64108EK
D0gUqKUWdcBhQRr60ThX3GH14PYmGADXPfyDfc4A9ufRgeky2vzejV1v2Kb2zI1m
dA/k4HZcV/0oxZ8HpiBLBsXFH1j6UlENVtBjVPCdgKnR8hfSaBJjFFiu3lAJwZ6V
m4+t6a/VFAHE83uwFt5loGfG/4ZS8OV0gEZqF6M8WJjf3m+uCkrLfANmOuiGTqj/
nPuCLROu2cybH6vPf3qiQIY4Ox0KK1qKA8i8Uu3np0QdsOua9yVLPMVdBMNITscT
lBJagi77b0LLZrzlF5mIHql64rsHOGzplpf75eXlllcc+RatVXiKjqUsWMRX7VOI
Swq7/RrYsrfuJWCuKeYGF+G3LXPJwNzM7HwHuKWHkPXDzqkmm6bxJ+lJ+Qpl4EgA
9cuCo6DzZBSOtgqvtY6sdds3mGOOLKtZJtoM+Uc+AIPtxufwZi++ltt7Q0N1P1Us
GGZoBRFSEAdjyE9zF2XCAGVM8FSnDEDqINIKkqzT4+KawMcJztfya+6nfL8uzgwG
afyhMleTDiosU2PkTccz4K4XIiDluFk+iHb6rPxurMS8NQcqLBIaMgW05ZWZKY+6
LBgApWJhUMKpIgYzyIH6iEwT+80Tz91oBEfbmaH7/R4S5Sxa67orcU6Gskw3iF9k
xbGk4KB8Q+WhU10bYmrrnGOHj+7Sg4xhBxAvNKl9Xr5up3UaQgra7eWdGLrWNJF+
Q8S7HcZ9yh3X59a77eyqyqd20RSksm3yAcoKyezYEre2IerN4+Uvm87SKD3EW8f1
01sMgaciGyki7dxyW8lefEFDCGAFHK/FO52vAzrt5Tpy3NqhISuE0Ohm5ro3gWPV
Vc4PXxBK0LIWsdQVNO040oh+yddsGZAYOQ+0BlSNlcxyz9SKXwZ+x4cjws3GGvlB
58qEeM8cE2ZGwdVhf8WK2pcWt+IlQOebxJURV09/MRVW4SPI6B4fGkqGtO0HA0fL
JVvKkS3dJ3Jh4qTR2EmmxAtwRQJG8zcaBqj073wESwd3/vlA2G/UiN95ZgGGudyP
uFbz12vgNk53Mnh9j6bwxDE5C/+agZ5yY55xEU97RY9ApmZhPRRykRz3JJdjclFN
i/Zxh3CNtdJcm/6iSblyewkKL6OsEuQCh1EYZPEpcjkL4KzQDCc12VrX4f02RAeg
FTr0uvAnTXTibFsbTXds8UOnJGtF6Rbo4afdkBitfKUSAUnmnhUuvoWINVnMZyF7
p3tfUfAekYZ3uzvDBtENgpWjGGPfTRC6lWce7dfcnFduo+R91FaFci51r48Ty9fB
2nuNMCyek8NSmj7KICEy0yr2TgZtYdeU2ZChwzsf6tVGkz0fQys7K9sNK+Ohb3db
nX9eQibwcD0CHYZOMfRBXL8x6wQcaKOWnBD8ndW462ZvRd9mjIyMd1edqFj2c0M9
+/dXSxNHuOFH4geggjVBWYDegU3R9CWnm9habWXN9qZqFQ3aak7kim8TbyKJDp/b
KMX0W2NVjxplDCl41Yu+V1wupZzY/LHHzi8cY61jvGX/JFYRVTzrFry0XTMLRvHm
Nqgx6UuaX8WIBOe+Y/ujYhL3W/IcoxZRn+0QlZpx+cv3pYx8FN+Jx446bi3WJurM
6DjTeJp9XFUVrQ7/ALyYbusPWWr6G/iaNZn8lndYdEuMWZFJkXWVcQ9LATEKA+kX
2V6ZyvdFGzGBTayKSL/YeCHrALxY3pUytlrImRgzl7WZsAk+OQPO79lZbavNTfcR
SWiHRkHahHz4SwxEQBoN3tPZDioidP/3jQNhSoqzjr+74cbz1O5dJJsFK9YkS6+8
0Z9SiQ5M0AvWwzP0urp7JvcwgctR3peH211QMm6xEx65v3Z+ipairvFoO0Wt3WE3
HIDxfpnamdE9705AHqTfpYuAMBmrqPkhmnT2cErC9p0KLt8QskkZeTZM0ihXYh94
Tnje3eCrdBsYA7onPBeqiQcggr4ZfAe0/e0rNdB1C/Fu9YyWklmhOOhrDaC+IXIM
76/Tyl3eldI3L0zn8nP42yETBjE7AqAFLiYiLdCuyrTIXN9UEsItwU57o0qfPANe
dc4V6bOz2q3l3Qowl+Byz59I8/lgHhPv8dvmcPXscrwLFvQVt5IRrze0TpR9kERk
zK8DYHPoDCZN8IrdGTkzOrLnx7Dph9yDx00bQx2/aXUiMV5jnmzoTYK23i+HwJmi
GHLCI/wOlAHmHIETO36yt2058kdtFx904NI8OG2zPm8IsRwXqKCfBmR7ZlkLbYON
LIMHDbSbKHdzYpWu7NwdQ1PmnSacV471wy8ebVKPElP9q9aFxOYBfP9mGRw87vFE
9eljQ3GflTJakBxnruILp4PCAPN4ELvw6frot6JV8gVcngLqVQ7H1yDuf4BB9uoW
dEGWkMQKYkzFaRNWoeByLpLE9MBzMxfk6rIxR/ZyeUAX58ho3iM+nB5nA5uCr4IZ
+Xb8lDr5XgxnsKdhLKeCMEAuOYOc3/J5CZBM/Y1XasZpew4xqogCCk1XlfgKHreW
Svz//ykED6rdqeP28a0S9jWN2H5oMdQe3CmssL7N2wlqK/owb+c5H56LLJgk0ygo
q81CZnZ8g/IBg2ZHXqW+CO23ak1gcqug+c6ebFEmySjs+AHOPg008ahcLXfou0qW
Br0PwPaL1VBkNkmrOvjv4GCMnLSFpi5eHXINpDiAcnYCEgn8yTU/no8MiPt6R2Ld
cVveu3thh1GkTktTIV89pxjVFV7gi/NFmm1i4PwF3Z57eSFGonWJNP/CKxcDc5o7
cI7klH64SMRFBy2HtMz6xzZe9rYhMCsvmSjloYQ3jxgASRBZrVLljQzNPjO87DmX
ncIYAlFFga77K2/XhKuCrLAFQrHfzqdJJgDfVNWW7t7HjBvZuE1iQpavidiH6GRX
agcUpd0zzCJE5aj1TOeOeuhch7HdI4OCtE4KrNI9VDHfYG5mdvzD0RrQQ7N9CTv1
4/lPzdNCI7htyIiMdqEvWi/q9JK2WLzYr+kl3QwXvV2nAxX1bwXxp4viPLBrUwNt
lcizgKk3V0aTjBu4tMdTC3PFQy80gtZM13/Fx6ChrKRVlV6pqDf3pNbvzA/yJERN
XDhmeQ/2y1S9Xk5BzCa3jj9mqcYkNPLTmeRV1NYS0SMLW4hPIHHR86DUtrxXad/s
SsCHgAPxe+IFnXmOxllAwwZo1yRVDoVdcm2y4vF6ZHxp0htCejDke62HIlZAKyZw
6FlbFGDu2alszteNiUbzXl6UTFama7qXZiPQvuDZP8rBvkGi9ga2rGTNEA7YYr9R
6Gp8BCG3qiNx4E6fXooOqW8oUhbZMGdH5bVxuy/tbkhrxRMPCtRIGarT15xKwl2v
Wi5546O/Of73E7oUbi7yVNaDxjm4vOURygNE/fJMCtrqL4Wf1znlyQPKAqY2QFhx
inUAyOxC84fwn9eBabmCZsy+PvfN6dBM9bFHc2x/o32DFXZ9hVbWkBX6TkzCLr1v
T40jqomCM6VnO6VufNuaoODb8j4nhSqU+zeOi92hRDJNLvlUU6x+uVj8p5h4433+
Vumr8+qCnUkE5QaJSRbyT/pMiyQ17g1TehFE+R2aqM62QGqJGDqnpJRdpnvx7hrg
Z9CZz2y5lLB005PwkqQCEWDibsOiSGOukFHv0HVwRkJ24EpYcuwuCJ8PAEMAMmHo
PtMMiQPQ+NrmOmp33hE4fUxjiYmEYTjJ+FIBX0POMvgRBBsnDii/y2HlKgdp8X3O
ZPycHJI7bRAD7oe/2OFyX6HpJr6PDRIaYWecORJBiR9Sn6HsZrqSbRlf4HJLfBDP
IXLIQZySHIdu9Jb9pITQwBJwiweMPctLsp876MtsWwdeEIvc5wAemWvZrZxhBB3O
rKoNZLfqY4Zdt9TXQMWGsKDSx8hf8zDJXMJ429PtG/kamRqYAyqUW5KyBVdVIq2a
FlL6/a46uHOYX658Ndt2mkcnHkuOgsY8Jc3H9fh7cgzwcKkDWM1RKFoQVZ771IFe
YFyAnF7VtS+yc0oDkwKiz8AbZe6gb4JMG7gadUNc13SdCkbdePCidaB4RiUzI0Gr
HbxF63adm/bWUZj/7Jr+4SYBa622gteGdNcUU2bJbzTCxMAm/lP6A747nA+W7fCQ
LjpEj09eT2Tc8wsj0HOTXbltGauUsCWBIOAgC2VuwvhLiFLCX18Nw8DizHBLkyT1
AO7SMDkA3skEjyt4gMJ455kbdJZzHpGzRiZIuJ0x++u0wQ/ti/LQE/atZ8tXZtCL
iNeotglTWGW/AKe0oGgq1kaokBZGB4K5aSqv1+yg3ArQSZTAbJ15DDKljFSIya00
rWYGyiaXzunKZiTXDPsY4398kxyyiXMlPLKuj5ZwKJ1zkbFVw2Y/YlF+nPBRCPeM
mxRU3KUKTi24N5BG21fCp9oc/AQJxD80VOvtpOj4d/PTyb+3oUKoE0mkZuACxf/N
fqOrKw3Z5SGEN0qb8dz2QcytkG0SbXn4vPhP3uqt7t4lgjJ9nbY0McrgIRgH00iC
t9UPFneYhEktaSAu4ea47YpGO1jaRTBJELgjWkPmqfhh587paH3opwK1T01GM7ff
zaiiYaSLp1YMbmr0trNNs68srkxhNvtD8zYeBZ8eUiyi0GvTMOQhCIHhaYBjrdVV
7ZFC76EXM6VRnRGOB6WnL2Ji06OU17CBNnophjDr1upM/zNycyL73S4aK7+I1axj
ML91nqhlOeE5ShpmsFiKGNK+MtNFUj3QY4eorL1ZLHG7qyK2L04reQCdM+uYeX6X
9o2lSdEwbkyGWE6i58uSOE+7SxHwQ1RqxElTE2qft8hLh0xVcuO/gWFuUt9Iq/if
valGnpJmfbvhMSDATC56JhXw+kBB9SPVxL6uHQRPmMj7qXFgi4u9rOxeRnyAfxIZ
xAR/uQQg+kLE3vZjkZaxvfl3DeYEpdHyH/a32svi3bJpP31HryhSHU6CddIrf5Da
2/scyJBffm8tkIlFBjWFYBVqUbvk4JQP5GIBWTskwk+PzfnO6upkMmc148qMQW9J
quxsJ7yNMPwtYtoGh81JEO3ok4yAHZRkuIdBn8MJ4MWo9/EJFrP8/lxEBcuRFcaU
EPqPJUcSYWZEekblsSsARNrNRbxCENqeH//Xx9nq5EDf5pdDBP16CSdS+rvtrluo
8SEU9KZ30aZbru+Riby+isuwzVKYFJAK/z6Su1rEOhyhEKXfTtEIWYKIsb86xMBZ
YE0qK8Yt+Gr+8Vuq1CAy8wx9bLsckaI9SfKNosAJyPbOpKvvHkwpjT6d1ODuia+8
MHUvaSeOGTyZBAoe1K6CYQna6YIpw3oGO8KLfQHlZybHvk0eQmfT7ggP75xWwrkQ
lW+IBWw8R7ttRVjUE4i6A7xmZ3SC6xp51LYf2jYpLEOmIOV22cr2EiBhQP3ch6fU
K46wqG5WpRzp51pb2g91qvND/6KFje9Q5KvFzT/qJq3xSRbss6WuoHVyTZbMnTQH
687qd5cLv2ZDgn+SN7071QlzsgBwXKV9YEoNVGpKl+hXYTlvt3/3syzfmukDdnKB
bEy2WVFK6RrF+QTloS4LpCTiM7G5d1re14pIK5+zsOKPh4faWc/VOc3KkHrfQfWr
Jg9M11V6PRn22q8BvbEvAH78TC1p4hgfF7OvKnEpbx6gU2P/V6juzAHO1T3LV1lU
6zGxBjnQ+kYFFZE/2Gs/aA+ezvru4+lUVZOpAfyo/NUQ7Y0eT00lUXVHXCXs1bFq
vNcmQ3oSvh0t2chuW8EnmMd25hQX2/PCj+Vn0Dm1ld53lSMlFQ4AeG0rVMvqQ8q1
j28dWs0koUxNftFtXsbQMNa2bFalUl5bpq4rMJESf6mD56oQfLbNPeASfbqb1KOQ
pk5O56lurjqpbzoCERzqDiDydIjJDBAd7tipBYMMRn5tw73Swtf6YpjCHqB9gL1M
2Y25D2hT2sYSw8TS8+megBnk1lte5MS7FJe9rA2dyiS6G+Ong/tIDXuKjhYbzWbJ
7UkHFyb2LsAZs4Tr1pdW2C+QbIHwC6P+haRHCcm8vq13dekTyl+m/JTChY7E3iJq
ikbOWgS9Tmuge4uafHMxpuTY44tP/6uTQS4Y9x8BSefjtXhpGUJ/HhGuz0R2y9FL
IoN9ey/K0uV62+2kZiSJmklzo3hy+l/6Z4NkYv2yyZcqtjdhaUOISEfZbXqd2RRo
Rb2b/Xdoej76wX1uSj/vChr0S+S/HEj5vNc5Bu+uRMfCsbCrYRz5P77FgPB9Zu4v
6WW9bYdGrHWA24ygD17rDjImavZe2Wexopdzxt8/G/tVhCXURrFF3tMZhYspp9D6
i2RyYhm2HZfu9/3WR5IB6QjRxVI6iCH2vg79RFhzUsC+ZcJxF/V+VKbaNJ/dw/f5
a/KChmr0ukDKVniWGNFs6VXlEZfk0gZ7tOaZKjRlbkzrC28LATwh0EsIBqD6eh1O
DzL+LbUyoSuNn8O9s13Y2+4ajgApM++pe9wctcy4hGaMHFCy1Sy8Mtcyt4pcjhE1
NUigq3DdLyIWz3cTvO7BbCty0NRK92A1Hc/oJyonoYbcrH5CYSNhz2UDEspH8nwi
eQIc2JqOWHXqOOLGBSd5e/d6eCV38n9yzO2t52MIn+lWddzFeFMw7hlVruq/ejoe
pIyeijdX2mWAWng4BDJnVY9uwFwYRX214HmHMJmbivfz6Idpy/1dD1cFRn6qBOfb
1ftY3yqqzd2RonEc1mU8yqYXA03BQ91/2VkbtBl5W5nl1m9qvpuvvTXzr6/RrlT4
3OW2wN4WM8mPt1pAld0+gXAhuKJf24W7A5TuWNj7PRy8hn8ASzhra2n7bkGSyHG2
QMG2Fv5UhMBA9B5eYGX4ppdrC28ibfJs8S7ub76aTOQfzkITOOfzOkDOWEI5xTRZ
LMlNl3aiYSDbEo5XY/3X9yacoZ45lm4wQIJEhGzr6IpLc+oTTcxZkBdblyztadAZ
Dsu7zjJEBSqoozxbRO0nYliFLhvRhY/tscrKKObeRhDKxeRseZUSFTEv1okwHvjC
yHm7QMBmaqG77P7JSmZW0f0eQFqAACLXGpPPCBE4AooweAN0aH7uaKEhx65ewDLc
c2o+ufgup/l0wyr4Xgw5ZskKxe4kAg4AqjYkNk3KJfax2FVCAOlBNdy7YKXkaK/9
be3KT15swkWd/hhetgL4a6lqhhkQNH41WHZI70hTf+8kkOhQ/J3ikG7goi8GxkuH
mDP9nzvClsGHO8ytiSBaxm1W6Ejb9rz1HsNRpFgiwQU+lWB7jRAaBfhT5cuvIc3D
TVEGUdzp/GRmi4ISbHh2JT9bmU8NCLANbT3IOKCuIQRvlP53xMg7OOxbwGhxajgg
UHa3M+Mw+IDMeboBqNSHlOGbc3pSBQWeY7bbSMZpFonSAmUg5mcTrAgdWBNbPDv6
gt+0Naxs3H85WMsWUkvzrrnhL8pwoi6nJy7lHp3NPpLb1cmgRWSOqviHrvcWTv+i
xTOH+VypWs/2dmUDBZHVN1CSxs5McVrtjreSBUD5cuyX1Jllq6G2ISL0xUWzfqQW
XTYwCnkmZHYy5f48rJPeonbjRkz83OQoO4hd69GElbKp8tGDWoJrbwjsx5/WnvtT
tossGWKpedTeCtuQwA1D/5fuw9N8G4+an96rZ5U5qXVRBq7QlEnbAGpNL+Oy83ey
yzA4OSxFb84haL5wFo5p12wSiGiYkUpvDnivtKUqaXyoynV1LOat0RXypjxmsN4P
nvhx1b8MpQqKsCT9J21/okNwVTVXZ4jV4pCCKGutapKf2N+9MOiRIA36Q8zcuIhl
EYl42ziDCaH7XF7MRmMMTCzCL+5hgufU/SP/1n9iSzX6ngDn+ZwpcvfrSdKJ5nsS
hMx4aYyI5RYEw0DXFNmghVhuK6yO7a0IHDV0ppzzoGt/5gaz45Oi9HFC+BrHr+8m
XqmAY5gDqZL6JcgStI+CiAr6WrromLa9ttd9XHCoRAW7+cg0vN0zuNBQ1+nLlYou
cSl3OF5rgK0uY/SMHCcT1BckHjo5ksfjHcv7Oqch0PWuxEw1XYZJ9yHf21IOH5lv
CAhWzS3ihHrm+xCUVGq0fAdWREOkBMfiRlU9SIQi1bbVexPXc4crgd0pMideVOU7
lpMRYp/UQAc/aO0i4Z2s2hUsIiUlRMG+jGicGQVEVIFKDm2vuFynIHgk3gGI6uI5
8XHFgO3+Di9574OX8EcIaefUtNdLCDUOXqd3SeVaIbgqa15WD2XUW+EncVYr1BQ7
9kCE1PBXie3g8N3PtJK1rxi0QeCXXAT0ylahCpbzfrVlu9Jnpqmn9/hIvmTt6y3r
bLVCtRmDUpEwXnz+Rh8CeMk9lBPb6glkGWnLWF/Lds77SE3Vfv8YkDGJ0mIAyUNB
SC/3nw5xiuXXQ4dkiYtte8/u9CMj9OYYfm97k/akGY59qQMe5bp3Nu3SXKzo2p1A
MlT7WoUQHDj0k28sFLeS+99Xt54NZ+6NLesdG4Pz+bXxRa8z7XXm8xyVTLXIo1YL
t674e/HYCCoPOI09sOOCd2wifP4U5Mc9/+sTUWd9Sg5KilSE8+Z9cDnoIRLDUycH
w2Uz22Kyh6oJc2yh1zTqLepMRQzTbw8JvLDL+6H7jdvi15GsnWOQ6X6hTw0c7LeC
vlJEJI3Yja/sNZKVxgAE+0K3OCUwv5jNnzcuFpa5yeeiPEi5/w747D8agUkbdDoi
JAf2/2eV51YV6aJWNGR4wed6ug/Q/3ZNWhMc90n3gbKu6GhRth/o0Qvjbhw3w9fQ
+ZjokgtwYwe1kQYykfg1vxYcxUchAfrc670uPnbS67YttcCLNKF0KxAK5OTqcWjv
lb0uYCvDOMlvdR34Hxk/NhCNQdHSLkHufsSMIlQUw5jif8dLoUO2An7XIt8bSrrk
LBgscijsGtPJeiFRaydGW4UZTXWhcMyKgcci9nx2fSAu/Q7BPhniJrQpwWSS0txC
AWhMUgtg+He2QBRMmAFzwaqPhEwQxNI2ScBcqPCd8c4DjsLtf08398gymRwX6NRn
ylfaEpe9pwXwUd5cUWgGbrcM7GMS4m2US8Jc2NfHddNlgZqmq/Dre2jsmACQ0iB/
dWKgn0JzWUiNOIwh3Y6upJQrCJHsDWxZVa8Q7TGTTyFv0W9by1WmzpD7BgYJTJQ3
npHCXK0smmoKV2uOI6l/JfrzTvznbsuAHoqhZ+yU5YmQoByoeRuLt3eLtqYIgtmN
m+OcavQY7KrPLyz9jnbtsnFd8cN+fb88SBpRHeVgD46qAbEaVlc1iq5ylq7MYdgh
SmueqrcOo/CA2Sn71E60Dq50wi4MjpqPVO2vXgRzolD4g4/KB8oMcr2JYNJ5Yej/
6+5gtodOLtCmguL7Bp4MvJx+Y59qrgtjtSXXcwRb2kCYT6YaJFUW27aBuKBlWjko
TQ7un0N3E3L2qfXuB/laqzKOrUZEKytkqi48b9ExQW/s2uNbw7gisstt+P2hJA+c
r2InWRC57jbQFeDZ/Mj/yXTwMtZyLzSnYtlks1wFYo90qOQyyF2qgRJsChwFLQbj
QINps1z1Jsvbn7qejdLM41rzhWvh9n3z1eiuyJwbBRv2Qi+msLqSJVhOAijwf3X0
yN80CueaVzDkz0u8uCfDznU9dXjjYXFcFyGU9MRS6SieveHlWWgwS0kDDbUIL/Qd
+92PiA0I3Np+8mFR1BsaLLvBrHo7XkPptyVYOLK3M7ciJVligXRr+jqEs4bW2szH
JisAwZFpcYwVjJH2HUlzkkrJRyn2EoA5hCMqMjT7SlphYc8tUfjaCwsl5pIYt+DD
QES5XKLaxCqKFnRMe8nQTJNbBym0pJqTzWTL4DXl6CA/3zIYCi3Na4YNa8sTeqdi
a+c/RGCMv+Ji0y7fFMTX8jrYB6twQWUsg4yxnzn+BwE4cEKYJerPrl45hPJr0zoN
BCFn58Vz1sVHc36ui65GSL/EcmJO4iq6hhj/N0nkkcnYa6Q2tQb+fEPpHs8AmQDN
wMW/OGPJK4dmQWVRlV0ZTe5P7/U2Jk/sbqOf2hE/330QgvbnKxqhONcOa5AsP/RT
5hhCiSZGS/PM2JjKH+UxbFWecEh2QgKQm4LgW3Tr+c2MaoDqrtpQTY1+i4pJdCZv
BZNgxT1/g0YvSlQe9ZzREkXtwHOKiOPLPwcLMOOLZAG/6jdI/Y/CKPZkcNRvn0dZ
vbzvL387Z6ZHZwE+Z5ob7wfigxbbkKSff830XzpaIlNUBHP4wQu+fL6CdKBkpz1C
puVPbMDS28E/43Co1vhTNsFnZgCHSuJAA2/v2r5aHfscS/tTqx2psVE6G7lgSYXL
b08nu43gHSbhK8VaIBZPCG3OzKP6KZvCVc2x+kGftjxjhtgCTCZpsU0COd7lZzat
j/WYy0KVg6uUebFBzxh0GgVStxdL4uFZKR5Ipb3SeQtfzvl62bBV4LKLigDZ3aEM
fGVgvZugazdD6PmtWpnz+09olzWVQkQSIMe2+MCyahzy2GCmCmAGaA91e3s3QNQH
AOPs/j+PZBLdgp631nHeVHD2HJqUpT5fZU1YadWyZbo8u1OLRckEmmO9PcQss6VX
TaX3LH1/I8YczELrQo+gugyqaSPikhZWPdGFHVBN8DK3P11PMExJDQl1xP+fdY7o
lrypxp0y0ui9pnMXibhaMVoeOGs0Le5ZvIHX13+FWJRF0B4/Re1FgNhckLC/1rRt
vl8nHghQb/BE46t3OtKn85wA15ZOYsT83iBJTxpfmRhi9LgUxTpO0h4LBD7AGd9Y
Cz477WaCoocGS+sCuDNsd02gwbaYRZSgHf9AaEteg5a2UsSZXls1T10SKsx+aIxm
WYco3iHT9Z1G8r9j6zhAI9ZyYpdnE5Z5ddHp11g8ue4BYeG7AVgJe10NpWDzby4k
nK+CY2AkljJWK3Lvr1vnoJ6JOWzx8H+m8np+gIVLa/s43xHnhVhs0QQlMrk+dNBF
A/W60Ja/CrcEAkzsVEuzQQNjXDCGj/Hmu4iPFPAI7pA52PWsJEw3rkkDpfzJ37iC
lCKYjANT/bzeq6CL43o9QsvFez9lPArhCfQz2UV7dyMU2BLyqFuiOO8uzpb89EL8
qGhZU+QnVgOaOiWdo+FWYDQ4mAMK3erL6Kcx4McXF9g2GpbT4UpwjfgesqK2VNJP
Q5+PQN9ve1vl7dcCvknYsKrh8Lmtnemg1HCMJ8cfey4hMWxwjEbFJr+gFQM9O8Hw
5bH+hp9cdaMLG1HlPkX9otZsKPaDyNnJdgk6l5wbyDTbs+ynOepG/+w05wxI/2Kq
rQ5IgbGf5yua7+Z+TkoqIV7VTU8eHNmsc1l6JigTP7WgJdQtLtnvaSdZLGc9RJPd
QECub27bt2WjIdp9ECGgrM5ldWlnHzfNdTfV6g4uWFDGKsShZ3R0jwMROGGPtZoF
p1vrBynLXAk1KnmlJnvNQHNziK4PPpnAQvTEbzM+9BE4k8JqxmRfqYM0bFw2H2WD
nNivVYrUWs7aXPR0+meeB+9kzsd2mqgaYwJaSxSJ4INYKI3KAGnaS/kC8tgvNKRr
CRX/eOpsF8rYS5E4o7eUoVwSKyY8lgHbqOvu9YdsWaYN8s2RYFnx0WlB2BQSWjyh
z0HFlr2eyhyTVhStCq5dvMQCPVxeFvoDPBcRQ7pN0OXBbSLJS5b4bDuRs77wU3io
+EPSjjLqFNv4TyORVBEHYH3hbXFAh1ZQNnwnxmRAOt143Axv2W40cm35sTUtbOky
ERi6vZySy5TZfu7NEN2cmtZNiD6/e49XyAa473Ywympltn1JbSKmUcS5e9PSGGuG
4xa0R125vugt2tcBaiVa/6YKKWC7mVOSTV5KYQH71H0fq4IWpmywx4WlY3t6yZ+H
OrKuOExyWzaGM0t6ijf9qpQmOLpC1F/WMmPfLJG9nRIwhYeGk+Dv6+qn8gDBnJTN
D+bvFlcINJnt4J1l/HFcaQzccOMCK5JjfV7ysRnYdRRHhPA9k/uT4dIpbNnPLv6S
e1cdP6ct79KsG5UFrUgLnCLxtBwtadUaWA8rKjO9XJhjKitKP76htHWgZmYaMsVt
ze9R1f1o7g10oo+MsfOtxAapkuUIojywYrGXejD/GO6UqDuNsBzJS6ArWEgj+c1n
gmQmo1vCgY1Rj9H9nffMViqKTALlJhgtasqwZmTq8E2HC4SrhUUUCMzVE042Xvur
TnuNFRrb35T2Lwr3pmAaKOf91XnMrXYPjlF2n6YIo1zoAqK34K5eELHCvPgL0TBO
98mUUSoTSkk02HPAtL3Z39nhP1hykts61FDOBmV8jZObqno60s3MV6nfE1xpy7DC
dHB1hQW4CuGLDg1+d9gTIUUv0AN1ry12BHVaP78ZY1TQ0c4X6gW5D/iag21EbT6P
Kaa6Wd3Jp3tsowu3sG4xbxDsDCPFCmYrd7PonY0pajtw2kmcrUCZv7/DsO/NNXV+
v96vUxST3K7FcjKM2F5/HwGE9rRxkQRd1TabYjZ6M5sCPfO9B9YAm8/dH2j4IIUc
sjgv+k8EqQw/Q4HsQLWyF065pVYgJQJOllZA9D7uAaGUR1TFq9iTpYyvFJ45eQZe
DbbIGMWy5b+P2RQ78a6uyFjtNTxIoAMesMZy+xUvR7rpv6Twc9BqbyF+hf7YUhdD
jttmsPFVZHommgMitZEo0IUerpxQCPCTkl2HFhlJjExOBX78xyxrUYEnbXG5W3WA
2RkIOtnP4I5JvRdSBWuDoQf9dNS3F0EJkJb+DLHLmnczNK2oijG4YklMOSvmxlq3
06hgseOhWil7Y7tRKMDY8uGzQmfwVQXYLfEhX5Khsztuxj4NtaJxJtfjsT6TZgeS
DDnLK1EdiRFBsFXzrT0n3aLL0d6DODwSJtPsnB75YZYC4q1nHWTzxCYTF5vqmE6r
tllYLybcwo4gUsEmS3UN1Lcq9CsC5aj67i7Jm8ArcardTQuITTV+oWrAvygyUIPC
8zVtyO4rqnUcPxqioZGoZSRsnP3KeG3oXh7SgshjXo+BNGY2tLFRA0a75iNVbcd/
+I6vZvK9FKetnCBKQJLL7NGgjGg1RKSunpYppOE/mBU0z8qrJ/T7ML7pH7ZPRzAu
7P4/iBOg7g6vtTYju9GOKf2EhPi+gXA/LPdi2iOe0I9q/rXdpFjaAoo8Fo2nFrNx
tjf6WjoNdY+UiT0vhlXHPpyGxlwOmP4V2vRSV4IOkHV3BYRMKATGH8y4qBdAyyZo
X6cyWusTPt286f+VwHSB32xlgTAyxUo+YL3Nz4kuMq1KnjZT6OkbaZNOHcoEJYzz
Vs7fVomjRjTtvYbCjUudf3bArz36fEUwjzzD37SKjEU3PwMS30B5xLzuG80XKYeN
WG0az5sildOrTSrw4NyxINyEgP7uRnaA7oLKfdHNCLX56AiyOixPf5m9xT4AjJpb
pvE9cfFQ+5g1/K1n8uU+e+2d6U4DoV3Q5td92vSU5W3hAiMeILxXDttgut1yk8jZ
dmyLS5c5EflgBKHrBeMG+6ALAKi+W9dJINXvlsP8/kwzjhI9caDHyTGHW/wHQZYP
3mob7yAAnrHxawFny7MUYJZImEZfnOvMj+uoeexAo1ZLimMVx+GrYJUwNA5m8dWG
y0a/SGhEzdsLjHQFI/Td58Ly0W6u8Rov04vNbg0mFD8shlxAfy5HLHIfs2uSVjlZ
WiXqWwqEG2jCUfUtO3Q4rxe1AY2pIwtf2zMaPQHPGPAFb7UaP/AER22bMpelnvkm
KxX8GW3+96gVhGfTsOVALtBtX7SRDdSYwwcPLALXYRXTSHkWorCvma+eQ7IxlOZI
/0m0krc0Jikh8ql/USJe1qE2KVwiLtu20klMzCy3I4XuGGwHnHVDok2rIQNIb6Rt
/eWv/z6uX46VjNywTR4Z3hSBdD1FV+fAFD244WFW7DtYSQhZQJLdEQgv0WlOMW+V
5OLe//r3e8toYCA157kF2FEg5X1MXtnrY0a6OS8aCHGajd+oXMcNU1u/DpZ94ySa
e4uW7J+Gs49whnxfjrSZQGKIoZZQ2cYxK3fInm0C21kavgvQvQYBYrs4MXSY7/Ko
k2hDk+AS3dYGMl6L3OYDP0Z10T9ZGLqIGerPYFi2hFhm9v+dJtP/EhirZHhlyeno
XTdUDwGfZnGrX4OYyModTVpJAElO0DukQAvM4ICf2uAhzfxmScELeDWwKqcijJX7
swXmTVvxk5YCqgEQP+G3UUw5DW3HsCVbM/ZK5KiD3Nj/yWND0TSneqxacyA9yYzR
0E0kJBJ92d128tt8nrNxLqTUmolQarxvY47ZDe0ZyrwW4joztkQkD/qk1EY8DVB/
VOxet8FxKFLYVV6daf9lT3QXfl5wxBYMiu7WBHCZWOn0S1P495XXL6ggdHiClG/5
5gbxy/tSWC1M2yy+K4ja9XOhiFnulvN+FExiOt5PEJU1GknpaEWG5jCz3Gi1Edsh
t8EFPAfnCRFIjZPidMNQjg2VaSqGSDnqQAQmOwLzbATuumpms3zmKp6Ocxt9rtnY
TVNZOJgGqNPITjoLTaAeShAR0Ka1mc7PzDRMSEVwbI91T4a28FyxUbaXlgK7cHT8
uX7lLwaR9tq4U5SbWCbD/W+vQvxQ9q+ErFXxKBmaPIH+p6O+gaGUWqoBM8qQRjOi
Kma3e8i3cnWkLr1lsN2DYG/5rQFI3ON5IdyLEyEbRu4Z1tTe2Fdpn25xkWGVQSOC
rQV/btH4ySShLr/95foNps0GEp1lezMlJtW0tsRxtiq9ecxvB3pbSzXMh/02pyXn
ikbhrtHYyzCKBhmgD+wbw20OnGEECZtU/BXyahIiUW3WJ74Ht0PoetN8lbNQ54E3
7gCHEGVOcfdcrtPCUDHzoQ0K7zlQHYJNyZRkm5dRr+eZOgmD2rLxJlG8RTNqaZui
tOnw2WQ8mYdkGclG4zxycziXhD9BwbwxGAF6WRxrWvbRnf65ZlExmyNn8D+plGFw
uA7XY//gWR0Ls/xQCvZoLVSEAf9gptKBJQZ1P7iCnpdyMFGbnIVKCh7mrudx0mlX
a17wU8drRnQo2wA7NOADI3m9b/PvSs84+frrweZjTGifoq+Da/e5BSIkhvtoTI3E
b8yeCo/uniljeTf/TvR+owkvFbIjTugdSmxcbdSRkvZWZnYcG2Ka3lZgk9Y4q9IH
wfNf4b4/Dcj+Z2hjLf++agCIpXBi/A8IoFTznUE/X7vv68O50C98DAdwJ7YDmKAR
xDc+G10BHdpMja5LrZMlF4E12VWLZ0K6rfaMShhbDAZsJuB0r2uDUoTrCLtxGBBb
b54V5sFiBVvGKhAHWUzSxfhr+prQHJTCNbrt/wo5LMB4zRCYwaXoWAQ+iDSLIrQu
iAdZxx8cpv3s8nEf04w1Lgq0IBipYsY/hd8jwwSRiaeuxNUwPscqTpvkSBQtUwOZ
E3SltUApDpErvQBVjmT1FaSDOp/piU+UnDesXiJIn2xDYtVJ+WQ8SP4d5iw9eaaw
A3siGAzn5EE5MUL+4sb7CE1Ltf5XzJrg0apWBEQmPZt4QEYMG5jZnAPmSk4IoaKP
QSg3xUZo98IainlrwMe7gdAO7bghDZJj2Hp9gVa5q/BMM9LU8L/QjQbmcekowXkx
fLKiXgLY7mGeQisQN5MzQh6fHUg9M8LZHlviUS9VCVFgv2K35RyrOrAcoi/16eMm
YcehCBR0A9BTGiB88VBbMNoGKl+JVOmmTmp+2kH+2cYo2hz/YYWoS6/6Qb+xRx3T
f1+TvD/Drad585APNnrZOZJurHpYIkVVXXh0R79uOgfblQvwHmD9JPFXITJVoAZa
qVzqn0bAoMkEJH7cYesi5OJvYLw0JvQGd8VqqZgKkzuvxQ8zLhSzz9OCvYGC0xXE
nFP6G1pobVjg880Qqr0wEXltPFqR+jqKeCb/xk+8fmQzvVPiWjvbaAM9Wq2tPTTY
IaJq6dMoq3vyDETVC6PfNDluqg1i7YfnX6k2tQFzfsJ3gwDcsYMCnZwwP66gQr0B
JW3o68rcYkSsgtY+YgEoPv0pTqcfeq2AQfDR9TuazmsUjFY3r4mxfxVL4OQ7gC/v
58P8IeTbz2U9Cdl8A70Iguro7ZvE3kfMDS3R44elcxssCa0bNwkPnujo2Vj4JKkF
aEKs7v6v0Ez32nq6Gos0pn9FXnhfgQERKX+8l1qDuLnnRGLVGeHTnmRmY+hXnWpR
LBZQb34iPKkcBvJ1E4G1L/Wag/YTGXQ1/WGkla62rRWuySE1bQHevt0Np4EF4eFh
wiHDoCib89ZQDFzYUHwakCFrJ6jD26vKJwp/zdz+c1B8zNvvVZsSVxoX6kWqeIip
h3V3Q8fNnZYUt5TQzOClu4VVi5OYrcNgWSLZa3Drcnxr9Xyl+LTt0g6hDoUyJp59
w73ADdXvoOd2yqMwUL5WKnLv1GoU+W9+hbYL1RcNEz1dH4HN5yiIE+AJGpV60S/L
Z6ggZ6ozMqRWP0Y6n7vXFlHPYJ5kjiTGextHGYxHF3DEKOolys8GjFEXVMAZcx9d
6pB/jeOQPzky4P9XFfEnffPbYe6Z9E8+ni7pHxIjc5kVzfM/oJ8+tI5g/L4K9gfR
dk5/9IXjjrQi0twCwHf6fecZaJZsYswHKLxHy1DzW02Xp2zvdrr+X0cThYHJzpwM
NyZZ5q4EOsLQJDbNUqxo8DbbefOHdKmb98RjFpFHRNLXaugwbhjG3Kjt4BOZ5TuR
L1aray9j7prZ31d7gvWO/k5+5SopXFFCAnX9CgU6dwrz9y9UIflmxpTiJ0Dky05Q
YebQVXkKOQ6Hnu4hzh6RwQeAv0sEj8cMMkxe6CVSwN5Qu8njpWaJj0V07fM/XOPB
PdioSmTx3buiM33donbpddh90ZQn+nwj/p4MSmhpZS2g3WAEVXfvollJoVIbo7Rh
lw33PsWRSgyzUVN45I2Xyhp5hPftphElirmDgvld3Ju8pA4GC/JmRV5xcvs5OLQU
XAxtPx+wnmE1wYUnyz5Xq4K95gAYHaClqvY5i16agCw3aFhpepHP0HH2y0bkJC6K
px668bGXaxxUIH8mp0ic8GFu80//cKzyG31rsAyUGikTErzGwvHSJWpUM79luACC
ZTEsTFq77NGD6xTeTcstlmVZ6AWPCnMFfqnQvaUE68y9onnxg+hbHwiblNbXzSD5
8CjyZr1xDvahpiBjPP4Y3qfyLzLY5Slbj7jCYwBQNxwuCcUJt101VD+POAW81l+o
YUOfADOUB9vLRDi/DLAdTBAdNEK1ZRRRwfBUG6ohkF4a8ShP6qzHePfuMHGOBxmg
a1w57HVmg/F/W2SP2IICdecF7BYpoTCEtsor9ZOWrPr78rj0PtifedXvTGDPHrdZ
fDCl2pTtKE6Kkenl3ztbl1P+D2KRJubXejjXlmUv/lq31FBrr2KtBnO53Byh3vYE
E2iCdgW5AR3SNramYL94PlNjoxdTCP1KJLUXMk6SZW7w/iVr+UxldEIv995s4jCF
W8U+A2VYvOK2vPZqDvrCLOgwXl95iPXdJrzgrqlyo5pAut4oPmtaK8zDWONPQZ4e
rKjbgXX/uurY+2tyWCtB7CZaGZwdol6d/fk118NAO7jWZv/eULe5+m1Mcr1gWswz
eoyx6yCwAKkZPHNHKSA77G6WU5GLJZHOaIO8FCzin6qAgX6OTHmbRvK7iGvzwjAm
JZArA//oJzSMCDT0UHP5YGLeL6xjs7Tjm5zecXOLtMiF4/bqj7KVY+y6OkeuEVCc
gvcM64xpEbw1QseroHjyy1iSthNQ7CbWxNXcnSFy2XpabcLaSZNU6eM9tL4yf9HN
x7hkf3RR+opD7/68UwV/g1UoASgPd7f/oZXsPCdAd9eczE5geghdD1NJ0gbZ6GVx
qS3ytp4wq/IuKJfxugTO0dWDaDl+5QhxCWA9dpkYsgtumJY1pw1gjIRsswFeXjcB
kxfHjNjHlAEbPRbQ17X45Lfbbc/HlPtkzp/yS5XfxMvTEIp4343P/UCdAHKI/A3S
G4X/oYDRTNPapvuvv9DzKfJNxbi9yOHgU8hqCmxjfL1dSb5LwqZS6rnhgtwCMVRC
eutwT9eeKERLwsGtJTlCSlE0ChVpHai+WRryBROxVyntawwP0AYPSu8y4W43w19g
lP0fb16MzPcb9kwcSblsdevnu5YnJGviOzwWX1LfxiUcW6McaFpDeO662zHtO8as
efL7AwCOYwMJkobkN3xrQcBaomTaSh+dx6du87T/f735+qhG+3uZBHRbC5jqyUuV
hYGfXb3F48ofTfPjav7ZGDxJvwQqtqEZ/lcM1FGzLXMN7hDmVC1AdDOtZpt9yoZC
gSrfRt2zbACkltTBWT7XBnEv9BQludv8UIPO9VpFFlKMGGyyYiIpFslCATTv0YEs
PB+bYuGkMs4/9qn0TDkUGRcIdzif/9ZkykZxKfGh1CFsi/dfa6gbId06uEXSSibc
olgeCGBae3paplBJWdu2XUzjdBdDBNv4Xb/dWesa2SZA1d+sRvF0aDzew21M/u+B
KtLuyScpsrZL85xT9CufF4LEwDLWFPUQHuZk89SLj4yDGQBnqP2nSzzRATy2qOb1
d6Ogo7tnel9zQXQDAK6SlrIltmc7G2OUUMHOP2GSz1lFf0eSjJb64oCupTaYVe41
qFjVV0BzXNIohgKfM1YFBczLyzshQ9E+V5pX5dGkD8QJYuCZ/wlxbHqNRJOPD+s6
w/FkCEZU1yeSb4VRpw6DMUdVhL29+wjRV2BTpqaDy+Waf4Trts3eCPcRs3nuzq5S
AdZJeNH6ieyuoAueLnbZNdMbauRl9+u3y4JwtbCyBcmhyJcKz1ln0ef0LicbXnok
zg6px2TepdLDZVqT9yfB6kz3PNE9aqJ5OAt/JgM0K8lCVofjhuOOzestW5z4fxN/
kwQG3R6VjYP6x8U/w0Bf38r2g/unNBQK9+NEPchThco8djrEf/UInmENRO/iZF7P
pAcq52HNmI+uvlmnbjubzu6k6H/FZWbzjzl/cLgllvqTygEueibS8hIjDlrZFGna
NSUb6CkpbS4INLZj3hLX0fBZ/yKGhSQEJJ+moh/K/3Cngtvi0YZkqpCUjZSc9tdD
WgscpWcGAE9yoezfQ6ZFh3gPjUgsD8+fns7CMiLqO00ky3FPL8EHownca6McYhk5
LULdfJrupdUOef3IqOuyEe0ywzoLm4XCQbF2a3iz+LTc8i3FgSFSCV4836w2i8A5
aWnlTnboybT4028NJZ2qsdxCIt4uEKieMTWlynrFN68mjlSJTdsx89SLUNIorBtu
d55TC8QqBtkq3o2UoUtIjmguiFPXzOsejFOT8u5IGmHe39E52Jt5xcsxQV2fjc/1
ELNMHJOC+sCwnIOmXJdGJhEW1mPseCnMOKmxU6NhT7wfV37DSe6EOKGgdM/sfdoo
NtWR8vkRAcG2asBDlW5bA4YA16hz9UahxmpyuiyTDJMAK1/+MdFzQBBHPmd9AhkP
BZOnApwweLc28h2cgODP5Erv+PhVF8pqGQldco/ZsIYPSS23yNo2+cMFr6IdGNZo
Zsq6lW1dqHgo7hNJmSqZHyNFSqLsvj2sjpP19z73nagj3w4g9qN0G76hfrHqoSQH
RIVf1LKbLymtb8LrYJZTc1clpKje6SAiH/heRVzcg+vwTTMHHDYMqvjVQqswo3kP
KaVTPrrh5wG/YVtxrQNFMY5+PLzLl4n1rb7Ir3nQDiahyi/KJ3JXGXKXIt/b4ByA
I/2dBRB9CI01wK4is9ld0TMD/lbxW+Zr8KsuGu/0V8d1MvxycqqcwXenLRVWpLOE
1UNZDJc/Wdlkwx4Ado/40WYzWnGfAN/3fXQ23i4coabzIIt4l5wi/Z0B81TOf0w4
BKKCohfEZH04JNeXWpQp/LPxxPg2S5a+I8l4PQ+flAfbB5gM0FNueRIMbabMxksj
tCQAaPs6BB3EG/n3+gJ31KRYErNx1ImFDRFONZLocA9lJvWkOQRi5reGrKBgQ9i8
KJNzxXi7xZ7407WqUdxD4QkXwtvpuF3b/Zm/hAQzhLkzvCcHK/qc44I8x3Q0NCWf
ML+WP/ackym1f4aeX1uTguZpUirk4FqeJxAvG687ZmNYLdW6HK6dvTHRsdgPEQ48
CXj4ow7jvA85oR75ii01YX+6AeC2mCg1A4+aYP7VP4JEuEVq4IF2I7JILmRoa999
7vy2FRCyGsymAv/0ka5twY3XHgrusA+fh0NMNjq32kiMQ5XbCNh2rSHJ2WPbkpHt
AL+WoNA5vT0IaXmogcejd4ZilRLlvCPmDjgVLQutlGKdkYc3nxegqsURRiVNrrmm
CVei2BZewcZrEHR1UM5Sk2tmW2Yjzt2FLBK75/NMLxzauP7DLzaAlA9nAMiNpdPI
YiMeClY29V1Ug+nRnYQ6YenKzg93e9dZAcqlXLJT8/V+8hAnoP+mQaMkwXRR3KY4
h1a24fIEq1LaT4P1RKVGMPOngi76qL+w5ApZ7zESScGbSq1ooLjPel3aLVosveLb
rfOiVLS+79wjrqvxtX3/oL4HeDBqW7mxOekbmoA4VIb68StP07bUen8XIt6zxr0A
To1kgHw6aJdb9TB+2ybO5ZCl/5G3+MiUZpvgWBzPUwoF8hExuFvN66soh0xiSHkX
UwZrZhpuy3kDnIOM+AwAhn3elrOtxfz+B4z5bs3cXOW/7GEQGI68JBWhjIBEQI0V
z4znjp0EiQ1TVwzfxJV0+0JR0fkNwqhw/q0nSg4UI/IckMrdMExgcdUTtb04vCaU
7ZKFBGooRb7kgGJTfiOM8iJs7k2jThrs6xU79TyS6iWDj8zM+ZWeWrKba76YkdgM
RLKvMMHK1KHOecJvHIkSdJkU4N2TNa/GvoSxrxYFwV2VDDSh0s+qhxs6PNccWYaQ
uRVslkOmNzl+apzWpZMlStQXxgj6Z9CBdZm29U35X+LdLLb38fMIbvFGGkQf0Hk3
XoDQMFtaZQplJAxdoxsof6vwOWuXrSOyTTjoVXx9gF/ZY0Hic3214Nkd9ySSe5iQ
ASTuf4sL6qXfN+Pvra076zNCDI8rSWsIGW5fpb88NkySDflK334FC5uHYLnndWtY
1Zzk7leuGs3+TwiudCd14Eax0Zb90NUggTRw0k50tBvZI9bbEjMHNbUI/I4mn07c
y1189pVUGWgi3r3Mwg/0aRhH3zfrSXLHkRaZKObPATPejQtIOEZ3Dno2+9hP7UJ/
7rTZSzOLspdxOzYPL75S+uAWm2jW6Jw+y9jT9bqdZGlR9NDfww5q+uthGRTWwUOv
gHpglxLiKg4BpAO9S7DRxrMZTZWNmKeZpKgJaJcIVz4AiTiFJ08DeDOGgjHlIOlP
S2cxJqyZsc/EpsiGbWRwH5HCQUdjAWfg+3uWkNIBxmjmxmjScKy+c5TYXWncocnC
jrrxqRo4iTSXeqIp9XSTgRrN4bcsfiQnvtExADWyIjm7QIguDcmw7qtIhF0VH85n
wTTgsnexPl3PC8VJ2+kOgdEKvACKcAmayyadI99dgQSze4bhpo0Vn/QFQaP8t8O5
F+VpVABxfOwqjKV7u2rF1LrOtiAQngdvnYQN7IQrlRRWCayzf+76EVYKl5ThpMXb
B7FHe6lWYXbwlGgWqK7cUiMiqNH7XQvQeFtmV6YKKonYpXrJ9EwhzpjQRJ0clrez
63Ax3rYSYoL1p4CfUWhv70kSYQGT+4dOz3qhBtKAbFF9JDHaroXYlrKb5+F9s36B
Dr0zrSxaHP4MMYNr88zQLi/ujXf9yyR7h4ocz8bHKZ1I0ohqntgxetwrVSuQwQcd
4GK4PIZvJ+Rh7yiJdU92ODyErOhkiZHQMltth9ZO4OsnL10QkTQRDbAAjTr7ZPiZ
N6rfTOKKujRD2227lBhYusdMuu/OnR9zI0DrjtfQ2vtNG6rX6nxnBjv/Ir+I0Ihl
XFLBViahQA1VZKBhodlAISFWVwcarOw544Pkt1VuAHFnhEgCdEL6z43VS6DPPDpy
+od+87PBADfoWPDQ6YGkPPrHeWfI0wqwIwAvCrPatnU321GdhGxBHRZSLhdXEn7A
k1t+bOv3KV3bDwe/jCNFheTZea5OGSIJy9AxD9jZNDbJjFovZJIrx83rFOHRtx+a
gVxuKcQkqzPxCKDg7qFerQZYRClS0zKyPFopXf1rFwhvD5KG7Io9QqVdeGFQA7Ex
Of8C/BCrYKk+dbO9vO+YMvWOdpHb1GZRxGB8ATjGM9A5s4HQHC7TNZ/UAGEzpIJo
S9bACMTyq8K9iGrGl+qtMbybPuo1RvuyrkK6kiNK004=
`pragma protect end_protected
