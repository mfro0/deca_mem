// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:07 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oMR7wmLiKg2uMm1CZiJNKVxAbiZrSCW3IrFAYkutd4bOuWnvk1Cl/C4PtZmZP9Ma
bEmcBEEPeHiOuTjr5IZxaA/qcie5/ev1VJiYQR6RqNWSGOjnbo9JEjGRZ9svOydG
pfQKRuRyJGfPBDIsqXZV6sni1db5kai8te9SGebgZ78=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5824)
SijV2SuHqS88j+tZI1WZNfT1kdchw61WUbkHSKn7TZC+nGZThmS8dA0fIrRy+USR
7OIpwAiKiRGWrMbDellTaxsaqw6CLX02wIMbNpPTb3Adnbnrykis67lEpFxh4T1+
mF7HkxOJ8D3FWgg99HNd8Ny3N751p2vcfh5vhxEz513BgKBTyAwGiwHPUcu7G68q
tocwZiaF1MBRnJx3OoqxRVUARbLTTHB4ayvAOSDeKp4QRSv4HDxdjIOQOS3+Tl7T
DYiETWTZYq06ipI9jLKQXZizEncBP6ItdxYF+aIrDmiqKIbtPdZEmT+P/wrgY7tI
VC/5DIdAMBTFMD7+BcdBB6I0xMl5HPfgPRJguhcEUvIAjymsp8cgCfhOgdfQ7xrE
PxUWF7U/lczaI3kX1swXakxMkqRrN3mGJ8kuAUpIEEydXI1QvWiTtOE9MdGtuzQ1
JGjp8MWSyY+ssXQIgXGeYDu6pE3+62XZiBK14YQU/MI7GuQ2iS11Bj1dSWiWVG73
St0bC7UR3/ogZYyHKtGrpPfwzi0GTNF7Ok6aY7kHDlvcWOEQcjz4HK8cT2cCwrWl
LsTbmjF0CUOm33D1DswPZ+9YjLHMx/PKqqkgEs9A+nYXUK7ixHdIgP1oGUxM6Mzq
LByqC605KovbFn5ccEEXoFhllqsPoLl4A8B6Vc0OMxgfU/+HxHtT2R2VddD5/Po8
oZsGw3pOxSi67ug+B2qLm8rl2vniCNFMKQcXoFDtGsFEck+P2dGtA44WUCyWlfou
6YKv+eH6mLFo7XK/jfcHBFnWh31CRI9nwI7ilkZbHelyZ/Pk37sLMWAHudQrEBM+
2TytG/FmttlcXGvyL3BbuHsUDdPdj4Or4zIMdVo17uFwI4pcKwckDgtSUYCEJFjv
WOx3cqlErD7qdDSo5rTwp3r7AZxwCUm+cWzNA/3kSn6RwtInlqay6ZkOnhiBes5A
YXw6CVywsGoxfTu+nmVAXkTqIzxGOqa1tyZq9pOziWSUcHMAuxt3V2lzQF+M0EW2
vTuu+7lACQq1DabZtewt4KQeImKHTYs8P//GDYotl78BK0qp47CD639jxB2ZjPii
e3ZzInE3F9g4UnfkaZSmLdg/C8QPmIHhk6sazygH/Jf6OUc89xcseUH9zFMP8hDY
z56I3FclO/w1wcrogpg6EIABlt/nAT0RsVG1dj0+GKnFEdVCorb4vMz1MDRmNCd/
67wU5W6dgvUQasWuihiS2ktR68k4YOt+m7pm5uGh+AgYKv6Ve3ijLLWiAjVuMhi7
o8YAFNU8P7z+LVXmy3bs+bMQT2wDK/KlCic4VHVMzjYXQnJWJ2VCTnfXmbtkJTqQ
bZNvQpvawJTOj9GrxvvaNe3+z9zFCtVFna6Mp2T2ij4BZgexn8tbUTPweWB2qfB5
xWFZ6TNJiigLPYvBRT9RoBluJ+uHBlFJwwCDRKiGIVZxx0NdakmBhUe9Dm3AKdKE
zdYX/KNOsTytJY3zAsBnwz5FDjpTodj9neATNFXoOUFr2I3jrWojI2qaqds9LRsK
J9df1b3B8p/P3+Jcg1QVx950SpbUBzCEyStWX7YD3s8k7dIH0QDSXwRhiuB/HxKG
a7QWKBPZvrmI1VFhzasTI8Y/gqmH4SkEQSbwPHutV4kuSRMGfEQ2hXGbErXjuFLk
evRJsebXHPq3Elg+NQ0fCNhxwJaj198bREncMUs15azp1vaR1H2oqoVcNGoyQ8sY
lOzR9TmApVnANkRMOtsud2bK5zTbOmupGpNR6Sa9NJMiq14TEA7tbX9k4RrbFglC
c7xSiOWECCzM5hhbr5IdmZP88I1nYsRzhaWpM6uNeJbDJ3bswuwhgjb143g+SwR/
sdCakrGldlqhfFpfVur8z9JGkvxY8erF5MZNU4NX9E+iA0C6A2KKj+k1Rserghx+
gIzMwht7UuXNzq4M05YbbLt3ahDpzLwrmsRBWJnHbDDc5Ve1x4mPJ9NsD4+sQ/zs
FtB19wATmlF3ZsD8I/e4wbcb+SJtLhFcDdSpWy+ahJtIE4BYuzV5xl8xXaUE3LMp
RdsPP2qqKWDJNwRx/U88VLbxCoIrG82c2UVzbM/ljsp2iraKhPWSoy/Xr4xADP17
es0ttKUGk/gZ0CqZ2WZQhBPtubjpDny5OFmWrbXkHCjHQgYJ684TYvI6lAKJmIfO
p/QzWa+Fa9KYDJHboTJU70eFdou4WnYCJ9LD0WiSErP50KmPC8feHD4AjEEHyryF
+Ul1L/ccSg7w/VmljAhSablW5M2URL+uVsE2oPROLIh0nTEnCGgirHr2FX7rQuQO
TbEs7CsH5URCFpW/T9HGpftmqSY+6l9hjEbYwHnvzmYO1sjvzJSuVy1IN0rm6fxM
Y67pXWbeYf1sDuE9Ez1VhKSwrO4mTQ9j/Hw93/Z0VL35kVw8vRhzsY2Fiwwc2uNb
piWLzgKyeqvIPlUp+zTGYdVbAK7InJ7x/qNjmFOpo7BGURjWJRyM91ZZWIezrYhz
auQet0Gp6rZBl0SnoFA807jFiYgKpS5cZAmSZhnjFiGjq3nEkPSbrPIJLopRWbAh
9iawLqMpNxtRw+Hbzyoq9nUGO4uR6Xy/s89T6QJyi6d93ErI+ltPz84+qfNEsH+K
NWTWOb2vT/BWSvQkSlpMo54Md03v/cF7EYBzum8fH3Qb9wGYhOINjAZK/hPY5JtC
nU/pPq3G4UDuRTZ8ME3FktzCL7JJ3qR6H9amsDbPDo/MfsKCe4rC2robIEtayt31
pDYb6wvPt/K4mIvZmBJguTCWlR7mJvRfhLdUkv1jbbfommA+JMoR6pTdcVBcBNcS
nAVaHiXobBe2Vx4I3eKYajrL0rr8bc4voJwgBRBtJn47EXKar0ZfRkPzmFJa/sni
+9EhUTa1s5wAZprAecfeVAudg7YnDVRsL/rdvVVEgWm81GcFeNG2LSL9OoffNCjP
h+2cCQqGJ99wd7jGhDIsaXsup4zUCRXe076xvn6ZrcLwk/BwMmmrLWsp0IOF7d3N
5JTa7pjUc3QictnMUBHVL3tLtm97HaPquEsW1pKtIs+cqpOb1tm/UdxH6wEqbBUN
176tIYYY6GfysPUN+8BetCuKLO+HwnUTv6EWisLiufweORF67J1Jp48WSjf0+kr/
wbf66AvW50ER/nHFbGs84eIiqNZqvsUYIOmoSkwj6iIXlX2YzxN8x8cmCE65wFEd
NhxoEW+/7WzTBC+WYywlEBSonE2Bx/9W8lgKI7DZFBlRZvJ2NXaDgyTUma36idXK
TkkUCixxJnN98cJcmhKlNYsXPi2AHMqeC5q4Ezbf1NOUOQtRHx8cHPOh9rx4jXys
LDVRZC6/ZatqglhZnqegDKlIcyZGAJ76U7ATG/AnmVH5JhonHK7JEXcRKuKJ5kyN
gr5bHgppPrMdDVb+0ClvNggBTNzlCQEUFqzk9PXyE4ljf08+3T/lHjwKoCqd5dU4
6sR9oBQzlaPbg0I5AoWF7ROMsRCS2aHzzIY2dikn94/Jibme4PfNmz+YqB83HSDj
gVpZDq8xU9K1oBGC+6PpSiTu4JDnyaRmt3Y1iZ1tpYsxNvJgIkgxBQTiy2oF4n/A
W+Yps0F83mq95kSWdzKa70L7II2tq3LNOACVPEOf3CQVv3PIl58TnB8EN8GayNr1
byrFEjn5VEDSHrpMf4pAYS90hYsD9kUJlewqRvO6D2g2Q9T/jjES+BYQpyx/luGZ
40mAtlFO2xNwweKPTi62TrP/eIDhPISFJ34pYj9jsC4Q6aBs8Pdp4ioAj640SvaP
DOCQwKX9JpEZA4ND3TjbU0RCYFc7SddjaWvKfiaY3R0kZjrvxSPaxZJQgdtrW6x+
UweTIkfqASnrJqHFmyzrvmZPjendB664hPhlHQvRt2NfbfWc8A3JKgh6pNP42H7u
Lh41Zh54e47qjBZFQFdEya7p7XU/vce+X4GwCPkibBnkRZXE+Q/ROyiTCaF7px0Z
4mrdzx33I/u5cGgLZmo03+wrP6eBleDkSBxV4p2JlDpjNOViDtRPdlc0UHExcyiK
tSMgJauuqfTXCfTiTsqvyIFGWxAF1tS9FleITSfO94E3AQwGmYsQ2oClCRs8UkeT
4WUzShN4pDb7DMcWv8G6BvQiMP0Iwyv5RmUbRk1Q+bO4pNWJN/+I63CGxaB8hWLf
WePmZm0XuGAzE1Uka1W0Gfm2lGdxfVIHNGoe7bu8Z+233TLZEh8GY0JjVz6LWVyt
m/j8f1AhSBpOwPlsAmI6EznL6UOKeSbq2WBY0Ob3u7pYH/P9KqPwxic/DoiwwumN
armEJUHp0xkM/j0Z1gzQpxHGmMgXCwGWd7/+DqTo0rKWf6rI8dzjE6uwMR56bu22
lEM5gu1buhhfJHDt5zqZXfLJhs8WCy1RobWL3OBwXqQ/sPFk9gHFXml2d0S5AW+o
9vlIQjY2QY/nR8RcAJTkL7w7S64mIAlip6l1LFaH8dJJQ3ZnUDZ3UgXeNCNd4Lb0
WD9kDK4wzu3YISmTSf2pSFjco+5ccSchPAMWPr6GmUGoz4fsDmGZY3hNhfyq4IXe
zZMSFN+7tNhD5zPXrxpvTS4pWzWaHSglF6wyVbC5yadzTeYel8KwkD1N8viJpEVi
5DqllAc32s+F32psWYA4s7vqfns+BH/ASteBbePNXjbfbdy0YDYeRQNOzb4OL0js
O4oJ+B2Lttbu8YnFCG12FsNTe+MobjY+SNvsuIJoNaqpGnV0qP5whoule3g/l6Fg
VEl41ewDJuJMvRqeD+TZIGCkD7S9B6xeBThKnr/B/CE25UnKZISzSyYxJmLAjF3I
Gcnn1tV8Nr0jShyTWGeU87q16lrpbFDVfnl2tjwuro+hh/woR/M2htdGxOVpN1/S
SxTXfUCt6YJbm6ArtB8K7aJc7lhF73CCzXFmL8h08hoJguURpn1pIKR+amrqqVet
JQjakKfQ3//ZviBEBzZVEvkQuB/rlBWJxw720Lrk2wp4QAFgQttOwE1FwDdsdcW7
9sbJEUsqpflV4Cp+5rAjw53/JMNBfylE+tx0QgPWVJsn+lgCaDkcQsBoAx6BEMbl
csynCrhUflRh08CDqhbKhwppkGUPV0Z19Kjvhe+Ejb2zTyvD+xC2eT56MXHponp7
kL2pYTsDebShSgo+sDRAiA6RryPF9ydf+GDbd7CC/my8wFdZSnUq5rM+pfbArX16
rBTWuRCoNq7jkQsm9F4DTeRCxJkNYvBAzE3k0FNKD70B8tZC4KPk023MZhVKwPkh
8LFE/q1sBKLx/4nM+tf3N4oka1erLMkNrFblT7GcwMM3fN8Dxce6IXc1sXFlOaf9
xgFwMABuxY7IqQL+1AtBSgCqfn2bB6zFhPxWJtpgPaLIS9ODxrg5OYpViMnrhdqB
M1We6/sAlCSjOGXuKuOpAsh3xhYwKXiPF2XgGv2Jr6IasQncjnx1ZtpkC2MJRlKp
tt78KRrhab4U4TSQ+ZZeGINqTg2hCHfN+gp4dIee29H13ey6iBE1WqvTlSv3ofQU
2uemSZ32mBc6t3YNSXz84Afqbh27CWkpb0Lwe7rw3Hzjx6SrTRgwUZUO6O6GvV+c
avx5AeHldnNzdxx6GViEBqIVwofkaSW+0TU/s0n8pdlLr6uB2/mWwJ9xDrKXujgg
Q9lQbMI1NH+vmtQn2Ne0DGlDV2Jk+KpaQtf3HD/iq+h1tme9jR0RYjSE7AqaeNuf
9Fc8g53bHKWexMt0Ih7djW/4SqPW88skbvptsYrn5W4WaCfzbm+HDF8SRwaifFaJ
8q1EzRZfdRzVo49O/BdjD3lRzCpCW/5ExBB+oywqrbY54IK4zgkK9lCj2dCljX6Q
ggY5BJIuIWNNW0TQhTYHwwjOurjWir/yt9pW2WAVk9GlHPtl/RZGPOOeAQG4x00n
rrorpvwdEUXNkJcTveQrHdhAXQtnCiT9pElI9EtRYFV/8udvqfrX0dWMkvdGxyQV
FQAA3Rfb17M9o7N8xst7nz7UgBkXcDOkgbESHXIUF/B7YG4rSy5P4BwjbfREh5pu
l4Z/kQaY3PxFsgwJ2769czXzSfaTaKw6xKkiqfLMbavSrc2wILkTKlkY+ztPcKhi
uElCClPRCZq5K4BtXsowb7Ms9O59SaEPMjuriA1QTGEvPTkF2BxYzbUq2U7PdbQp
Lp+GoGGk3e5xOqicmsA+KlLmo3+5hA+4I3ynlnO6ThaSzEQlm99dsklmQGbyzKS0
VFgmqO0OuC4ND2AGncDq5zk7DnrV4c93aUdObtXd9ZZoJNmLPoFHoK7IUmPs+ro7
g1tzEvDAlskDKBDZHoUczcG4Ixq5lnEhHRRRLIYct/o/RACrSgWfks9bSd6tsPVL
v5ZRQVXXXgj7IxUvY1zrcb148Pnqj9ndU/7PTdM0HpiZnmaKaGPOim3nRuyrDCP7
VF7YskV5496bSFvfqPemYtJIeuuP43pJ6MucR43cNtq3Z2QTUgo3/uKfCs34Oyi0
IH+F2gzbuD+3qlPnm2MxKagImwZph1TrUE+ACZK7bJC8aEFb5gfxGlVGlMfRwQWO
dIpvB//og8PV0EL1rdELIvcRVN16byZ4xNebO3etmVcoq3heguNcEB+RQiSR7Ksf
YPBHaYNdciPW7ocuJRabE7rWn2Eg9UgLHeOy38hsjKRGxV4euviAatGspMCDcR9R
9vG0CyrirDqShDe4V+N78FV3k63s8UT107F8RFS0DqyuRZgcmsiIuCUw3bPhfqbY
67hTw8/AJkwgAsgQ9zXk8tLvdC7KDMNU9AToWYbpoxGOMQsi/pHKcCMkG2KIQdHo
DRlHPFS2VpSq7yCHeh1JUIYucJ79TrJL6uWzPEpMHnNQPUqKXBJIN5gG1JoZJsFE
Y1Cfu5pPqM1/Pge09UzcfpqSicVaazik4EQ8r7N2moRCvarV4OMCBq56TYfcYq+g
V/eDynIJ/xl3O33+5ZEREnKCaQxoPqaglSwLtnzch266gUVBtFYbR8OgPuv0Ce0P
53Qq9lxvHy8xIWB4+aWnTEOHf9WR4oW3pd+dn2lfDYevVMImPlTvQXq7Cav1gBFT
yDrWCdFzHiyxYdSSg3eWfez4l2P91M++RRWYM1uhT7wyOh+yS0jr6gy7h/TYSuf4
USLAfkBUq3r0BJhGSJZph+eF465KjqoogKfSbmRGJzkzkJtWR9eiC+lIt8h7bCrc
wZUUv3rAGEwqvYU1qIIGCbYCtr/zbakQOV+UWqHmQzhv6mJX93BCbhRwkier9j34
bV2ge7sBfzFBHmAV1oIbO9dweUDMu1yxHw7EHJJQ4S5/ZuEndqfpE81La+ehvAgu
BzSvAc2LhdpR6QgO0ubPuDeaYVc/wyshii8KNPj8uJQ3fgs7UOocwNP6RBJ0Fnhz
tQFw24TaCbsB99ADb36B0QdYxE9ddx/0xEEFBVcGc/OeyRsJ6npstzzo5Vv+HSW9
nQEkKHSQybGWkL89RnSXnEtyJd8c78vaNriaEreOxhRkrUlKBpDMMZ52YRP0ewQ1
6r+GmRknUXIsaegWfGUlZdjMM4idc2X6/AMpcMyx6KBVkcGcmmf7Z5gxdcnHqOTY
aY0O93PsUqJkklkGfRDyzN0qfHx+ti5sE+bltyyNY/bL3DUfuzbeq2z6Qipo2fwQ
ZqReDu8GLYnSUkz6Buchi75pj1snYS6gBTvmvTUWBY//dR8+s7R4e/Tw4IWowXkY
ci0vGE1cJ0TW/Lq/jnHc7E2QuxXMuvOVerEXtprMUb+7kxolayHUlEak5BBIYNAt
6mcLLB8Pl+Z+MPzAPUSXCw==
`pragma protect end_protected
