// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H]H-Z:K36QLW$N7VREB=^O+/<N/.%ZWNF<G,",HF-AM8?HN5H^2)A^@  
HE2 O? '@%[+F@!2>I967[D\J87[4<UZXL6/KB',OM/E# <*7\FD]*   
HBF@KEX!5I>/DOX'XRK@2H?TV+DT,8Q:4[^-;W--OUALP%,%@#PE%<P  
H2S%6XCBE2BA:4]X=0]XM$TT;!;Q-;N"">L!+(M WC3R6QX['7L*</0  
H!-V)Y"#,M: V6L6KR+YG^Z&TJX TU1"31MVVDGP+'4;NMZLW_]MWM0  
`pragma protect encoding=(enctype="uuencode",bytes=13744       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@?4FCQP&ZQ(/$GO[)M5O-!5G6:,CGXW7Q$=/Y(YL?<)0 
@<<)I3DP]UP@9%7WK-5)1"@B42+*)Z%W2CUWR0Z\Q\Z  
@>TC\#6[VX[R2(W'F.U*8_1Z>!2.,%'3^9Y3;' >#LD@ 
@'2[43A!#'?,<Q\A&YJ.6*9>QR-_8!Q83FR5V1_H#=\X 
@9X#9LD;<Y.&9 ,O=Z^'@1,AGDU-="* D@QLA4CS2N^4 
@KS<#<3\?.O:*?5KKI(?JZJ+<*LT20L10+5@JO\IBRE4 
@/XQB6X?Y%.H%F/)[4I""- [X1C_9.H0[&MU4AV:R8T@ 
@FGZ'B+3,"LG#^H0TTFRO!D\$PEDMB=+8I-/Q4C6X)S  
@Y813#Q(VE"#''N.0_G8 YUJCQ2J,7D\ (?63Q\N&9"8 
@/TAXIO" QY2@HG5)*RQ>$"3,<!P-AY'L\37$/R+L@O4 
@6[33'G,KMU"2JW:5GHMV@L8X)\R!#S,J^GU.O\3E6AP 
@NT.08BO0Y>E.0)+?P ;!B1P27+V2H0+']7RZ=R8S%?, 
@*2FN(--W"H1F;.0 N0$TX?W3PL7::[4#I!O#C35%.HL 
@,E%L7Q#3>ED1R:VFP)6G5]9$$@;=#?X/4ZC-Z+RD#%H 
@)LRT!I$/Y/#T&EJK:QTDD^""(U+)3V=N#[T1[:C\$4, 
@E]<-;]/7J&X)N*18M7K?$^V77) >>O0[%+E9=L^4M0, 
@AWMR9R'ZNS\(EZ$BF"#IX>Q2=R=7DV6/]/4P&'/DM9D 
@NQZS\Y[/$>?4C.+&Q3%WYTS/ROD+TZVRE6/.[F/%D_< 
@7. Y578R;SZ0$IBOD$%$\B$<K7G!Z>$L(U9#91XH0LH 
@,J&=6>NP)B@JNJ;3%@'I:.O]#G+\:!U,1'GDO<E'DH4 
@8VSNWRZUSI?O2^=WNEG+=-H]3Y5P'NB.ENL=R&FGS$( 
@?$QBGA8]LJU\1&U1MLPNL$UG*=D$9>G;:G!/B8R7_B8 
@!CI+/FMLV7N^F&/US@%93NJQ#I:GL@UH5\]83>1SLE8 
@*PV-/2: GJ/E+-<R.]@&@)W-N )XE/DU_+88*FU(CPT 
@U(?SUT]W>V_7P)[W- K-M\@\P:74I(YE8AKY[+.U%_$ 
@Z/>@17NS=?XQW($4\/M;<GY<A/=]E JQ'S>@6W4?G;0 
@;<QGEAX1]B#4O&:M=+]XP5<6S8O<6;&YTY5\,\WEM,8 
@,^]!HKX"GH9.%KG<O-NBU<H$H_L/0-'@"^[Z.P9@$+8 
@'#WYTUH+-EVZBM_R3#P614.A;M(TH=NMGG>K:,_/R2P 
@H=9AXV?P"LI7(;>CF^HXO$EH:T]HSU3P\RPL_:[/^@H 
@ 4.K0W 9*'-8QJ2P1B#9NSCDYIIQWI@G*W49).=Q(>L 
@S@A=EOJ]#XN<]9K\6XWR0 :)X+C7(ZV%QT&>J0MKGET 
@Q[OYL)LH\?[TFL^*T UU,0OR=E!Z24R[0)_6+U[_T#8 
@KAF5D5V"0?[LB$?R#;S_'17.8\K]7^7HN?KW"SC*=H  
@I,J6[TQFB$ _YJB;2GD"ONE[Z2'&5K&0R<4?Y5E"9WD 
@J58_6.*@;$G<A;"L%20.#RJ_YZN"M"MFVQ32D#3K=I@ 
@>Z/G.1!@<&W2>4/.J6@<&P_ 9Q?RG,J^:;NE4,KQ#^( 
@:L=,T+WC%2FS'J=LD'(DU[*Z&3;?X<JY@K)*EJ<7TGT 
@,F]O/J L-0*$QLV[4I!\,=-,W;SDKQ0<Q*8U0H=ZU[H 
@W4N"DO"8WSU[(!!_CG')X#GE&RQC,(9]I+Y$YFE=+]\ 
@A@!$%G'%03>3?O!WHKJ1HQ%\4?41T3ZRH)R3H/<KP7( 
@5!<=FTB6R<R@B0=F =^HMWXB7E]#AZ/"5FC*,GP=6", 
@H'@?!FH22;D"\J_L';KK">PY@MV60!6K*A :!NP=3$8 
@&#,.O)D)Q?*WQGO%AQO?*RU/O\%]0 $*:D/*>(Y":/4 
@]WTD"CKQ+==5.BUK/(==8##GWXUI,/'-5QH+.HO&JW8 
@%2HYXQ_UU/&Y.2)4'2;FL*2IBA(JJTTO!2#+RGR0L1P 
@J'K!5V>8VV^NK^)%N7IDK[S/37FW.>O+UJA@2 .&_Q0 
@L^5[%\F;84R])JH.4)R&+=J#<+"XZ#P<((KZ]55!X9\ 
@P9S_L]R_10RMMK^E#_(_]A3BK$6@[M"%);K(=VO'ZSX 
@BN#D(^("CO\$6?_H0*QHN&<MN8&6*(T[X0MEHO*O8U8 
@%#\SO%9 X%DG9-KH/3"/7W,[DMQ9R?_-LXS5T$#-:KD 
@I1_$=@$Z/8.>BY <]-B9VJ89-6)AF<QHDYX+07*51!( 
@>W&B6#/)]*YS\'C^&CCGUBE";.)'9[QC@YJBEK*4V(\ 
@X=E&YFF=+X0V'2Z-F<-K%"][R(EVOF\M-W/4KMS;0;, 
@0 @VS3)]. S#C6,,P$9I!2-WD1=XGUJ-;T.9!,N=)D< 
@C1UVSPK7: V<+@4#%AOQ&9,DOHRCWB?!P>MO#;?3;YH 
@2"_#</R]NIB+R$>#B@7F:;"H*8<DVRTB..._+AAA/C8 
@DZ!.PQS2K+]8A") F\8OP+)JN/W>1JNV8$J$R.:S"'0 
@D5TKQG7 I.$860\"NT<C]&>2WR%-_ND5]3">,TI0%M4 
@:(Q(:4'4,%>PH&P;?,0TAI$_7[,$ M?=Y5Y3QYU&&<$ 
@I6!=X@" L:<=![F;!'8?8S'#T50---EA*#B%=EL\R0( 
@HW]^]+8%@QHJZN0U 'MQ]KKIL(N"G:N.JOGQ=A2(6NX 
@:;5X>&$-?"K&TTA[GMQ("HN(XK]L)0V1A[K++_/DVQT 
@XP8O\C /"MQ"^L<4D_E8N11H^0CY7#57V"/9$C+1GI\ 
@8ZC2+\R@N&[G3% [K?=SJ6GJ[ONT/[$S&A#>JB'KF]( 
@7R1WL)K\5D)XY376RR:17$^?=BC3Z+<FQ/04&;Q*DTT 
@,@4N"P!HF",2G-BS$78*C]0&P-ZV0=:RW%*A:<GOT/$ 
@,$B=@8(44Y?VE/MNYRK9B.FL9]:THR)=U <LAEEXW=4 
@7-\JMF5GDSBSBB:+?L$T>E%T^K8U7[U48M\]T+8AV?0 
@Y-]0+^ZSKNWQP8H?1+__!>-#)M!#_=4PQH<, U 5<+@ 
@JG<O7W%;:41_OB&I)8,KA[KZ)6QOY,GGIVJWR2N;+"P 
@8+>KMR1+#N)PX4_X#[.N^"9$T5YA"%W5!OT5-*;Y=L$ 
@K4R5/!JM[B#$TL@-(,<GBQFKQ^S_B0Z(%F_*0O&=*H0 
@Y+@%S;")D7WJ?U>SDIIAPS\_2TBYB8'/3E*:NFU9?_4 
@9QC[CO:%B4XX<4/47P_,:5+:]0/O+?LZS@:F?!ZZ[4@ 
@[U5(OB\"ZQ.C'KQA[5TJOKW_,,GE ")I;EDG@<M17X\ 
@M%#)R= *$P?Q=8<$RMV&D6?D0+ &EKL-&$\WW!_^SS8 
@V1 T,N[6+>D=#K7Z&FUQ)C[W-L:K">ELX][[]TC&E;P 
@Q-ZVZB0 V)GWI/H"AP'?)I:HM6E,XZ+NT:%^%KX:?*D 
@SL@D8",],IAU*5.C2)HY])'*":-S&*2&2#!#;-8GVK( 
@:^/2:O>AZ#VA-'5NQY1\.RW4<8,EQ3/0<^7 I!2WW+8 
@N&C.'+,X0=U:E-__[P8:^VI)J>5%(7BS7T,-M3IHS/T 
@NV5Y9TMX\0.%U$6%\ >S)YH0/V>QWZQOLXT$-UGP!J0 
@R.FP0/6A#(CO00$/?Q$4F[")^HBU,CC&[H]*OV)G.J< 
@6!OG]:5%*0\1_P-O4IABDT(*6SJ273"V[N !.87\XC( 
@[\"X/6*"/R91R\?&-G Q82<V'<6C2]2]Z-61;=A!NH  
@+?W5G@T>!->UFRJI?'^!#\?V0K9W)M>W:!6S4]PR "8 
@^*60!5_IM>FS"WE3LNI)HRS.-CC[>8_+A:XFFNP R%< 
@@=Q;!&;* #OYRYID636Q6MRKR*--<H!>U[AS+@G'AF8 
@.O&Y$JGK<<07B]>#5$%"<4H!9\+M[OF/V2$C.B0;>AL 
@33?^/0U^WUK(":!H)EKKM7PIM<W:9'7G4\\!>T1-]SH 
@'"<68N69G9@U^QG.-++]9\\Q:>[1NYWX=Y1#[5=+!G( 
@BALC@O<DT@'M8.=S>.]W!=_$P_^>25/=49Y5T];07=, 
@?XP?F90F(;&K*AAA!2&_:@7"LI],M$,]'J)'3?$V3^< 
@G(T/@S$9+CKH+\H*!?YB2")<D!7"&NYU][X6:[52I P 
@+-#U\@326UCA55FEET7()VI8K#HVRZSN@TII@%@D 2D 
@+C\=WT^M7+(*O;6;%=K9OA>$%$[IMMA ^NXD ZOC:<X 
@A363J-?@&2OE.E_(3";X_PJ5R15#%K.!T"'7#,\!=XT 
@T_@-F@&U$0/++805(H7C-"0S0%0JGZ.Q+C#G:,?>D), 
@F ?#Y_>OC>]<&@JD.C@03ZM+7C_P,ROTY,CK^K=8HP$ 
@F&+I*M-"N^;XCLHX?]**,2.1(72H&C4>$P^\QV+:"6P 
@'Z@AB%8Y=<79X%<:_RKURI!Z&0QIC#105YV_;5 G1&\ 
@"D&)77$J<+"<-#[S0)F=6NFK"3C1T?-'W.'J5A(CGNH 
@9HL<SH.84I^"K/23KDQ)DL2GV\DT0"N9[]U>W@KIN1$ 
@8?O2"@/73!5!?R(;@)5\'G8Y3PLZ2<V1[:6^2//)(^4 
@:J_A9=?'\= "S_<Q5+!S1[V%>H/ATU^!)J*] CB*41< 
@C<)^4YTB>T*'*B/J;A6Z<B,MXU2D(8!A6*#7P0D#X/$ 
@D,8W^^(F-;][H<DQ^A8HV&<,J2RO"/_#G,L>SEW_)&P 
@'YFA,)4IF 4$3,@,H<+5<Q2X%]S%+8_O>S_JC4?6UJX 
@8A5ZU6(!%KB&E]C MA7\ M1OB('8_(R@,9#_R[Y<7Q4 
@A_5@2T?T@'N]WJ\(_2XZ#EOTWX6Y7]/^&NA^^<H.EI\ 
@(T]E"DS0D"BYX-N&[G$L[,I0]EJGR\B#)Y>F*Q$9FY0 
@[XPZWNZ_\G@A954,(:ZC:9%FSER_M>)/NVNU@G%[\:X 
@A=BMKT)"^HXF*]$6M@D_)2J,"0QO4(2S[\  HH#O/Z$ 
@ U9\/,6BZ7K5%LG05<R]O%5(!T.@9_0;Q\U&1''H<@X 
@$%)*R;1<<G+=XNWY<$KXRXJ^(Y9EDLXM!G^CZSBH4X0 
@CA(SK0XAP2.'WS74]3KSIUQ &>[%B\8RRQ^Z'G<  KT 
@NP7,G,Z@1\'81#[*VFP^GR\L4_I)E["D0<&^1;F8\'8 
@0?>2+-=$QP3"'"H"_MC;+.J10H<;CUJNJI'CD%.!=^P 
@ \;%)O@%M!.$2=64H5(<.2//V+KG;P)P54D-K7:8F&0 
@'4220PBP![!\&8>XN:JYZ]/FSGJ2TLYR\]Z:NVE?W/< 
@-\M6GY&ED@VT)T1BF2_>G+?6'IAO,9S=Q6T0!04-.UL 
@:)@3Q_]7#.4A+2/;B#Q^?YIJI*IW2*(*_H*<R#P]WGH 
@VN64W?M'RT-MA.H=R"<?;58(J75)SL2;[+ZSJ\!A7:\ 
@F:R9H7Z?-W-0Q6YI$/_FVGCX-U^[>0ZV42!0Q3H8IJ( 
@/J1[?@D9)+.K+*I8C?S(FWU!OM#4H'FFC..'<':3\Z< 
@VNCU=.CW8NM+C@(*HPI\?P)W#JN:8MYFZ>B^9'@)Y]@ 
@21$HD2V=#5+-Q:E#J"LC.R\JH[.#;3JG.Y *.'*'.S0 
@S=[="BK,X5VQ=MM9&Z%'X#)(7_H^>/R@O2DGB<2/<#D 
@7NOMG'RH/7N47Y$ O)S/$Q;9=]7<\A (R.'SPU^J:>4 
@N$J4FZ=T,6"+ZZ,C=7EH8L]*Y;>M/2Y;Q3(_TL=G:^D 
@=BDO 7%.&DBH91ACC^GIW^^E/U+..L;&E*[_1XSKQ[X 
@[D$'J!06'U>1<<;"$GX)@_EWYOTWF+Z#_1L[&1-%]U  
@V&O-0^E5R."Q8F18OF8W3Q EV[-8$?MCZ=.8G@\7GOT 
@?@DRG-O43H(8 AMRQEW=SYWB(58X<,E>[Y,S5^>.@H< 
@0%DT!!G.4V(S,%PZD7U;&_\35*!F\9],TF3SD<!O=FH 
@Y9RF4!OLS2#2:W0#_RRWZ#R8B _;(-+RC2.?K_^4Z]H 
@$*C*/%*S<>.6!PCL6*Q5"@K73',YM?<>HQ*WK*E"]68 
@K<S.P(H/J]_?T"+5.>G8R3B-=HH/(C8($F1NJH>Q8$@ 
@TG)+#M_):ZN$Z1"C3Z#2EDV:%D((A6C)?6#H%FL@P>\ 
@O&S/V5]84BTR5&&,#"U-,S ]<=?[U]V-$(X\$X\J0"< 
@J1?5YTB));HK=5#?KJ:H4#[%](T&&$, 8(5%0D$.:!D 
@D\D<A#U-$]C;E(P:=U9!YEO#D! &S,@:(G.!;02Y3-( 
@*X7$/JG;FK@*)"AZ.W.@@$%5L9&"%,0;Q$9<VBV,YM( 
@K&KW2"PR.2S'5ZN6T>>D0,"DAA[\<UJR%6!CA>-%<Q( 
@-6T8U?Q3.;?F@Z+"2]^VB^TRLPV6E:>> I]#%5>$D^@ 
@:Q"6#@&NA'ZS:!DU![#9=_C36&Y#)6;APA9>YMJPBI4 
@=1V81=;<^3H(G+SP#OX'D&UUSE=2:NA'/'JR$ U#.80 
@[H>,,E<?.6>C$6*2WX\+(5<LZN[^U)1F>&3-0Z!:@[$ 
@KTN;?K3O$SK)Z-E9_+.KWQM=T*)3WWW,93Y51FM,>:8 
@GXH\)2)EC@I"@.8U1S\F4'G/*1!(.^RT?"1RC@":A4P 
@XVB5R![.:&5[XQ<_"/A([Y^S@7_BDK=X&.9!NJ:R_J4 
@-IE.4Y'=JH.*(2BU/AIM\C_DDPBDNEZ[9.F5](FUUML 
@/9_R%?.J;^=2CG1+:#R"XQ?>3,N+GX,%AU27&2H] \0 
@PYC?[1EN&6]P[YNYNYV!G*45T'?_\W;,),\!]7U/J=X 
@DG%R!@MNX!.>?\>./MQ71 Z&F#FVY)^$<!6P ]84YH@ 
@,#PP7C.DE19&0M1 YQ=2X@&(\L ?&C1T?RY>TQ@=E*  
@C87&5>>1A:"/Q::&G$9SS.&<"TQ!HP=YH[ ?ULQW?Y\ 
@N_2[]4AS M8#RZ"RS#BEL3Y^&R<W8![B4<%M<0^\5>0 
@BNM*5^_1FEU$"%F <=6;LD+F8S41GM2Z;:KQ>E9.C!X 
@UXI,-53S(&*8DKGXD/9KY]PU];FB-E]0,!3+/S,@NE  
@"Q+45031);*GQ"+H.%CO"#+H2.0/.*&<-W#E9J_U*&8 
@1\,#E\+Q\ PC!E"MZ@7T38V9Q.01<#.Z2\LWDF_/:C8 
@O33"L-9D,- ?'OCF57W;(&A(*W>@7KS+UVVC=E(CK)4 
@RGLEP1@;3FS7W28J=&MG86AC41U*CVDG+WZ[Z<(9K1P 
@F6_]78T%.TY*8*3">#X;V;90-=D<K'"K<_[(N' ,+ < 
@8W<F>8<8IEN+<1GE/0CS#?%.3)2Z#JBSVIU_OS#I:"\ 
@^C\[*^/<4&_D'(I#]1DZ%'4PC]E/#V?HTB\Y8=5UP>H 
@C;/X@7>V")9_?F#XO%=C+MC[S^21M_LCA4+C6%9/H'@ 
@Q]#EGJ!]V8R- #J>L((A.?E4;HX1^_KA&Z17PFG!.$T 
@4W9CZ%(ZWE4%*HZL@0O^4]"W8)*D"N9?(_QN+E Y*(\ 
@+P5?O+1H#61;UERRI$2WW$=FRKW*3+Q:ZBZM7K+LATP 
@=-E<)KS/M[UT^IK%F\#WP8V26';\U^;IEOHB:5N3TJ( 
@PU;!YA#>*RN-KQ (^ CLIY3(8LTL;&#(@'$XIEP@G8P 
@@%\$Y,H( "A0%@3"6\T<CI>-4T!J&)G>I0J9GO54%Q  
@ E<^U_6,8\?".VLQ\GA@!<X^"2%9/**]K_.1-OGE/N, 
@AN5<ED=;&V7,$##M\06@FXW6UG9D2%(I%Y@\\)9JD<  
@$E@D78RK'JUZ5HF"!"RSJ3D9;ZWG;:DOK+I\1W/AX_T 
@  47#;KQ4>\P432'?GK-*JF'@_,?0CI.>V$KU!))/.< 
@0'Y<R(N6O^6C;Y/G1?@I#757R+T):\6AP(2$U?'L)FT 
@M=6>,.&3@I#DG5HHV=A4ST]8);,@D8]-X?MN&[&VC+8 
@32UH[<6*VT-/PIE<+SGO9(*&N91E5^!G"<2 %E(Z=@P 
@6'7>_W>^+9W0]RHE.<9A@ZP8V8$A,6!0:4Z5\XKW 9X 
@NPRM>I<ISF[IU<_YDOKEK]XL*F&6+9"PV*'=(-W4$K< 
@7M;'5O)1A[6MC5S#T0PVAK]Z?HE3'.MNA1V&#H>$<6, 
@<,-V]/L/7Y+BFHG\9A;-@'3\^$"J&ARS&'JC;/2.(+X 
@PAQ"(-9Q_1P>J$XB\SDZ5)CR97!J[J8 ZB?UV\UP4N, 
@U/6X]-+,/^$*G)&O%12]IKWF?>XC,@9QP@(%&K**(00 
@K2I2UW'>FFY62Q_99DK.0(>L\^-]ES,Y#BW7  @M5^\ 
@:,_KP><1,IWQ7 GL,X+T2#M2->"*P,DA\I \)E+V%_P 
@(VM@84\F+H#D&<2[$)%A)N;H-@3ER[0:N &@;K$< _$ 
@?U8O2U4$-@/HJD.5Q,1(GK5*,TV_LU=K>$V4Q[GQO?D 
@625'U7P43>@IX'@S=_=N=3I8.YL_DIZ<:'MA/$>M]2P 
@8N82L*QU5OC#O[,_SBD%BPY S7.JE[A"*Q20Q-](Z#( 
@O8K%M%$95-#AQ(B2Q@,4%K5K/O*T_  $30#*A1<M$0H 
@L(2!/N6$U/6]M,!Q<#8I^04(S%FK6)D)'3NL:Y,1ELT 
@#AJ-MT^[Y\3(4 #$=:0JQW[.OF(\"MNX4"CVL6=IF+  
@H+SW8TCZCE#^-0H6S48#MDNG!WH0H0<]X\G8:!>QR/X 
@7(U$0OE7BQ :>TQP*S-1-: &H8S*=B78NIA-X-CB]!, 
@[]<8G;=2LI9AT&#-<!R>[] 65(AVY_APSJ6X^?O-U7D 
@KS:!9MC[A<<8[?9[+O\Y!Q=$+R_L:G3WVU$ E=[_ZP  
@)W$CS0LC[+..%-- 4\>BT14[Q?Y\Z+*T!2HNU>[<XJP 
@7O)]X0.0Q:0JBS"H:1*D\B%P'N=BY4L*-=>U\F]O<6D 
@/'9!E0]Y7&&.M+9W[:-P&L\Y[HI-\)4='$PB,9BS;\X 
@,NWH%_6L="V%Z^T+P"INGO]*\EP;GIBQ5T#+:2OLP D 
@,_"A!-_MKO&RL/-UO]/:8YIUO:RGH!V"TCZ8#LNOD?0 
@S\21AELY@#I,J67^6'=%E<8\_HB17.-L6/^<'%![*&@ 
@N@<V88H,$F@V;*,S,(1D-B@]<#]?[+>:"Q,AE9"=E3, 
@ L:(<7W5CGRN+3MX:S]*NP-(R0]KP_Z^M\[:T)^I^?H 
@+GQAK<-?RX0R  ';KGQ9]K8#%KYT;YKCSZA_S^HDM7( 
@[6,R==Y4'CRGD2CP:,E!FU_A0O_'0K1[#T*8F$)Y+NX 
@Q$/K7T<)+O:/V[_#S(S2I<<8UG#N-&)8(L"Y('SCOE$ 
@(M)"&:MA:1^N&,%X,\.H6_Z%9O"@.LN3D6<XF9]'H2H 
@K297B,/&F&9LC6AF-YC!;+(SU>%+$(??2JY]*9!3[-$ 
@S&G=8)!*9GR!@8JM]CGA#SP%*26].S*OJ%4=#OO-#RH 
@"$_+I$+$BB -NU?EMFHM:.#^!MF^Y GP YMJS&[MZ3  
@V[TQ5K"+NDSE3OQF%[%(<#'M,]KB0FV699: $,2GPR, 
@\9JQ^IMUYP+Y>E5BC3(\1(!^DF5Y1H!$ D&MGGYD:MT 
@30XBC<:P+F=4$4--%?Q<Y8B)T#<K'9VF:M:UW+3UT:P 
@&LU25ZSGUSR-Q"9?;RX_K\X3GEC/R57'']G.394J?<L 
@0.:^A5>A@ B&$B;Q5!-ELIT%4SZBJM%-QKB+"/55J^\ 
@9X4L&!CQYS[OF*+>!_J;L".F3L"G0YF*YN2&P3+ 1Y0 
@=7!E<5.D+83<=7M&%O@_;X!_YF:=O18Q,P5T2OL!0A  
@77[T.FC!048_ZO^GDI[>Q5U,9CPN (I:X$2M8)-FX4$ 
@Y<SH9'!A5%1C1_/'H1ARVFN81Q5_6G!J] ^%A"'U=D( 
@)-SY/FF[KFBYRIDU 0"#'1ZLEYY=0(\*J6(C":R[(5< 
@<-WYK@B_"?X-!)"?"A-"[3+YS?]!NC0NA(*>4$DQ:F@ 
@K%=.//A!UY7>!!0HU0AFWHPSL3OO/U]?[^75K8?.=#L 
@@(7%)]CM U(;OD#OL_%&M@NSA:JNF;@H?K5X^.8C!(T 
@\]\HX0S838=Y.)*FR#JSFE!$TT^SJG_EN5E(H;FY;XH 
@_NFNWNSX;-M_6"M1^H-->M\9;C=3+Y+*XK'B5 ;&4(4 
@!+S&?>P0Y,4AM&V\G+W8:MCO 8@I!GWG&X?%LMM>?%\ 
@<4JO;TG5M=HIC*KZM-E_XYV&NW&U:8)T+RS2&;?M!$L 
@))6*0A1/X* YF([RM#!_SY^9%*+*,T)>0H# AS2J(U$ 
@@0S$U@]O*%")0%UY4,OUK/,[D\BU'%=#;V?KB ;3_*T 
@U]V/DTP@X^5>B;N$XZ0X[$5>UO75C(VZ.OPOUOW&<E( 
@O#QVV_U>U3NW:@@K&3<+.N.*:<OY-?.8 )W(Y)3MQD@ 
@1#1D+VT ).,09QX>!T;_0MKW;H)F ZI]W3)_79['P/0 
@2(>$SBZXAB'>"/8:..AG#!&RPD\U)< MVRUY4Q.5@Q< 
@>?<;>Y@^J\+<AD'=2LES_O-"+K/E:N='0[3(G7622^T 
@U:8\4KK(,8:')7^05><+4C/,7M+L2()J_,X3M7Y[ZD@ 
@QQL$=Y!=4!D%Z=#;)(8?90$7)C$FL>QYJ['O$_B>'1T 
@R/?VA,A))/DP:3!U&S4M!-O=AHK8YTLXC6?TV?J1G94 
@.)W-?.4"T>CHML<MH97<1^&(R+GMV)IIZZ\-T)*5@4L 
@UO9"N/](P/XOX 0;EQJ617N79#P+UYA_8!=7;ZM8C=X 
@O9$/NZ?48FT/BZ(-7V0ZI6*NN0LRA/#B\M>K1KM%UE$ 
@N[T@USE=T]^-_M.^?<;N/:E,0)H_"_U>?+.92J^(S7L 
@T&,[J$V ;/FP57T]5$$0"B[Z*4+VA]:_'7U@(!T<T(( 
@F3%EL- :PO:QJ.U45+UIXP'2EWC,W9SM0C6+_ >%+6L 
@'TI/!WAA[?)9=2WF8VX5"8E;J8 :F),^] ; D:Q@JJ( 
@Y0O!]OA3ESCK[S&DL* P+[\/=X6O]8D_Q9Z6G4==D[, 
@E@4.CC6/7!AQI5G@[@$(R?_KZ)%62LWPWFVF+K',O_D 
@SXKNH_\VA&5X,,KXB *=J4)YQ(SG[F8:88%+_\*SK#T 
@\4W$?F@4^9H!EX3 EP=T4[7 WKDZ[DB!C,3U($")O#\ 
@LQ=980QN?E2LVVIW1IH:UX&Z4]4'=?BJ1<\N;A?J1$@ 
@<IF84Z?>+"UWQ*V(Z&/_OKI*K08S(',HL.XP5;Z&P_, 
@!*FAF8LNAHQ,+<P(K'Q_>[&QR1@SD+:DV*!LB.B-6^, 
@#7*_B@UEAPKPRI^ZF6:8X6VY:,'1BQB=0F$BB]_;9SX 
@:O8SL?;K=R][JO? \N?"M,6+X:.ZJ:+;E%<J?,:RMI( 
@QULX8ZBT!+BRVJB5R,L#L10JHK>H3=EYX7*:TG@IE"4 
@][L3<DP$8B$^NSP#'S#<X1%QH5!CE5@P,W_>!79R+T( 
@.8?&[J3/!_^[[F4-&25>20X&*"ZXM(RJ#A]_?_ :#B8 
@2>[4P;S(Y55<DWY0R>MIG06HCX>7XBC.Y9;:PC[4O^  
@R PF.SV\GCY-%>=Q+-8FEC+WOVRZ<.*=**"]X=F&W., 
@VCO ^3O/M04?)VV&@:7^*"_I+#-<>&0@MT5L$7)^1P0 
@L/S430K\=)QV._S)%J)+%0:-_S]OD)GHG=2P91/V]B$ 
@^+'"IH\J0/I<F:>%=V&F9VE4XWNEL+2M"TJ]IEEPRN4 
@^\9+@]UR <=%=+'UQB"K:[PU=P*-6'$;-;!21KYT3T8 
@S$$V<?PXM(^)PE?2[H5P#F?4Z'PX^0P6\.K]*.PT%?D 
@OJ4M6+RR\&_>Q0],:/Y;[T-EP.N>)"V@>JT(UE3 1N4 
@*MP< UELD2,_1]E;H,>I]UV-"XXD"3#A9<X>N$>.FV4 
@_$A1W)E?F=#5LFS$HEGJ_(#/_Z'0/"71<H%#^_3H&9( 
@%!.72,QY0M]ZU8>LKA'"3.'"U3^_E?"Y%7";5AQK3*\ 
@\F0257X-2^3S+1)F-OIT'$0=@/#2CLFP^V*YE"!J^O0 
@3]9&%,4&YX\ ND"/^GJ"7>]M8H%$F,H#/@[[TA*WSH( 
@2"!D 1&=]JZHG4#\=P09.>6B+M,+WW7&W PSP)H47G\ 
@\SY1UQ'H$LNR2L0 NR3!D:Z"D.O\@GXW60.F[N^QEV$ 
@V2?V/3A0 -%]\</(O$8Z.CL%NP0<[]'4B:V<R8#LZ00 
@]?E(B:V,95)2G?1[(CP+70N4Q5_410FF0:PL&*77.@$ 
@*P]2RW"PD^Q+<',8D$)BU36J?SKP$?5_*@YN[F7"_U\ 
@L"R@IV:86M4O+0,GA=(+"$_>T" HV872 02DP3^6?&\ 
@#><2W,UL]TEZ;0B?MEE9>V4Q<Y0X1O*.Y'<5M( $ S0 
@[8>VQM,/DDU=Y\Z49%_R=-[0>5VB13S:T?T1TP/,;S4 
@P0QSI1>[08:RM<9%&60H4:[@05WA!?"4HB62^3WU$C\ 
@%\R],8V%J$S+%D^K$#W!3$-^.=V]Y8?);OT6[NZ#O;L 
@4HL&Z CA/2-__*:4D;YLA. :6BJ9^O@6&@VO 724P<( 
@?_#*9%7' C]5A;(Q'88VQUF5*1&.56>#R*]DU;(:8G8 
@WMMC<('"T[<@IQQI;C]LF!33/$!@\0OL^K!>EJO]EB4 
@/HP\JVCF?9N-"D/BSE')"@>W-RR:3>>)K5YK+0!GO@  
@.7SU*".4+Q/(37BM9*',J"%"T_]7^/&2Z,A$$DI-7B$ 
@0X/\<_? =@Q9 S25NC(],>NQ:XR:\.%GW0GP"V7($ 8 
@UX(= &X9)DR=X!"02087C\?&AUVZ7]0-80 23&B])\( 
@52<^UH?ZR) 4V)&DQ#$M,4=1Z/1PJ^X^=()JT,HHP=( 
@2(H?)M/!VZ)_-P9>SLC&<=P]?&R8W]S(/_@<)GF1[&$ 
@6%R^QXT%O!J![,'QE,7O*J9KVK7(;*'";6@#"QG$U@@ 
@,4[,R[+T[3!,?R\48;.VXI[J@\-+<TKNHE5KS5DL6-T 
@C&1>4\]8-A;CG2[78,59WJFS84^K8[XFA]ME.9PX.MP 
@:L\G//GM?EC*J^A80&7:R"PXI!0M54YRB^2T%G-41H( 
@7-V(T_MU3Z76$YRUJ7\?N1.RQT1D", 9DD28.IU@I<H 
@-7'PRW:+_B"M&U^=SIF&RSCY1&Q+J;WM^;'B!\>2?[\ 
@:7,24U@1.DJE(""TRUECC):A6@ P@BW5RM0M@\":#60 
@Y#($O8W]#T'B74VC+36.CG''S:M#<H/%T-J48K2J4EL 
@%9$@<0-;$X?X>);EMV,C&_D&1"Q,R;^?$(]<-A,8*&0 
@LT$V)'DP1$K'=<*JV;JS+A2'T,5&% ?AD_3:0-=Z"\0 
@]:Y;-G5O:KO'?N,"?I1'"6IHS4>41\P4L.^WFJ^-V/< 
@A38'VD;_P<Y%)98U0R(1$_<(#@^,J5HHP?8=L9;6@Y4 
@Q2T8%<&^OQM*_^B^:M*2S;5&\E $$-@#')^"9(_*VPP 
@5I;?]0>7/;+L3A.A:E";?B;@,\4/_C/8LB+ !&:NQ]( 
@4 #&F:BV[O@@L(7XB)  Q"P2@+X2.3@H[:LT3_&=NFP 
@"%&Z6TL\\B35L+'?$8+7!4$&F4T]I0ZC].D;6C(\RQ< 
@W1CW82 \D&R(._&"VVPZ[I2I>!*QSC]#%OF@#P^?E?0 
@VI3G,OR0#M]1F2/VUC-)],(*F5?*W1"]=G$^G;8A[>@ 
@5J]*2;^E^4Q'&Q33?;A--0A9L4_F/543?IH>>;&G6>, 
@>A,KB23)TX6AI.=KIIR*WRJW_["DP'6L$!G_'V\V*(< 
@<,IUK(Y=4+1%]MX<GX'L:?0V,QHE>L(&[;Y&S(1N\4L 
@\>@%/[MVK#N>'^3_RO*X8S@+6PAM]N>DG]D1*G:$@W( 
@ILZ(@T%@^KQ*[SG^6Y61)A/B_7?H[C!'Z(LF %-5$Q@ 
@&./Z5](B$-!H[^I[=>SRZWE"OE^)9"E"@$-AE0GF9Y  
@(NR<5FS%,%V<T3U JYD)K70#;#:&2Z4^1OZTTU>.TD  
@."SN.ED*J"YK[,HXA-8EG4N"R5'0,ZF5W8MK&,1J#?0 
@5+FRL7".PG-E54,"?(R@K[Z@U5"SXE[\Q^ G!SXAN6( 
@<NY7SB]V<.\E;N%!/)H^6-O"@ZY[BFWK8ETI+49;M<P 
@<63O-%0FH1B'JVI.)$]J&C) ?%0OL,42!9(PYUPD=E\ 
@-:X'HT:Y24&OD431KQ3TJ:G'*]Z"&L%-G()38&NSR(( 
@%VCT?23_>"2B^QKB"2BM-8>A^)7Z7 J!KXV7Z\?+J^@ 
@*<36[>SWSP;\CU*FTG)% _*+X7 W&(%MP#<RO96Q\^$ 
@2L-J4IB4MT<7!?HTP)JJ-R"]YZ#>])\DO]XBK'P_<2X 
@<.*Y+V2Z:&QX!SZ>Y.V1:%!<VL-LZ>R^'0[[\WYNY(X 
@4U@,/WEF*?A*'R$*>.Q%[_T;1_VRRX&>YT-5D:+-RDP 
@%;,*RY8K!3/O!"2PBU9Q:27?:,"%U 7C1^X@JA;ZUP  
@. ^VDE<&9'D"OLD+P<]PQ2+.J[Q7D?\/>3;M5.OZWU$ 
@! 4D5-[8:TH.GOPDPU<T2M!H]%0([!-GM+PJ@IKRY!0 
@KE#]CU.PYKWC&<<43G]+QS5U$19J>#0,WSL*0I D2?0 
@%R@"$Q#\/IEX .#\'"QD-NO<;BS$(Q7.*%;NG^3.^M8 
@&# IJB\G4H)@LQGMN7\-YP[_H9,\BX0$*>(8MWE07<( 
@,K69=KU[^2D85*ZG.^UTQ2A>1 1(F54*NXO 5D=]Z*  
@'!M%@"$X9;M2^7>[V.@0KJ%78."NISODEK+6G$;53$L 
@]#C*UXL:'0LEW=80:+!<-&794T?C,]Y@8#X9@HZLGEL 
@"#GJHTKR_WA@KH(C1]O[W\*4W(S[S%2OY*<.1^\JE;@ 
@/XKQKHDRH"=NUDY 3J[OX!\=ORX^ 1Z"BR;-"N'B\<8 
@&K/<7@-&1S3Q-2#E!@E39KU@?Z$BWH,NEQE.E/LS/)0 
@%5Y&S03<U_'=B+ZJ (!X>0, O9)H0VC67/V<1;P#E_8 
@R'E@]/<;AZ*'WW0!\RM/H4AO)^Y]]PPPHH%(L)Q=*$$ 
@1:3U:UW3*C>5FB@BSJ<KEIN'+\!_>5')RVF 0$,LF(( 
@?3U)9<L\*ZO^@FQE<DO]MC9SA8G"DCI"* YECCH%:UX 
@71'^T\!\F]%]!>+G7*]!2,H/J/94XS6L!M&7Q&ND;HH 
@Q4JU\BO*49"#"?UJ/*LD,=@1Q2(.WG3Q-FZP3J=.YCD 
@N*$)[2#)-<<&?57(E:M42XF/L_\%2@B-3LU"-!!@+_, 
@[Q$4.8B?CGP[9T"T[,T<_12A?KCWQR]N*R_TZ2O9B$D 
@*2@C4:N @RCBQ9[0DK?*(T(3!*)M%&>EJM\>@JMC(/4 
@Y84<S]A'"HE[8S5P1>B"#:C"H+W ^,;F"$GA50!]ZC\ 
@AO!_J9I\:Q5;HP]6-9:6X\0:5P[.*A)IBV!2;]?SD60 
@B1\C?D8S="Z$181+07EL..FP+>M+4!HG6>9PE"';OV4 
@.!TVDT[@7#AI^$]SF%&=J]C1OIYZ'NE=NIZ*B2AD+U@ 
@%&1]O$& L^\%Q\)L)M$^^YH1U-*7"ND/SV,G9Q?)VG4 
@T75[.4(?%8,T44DG^&\ININ@EGHR@#(O#-H#F2VOAPP 
@%_E[@<*Z@CCJF;11-7<_YY0(=:8^Z)GX&?9MAZG;#GD 
@G$B\DP$2:!AZ7RQ7+(G)%AO_2Q/(J($XB3KQX/C\%>\ 
@"] 55-?HPSB,W@SG^,!;-B"SV)\0Q0.8OZJE+-%&SY0 
@0S,:A 28!DRM";@7.OK D9LM.Q<JQX',*"#B;AE\ TT 
@IH\,'MJ?R5!G\$"4Z,K"4",?Y>LFY2+. %Y0^6U7)F$ 
@@!HZ10"2V"PF4?OO/;0P+)VC\:4"@?%R?W/;["8*ID$ 
@?1]*WO&;&W=M\U$CC(N.U*,TH<V@G*(B&-6J]NIL(G( 
@'+87YU0';>["#--@%R/BO.GA[[#KY9?9^[^'<$8V.BL 
@#YP=F:I,2^%0WMF0V)_D7L.WD<U,7RBY$%]\[7K 4BX 
@@PL9=N4?!A@[C23V T&JLDK(*0MX5=94I$"^?_.AF?H 
@?"NK^<JI3Z$8??B)M_K&0YWQ]F-DDFCPM#A^QP'274, 
@,$?I1VQ^(1#_IYQ\35<;X4(J61F:NP90<.+MV%8]WYP 
@8M"'$TIN\O>D[O<F<E(3?-B*29TT!/W P<E*@#0OM=@ 
@S"7,]@N^Z"(D[V=#?P0%MROOD?,!/_^QVA-U@,%GE:, 
@S"6&#H3X;#'(<C/KY=^R7#Z$-20VQMFFZA ^&=7A]], 
@CV_0D+ZS8?.>>A\-KKMLT /X!4?.B08_)C@^$:#4L#H 
@\5W 3E<;YD8I4]40B8Y$:^'!.30</55!W5,? PU'EWD 
@/A5(_?<\D49S4W\7O8NPM3$,F(KPT,<MW=G7,&7&(S$ 
@22G>39BTGF*X%ONTNQ&!N5\DY,1THWL>[>/]_UK46ZX 
@Y1>\E^0R83 [?C_WV"_)HUSZ]X:=8.A-FFUM4_B-$J4 
@FSJ2D57-*_ORV046KIN>;J5ULNWK'::[4I&K">GE37< 
@*+]R)?^"<>&MQ6(MG"DMQ79Y2KDNO[2:PXHO(@6GF)@ 
@27UQ>YD3P#9R1,$06"3!XBL#0/$0?%YV$]XW*(-W#&$ 
@+4[E5:_!W]]]4F@6P_/:%KN"Y\*(Y<'&B6D3MCV3&:( 
@Y:=G<#GG.3L\I"^"H@':73MAI\0U_N;K@="P $6REHX 
@]K7[C,,;/3=]8"X7P(SNG/FE(A<_=S?BXE?,AVSMWNT 
@^V[WC.(7_!4 5]S;T+FTV4ET3LUBC+ 4U-(3CFZ,49L 
@XR6C.5PJ9PN&!64E[/QYB:'V;HU7IZ8]1F#_0.W7UMX 
@<?N!Y<?3>RUR7(O"7P_3$#6HP2>)SQ6?<LX5<\$3/;, 
@%$'4*4)% T_HR["$FRUC:^G"T5ZUNM,0YE<.<Z<P\$X 
@95(][$]I=W0+$&DM_/KAU1DGE<3.34H6P$;/_&1*FB( 
@+MT4NUR>MKPN&Y-3E\36FI90BG@M</?2*(?D<N_=2J0 
@Q=XL@^:?)$R,M22=]*,K(/P(80"FR:*N!(.F-:SN$H@ 
@./) $%9<=4\LM][8^;D,-C(OA EM3W=? "!;..=NAS8 
@[9@!ENS@3D>P\V9UBY)#S]RR35/W4V1\JFP5<<8/TCX 
@%!TUK\'Q<ASA3+#-+3GU/]#VX/T[V@Y?NZ1+HF'0D_L 
@*ANTZ?,>XW,X5&I-+&W.;2^!@/P_C1DO W2VI]@;UV\ 
@Q_ZV@%9PTBNM&NIKNH"XP;8?U$6SGT7*9\/B2W]7S@  
@AZZPINA,C*"C.'(]O!62;1R< TNU+(8)?Y+8&G/]_", 
@ZYS;L&;.A7 HBP59F).1D=CL ]<N^$7TL)F6D5ADQB  
@)N\0N_D&1":0@&VB:^ 8UPR[MHQPJB15V=R4/]NJH.T 
@0X/DE@3G64;A,>O'G5W_:/^?+?W=Y$69C7/.)Q'+8*H 
@5"Z1 "951\L% _-0GW.8-4#['W_>U7E"=7&),E /Z54 
@9(J1[A<W=>\;*PCY#AE*<RL2<D6EWH%FWOU/UA4\WRD 
@-^\H. M0=O3%.'_YXTS"^&RP<[*;@TO4+<M9,BPP$%T 
@%'AHS-4CB3.F?CW#Z#SDN WTM>Q2K'=,60^+\;N=>JX 
@UC_[0[BDK<RLW0[6T/N7B"5L->82-<BV&F+Y=6B^N<H 
@6M8=U&Q"2<K]@G9J[.,GS$WMW\0G0@K\ICZNAHG2QT8 
@W3<BWLX$87.'6C5DF---_F;54W,[QM8GLV.)*V8FB9X 
@$9D5A<S=A:(/]-NB?O/Y[Y'WLHPGJUTC42EH&HUN-Y$ 
@A\./]'<<A5P,PO<&V+FV<3>'Y'3F"G3; T=^MQO6&PH 
@#0_'.OG:1!OP%9,+,;$72BCZ29=P[>BV@>]=TX/)][L 
@%GRWSN<#)'[ILGYSMN.X@/K#+V\#P94:(_$6EBDX<5X 
@CB96X%*(1WNUK!%P\C^V+LQ"Q7?%7>H&?_L%PEZBC%, 
@M'\+8RRT_KT>*M)1H<U'[S31TJ%^)>72JUI=2]<+P^P 
@\LBFQG:40&G?J#B3:<#1R8-I"( =9[H=,4<KO6>:'NH 
@0WVY'WB O"B?3+T$H_*J#^NQZ;\K_W2BQG>((M)ECLD 
@YSK#3Q\9HY9]WHC<YL/:7GKO2F:LUSU41/3)<Z_1-7@ 
@C#-DZN%AU"[[:&S]T<,!YN,X'"?N]MB,Z4'/\=<;U@\ 
@#/ @H->".5"PEOW^&&WF/O.GR@T$['O/#RT BL8Z1[< 
@;I90>05I=OZ5BG*MCU^%NBM^F\2JDN2UUG7M^OCM;T8 
@D3U7 G[%V$=OO,0W21]"MJMWW'CO&S&(-_G(^Y.;9$@ 
@7SYBO%)SM5Y<059/F&'ZG #-=E6+!1VA[7$5<2(RV4L 
@TFQY-7,1V>]K@4>Q!_@^=1QPGC.* !2Q2^=M^,:I5A0 
@WZ1,#-L9RWO=O#@Q ]OA?:!T5'V,+7W?*JA:\^_D;$0 
@,4G(3L.MPO5T;[/?XFLA1DH=6"7+0EDY6^9^GO2+<?P 
@I6&N&]FXK&[:(\MI2.]/\X?7.KVU1\8"2&/QM*'M++, 
@ KQ^K?.",'+ KARYM:\Q@>=3HQ@G/H,B9K^BMK'-2<P 
@K M*YVU2Y_2D-;T=<[4^]$NJ\J51?)+EF>L8 :UG!&8 
@*NM(;GL!>=Y?"R!L=Y5H$[P.8G>5&?4D,Y68=?_5F!8 
@@6*+K;[MHII(%LE\ZQ M*<$=7I[TF(OXJ0+>0.H)/JX 
@BJ$6E-4_73 ;5+>A!@,*I.7;95._#(+I53HUPR2#)", 
@4$;-_-T!>40M4K!JH@KN*ZENE5G4V]E @T#W;MLCM$4 
0/H))NA($UT1?&6%Z*(PH!@  
`pragma protect end_protected
