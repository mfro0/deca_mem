// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LRf48I0gVeOonj5wHDdZsX+KP4/5g3ku/rUODlEY07urDx+JzWe3Pv9/JzwgtVcaAQw063gsjxR4
AEBGRhp472jlh8gTOSE2olD6X8L53Sml1aTHHFYZtk9XAf8yYmsyEwd+6ytyTlCDP9a4arvGUqKF
XMMsaNCuC1L4LODOfa0w36aESbN17LJoZsXl98M0wu45gVPpRAmMvnkc56NslxicezKHtCvEMFt2
6KUU9A8k9snnEL86lC1vY6F8reIz880eDfyNYFpfxnGSzo73E9N4B+nbxX1s7pXYsynY2jbxlgXC
bISnn1kcf2Sk3ZGXTN+LNfseltESqyIl4DXvSw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11088)
3ISJnHpFh4Ii7JBOBFg/x4DpYjsV7CDtRfmsFNYzuWVbb5PTql/u8EjeLiXAgzgTabN7udZVpJ9J
HSgyMUWW0fKUqRlKiiuRlMXj6UhZ5e/AdQS8TnSCOg8NnP7ZYcbtJbpR9M3lTOtGVYOT775hegve
zDPuEJaI1U1QIg0se7aJ0aXJvXDXYhpj701bARbx6MYjHFEpuCW/2i/RNHmAms2uguXSXbUcoQoY
jZXPqBZ1ynE8AKHWbyB+0+CZbJg0RSBoZ8Usb+niOIHvf+Rs124cFFKJ7+lil4YH6TXrNOv7I11J
QhPl6aY6y/NyrxscnqaEpDFTLCY+Glb54YTLgYtDNLcqXjJVsu9LQQja4eK2pAMFTJBYEDZXzF6Z
KP4u9cR3pr3BpMXk+dC1TCQYgR5RKaDE66U2vymBNX66wRdIh3+MWg8fYwhLg2/gVx0AGdudlfBk
QKM3n1EcZMu3lG/ts7/cLUoUsF5hGHlqYeFcPfavSYfNiaQmFKVnlwoH2ty0cN0bv8pJo+GDWwIs
aZggaFdks10qxqVmikw0+36dTasKk4TPd9oO6UEdBYVe+TPPxpDH6X4hYa8zywjw885PO3UdGj+P
IzYcFbo3RyFVQux72fNVYtln698bdDYby0WH0FeDa6gfkeKusHZzPLNpkBXjytXrazf9+x02aoOm
CIxBp8QZTK+j9n6Y7iQI4oNH8drY/YVpfuvf4uE07lIwP5bYOVJt6PcdtP4KGwuaROFqqr5kwzPX
UZiCd85pMbDqQ34qYt8REIC0A3f02EEKEQgBEs7gudUKXjmegXReAnYGRT08zM90uigggOx+txMb
Zd6ApcgYqk3sUNjIuz51YPqbWrQNzYL6fRfWF1rHxyTSyh5q0FKQ+sAVftsCWc/+PTUAqSvLdFJd
Guid8I+yp8UtUyQwQhFbRvrdfbbPt5UboI3kHfk1eBFxF89MLnnNwW3z8Dj3r7brR7ixwATk9kYf
KfSKkaTrSCvSI340dM/5OuUqfEgNI8TDVcsMr+rRCqn7AIDAuzPVvzDF/LRiiHVT/wKv9+vrcfVl
ROvsV1KzAH8rwX+p1M9RjDaxvk9OVZpPE/pJf5hKaCY9yTG00p/Tbm1mDLBUm0qKoqfu8N+Wp+3c
pf3+3zZcBgnb4uRkbvZGzdKNCTFRu1oXwleiaIRs5t4jWwFAwl1OWAdX3mslWC7Kx+N8VFR6Yurd
K+di3+39LejiyVkwC/646s0VGbEFKMjY5tgtGH2lZnKkR05v2XqgaIKqHwESDg0f9s5JA09R1gIT
L736C1t4se49FT2Am9Uj+y+XAPoEvIRtMUpplp7Dpum3wFb51mHL6M8I1wq9Rs3QftCJfORFyndH
hcIiCxhqzPvasTyPhJDW8XDKVNnQVxgqi3H+5C0ayaeVJhfaXTHbuP56PvMUxuwKdwgfImSLmBkr
KIsd5io2BIYbs6L73N3Rkf27TGo94zGxyw7HI07RbyVUP/CUK9N9pHJn620fAvTvP5/lWCJ2Cr3x
h/Yo7jrarFbEJJC/MsrL4k2eBBAiP/cqPu2+8DeZ1qStNpcXg5Pz60IiI0DTKq6i4CI6eCy8YSoa
buSVn37NJPZwY3I6Ossnic9DV9S4MgYlrVFUPp89PqjapuY/SjhMqUn7QvPPCiMvoDMY1NnmxJM4
zZdyKwBpRqKbsParMeJniSgqm0lyNo5kQbeHYVNX3JUxizx/MKRuibe1UfgfXLXgQeMY426RQGRk
yLNALpwhnZpF06PEfbftiPO92pNbGKCp+vQ5bknkwXX2x7keFGeqNUlYgjLdGU9lWb1CyVcv2fVi
3hCQuboeUGMMjZl/01gjSCpb/oRfAlsXkpjteJdJhbT6ILeTaYxElEdwMW8NdCta0wdyV6sjbhI1
eInEZROgO/vyWA8mA3AACM4wjPLybaIAcO9hbN0ANXdQ8gLrFQ02XT1Cw8R55AiZuMwBM7oDFYdb
YBsdKxX0LFBAlHOyvH195wRY04HxUCGfj7ZailUB+7NS0aCtqenoKsvaDhApqMfLlOoJzKrq4EAQ
paE2dL5vj0avUtgx9QTcetkr3HIoSvMH1gCtb1Ek8vXxcndn5/IyOrsFf9LvdlJMDUOATV51YqRX
7Zzr0weCNJ1g02y+6s+LCcRac8UrFv0CoGHn5LVK172iLqYJf6SoBDKm/w8+GxT7E7VbLV9OBSm+
EsiERvzvThI6rBU6zd6ec/iyHV55dMiqI5sQj62a1U5GGB2xmFEoClqd5eSofC7V7qNNFGYa55kb
colx5yxREeIKVsUGkKxBnkijq+p5OmrToYmX7E4PvSOg4pSmVj3eS3W7oOARNu884pBW97zEUty0
3//79VMo58RWz+9zeoT7Y7EN8DlLxYRcixz1uLsXJGNSpXfOHVUXSGzNqE7cPzPZd1v0F+yjmX+A
TF1zniGYigj43khkjrghmNNvNAFpbkuZaO/KubHJrHzvLHwItWyS4tFcNUxLFZQGAZ5HrwF/OrSO
ViI5B/2DbGOju60TdBguUUCzT6WUBBtltOYuyQh+HSzk3x0Sde5JsHmDm7VIISHeyPpgzxsxYz2N
+7yL/vNWcvY6X0ntkCpmEHC6lfUeVQMn23ncHvwwKTsBV7RCCw6T8cg7MuBXQijagecPHVxvcqSc
UZkpdcJ2JAoUSWOl+j8IqtXJNBeXyUoE5rG/+jOE2hTKnDxllt7D6Yc/eYUX65wBYGdlV1iMOgH8
kH+CpprqbyqXBpEOWMUBFb5mY96ILPVo5PefdA5MsQ7CN4JMHLzHyr7GxWUeQiFeygSitNwAhQu1
IxRAU/k59BcR4D4zLtT1tYHrpwwjPkyAc2J++bgCF7hKtypNM405zygNb4KRsrIGHkvy2nekWFny
Oq1S1sLo3bjb5AfAAUykqcR8S2+WrgUakhFVtZMBGUW7Mx36uJXtwcWagmV2SW7mrc7lPaGtiSLc
zUN74BBUiUjU9d5vSAGGZgUJYhW+mzevca8qkf3X3Sj3TushWBtJbXdjN6VCuFzUXCv7p/oZ9m3d
cKp7ohtwpqvmYotFLPQA3PTJnZUZMj25VFnngfNvXcLOIr4K/D8rvAI0q2mYx3usgwClhSb+FKeU
Vll0bjPUBQbcCZ+ziDg9r0ZM+iYuArlfs9z3G6cN68DoGYcg13Xj9ym8kKJE4MHSdzTZIqf4pyss
NIBCM2IamdDD0lp8/z4vXbcpDKTPBAEcsfWgr/Yao4M54UjBlR968hPOqG0YQGhWkfrDQCOJwEsc
VYQZ+139sRjEApzxaOtAKSgtbXW1X/7zFC+S4DMNLWoPLzDTLUGbmhbJXQZqY/s8ORlmPk4XgpYQ
UgkFlJqL4WuKvJOc3JxXAUbd7XCe1CJViXQBpWTsgfLFsgC0z0G3LOQ2K5imz6/VZfNjy3L79eQ1
f41honVlivLR6Upp6CGr/h5RKjhobLqC6gdXdTr9LRSV2oUZSiNkIFftZRvWVqDz5WRrJLEOXFXX
8Wz3w6eDuJ33z9RHk3WJTWs90mMhW72WKx7r+8B+ov3qsm7EtmV/XSBki9XE9wdtaC8JQzk7EQgl
Mozd/8sBDuzfW81HkYCbYvz2Vhs9q7E+jJU5wlu26LziI2qtzVLYnOfXBGoIrbTWy6J7hLpzy3BF
T3CJFYdeKxnMlPQfrWw8ADC2GH9MovdO3ppoaKa+mfshw72G7NoWSe1lcJ0SGNi4fZzXVPeUKp2m
iaDNB04SNsFfFtgWFlk371U5i4VKqndbLx/O73f6Sn5bSDwToTS/pjzHAekQ1nWR8pUEK9RYj5VR
AiLPpFDglN8z/f2OQTZ4GXFEUTId3eTXi5QXB44attZrLBX07tqGWPPDA7p6o8oAFMIuoiHWsrUh
ho8UB60zdCNVx4T7bFGCeZOxlJ+W5GfCBbHPe9upfBfw1m4t4lCy9LKrfnZiALdAyaBXtqVMampW
AD/G5qLUpEcxBTdgHLQC3OlessjsDtaHQfXqT+slmq1lPJ1yTyCZb5Khjy0SHxyczrb6BWZzLJ/7
SW3UN3uENzBVzQv4NoDLl+NuzVccdFOOLLhqM7SLt08ebUZS3FqiNX25jKDAXOrtPulMUeSHNrp4
PRcJIGsqUlh6zjWhtl81LttWmtdzTNN3PA7vut/B+mFmdNkzc4sgGyjmQTjYLynTUNoTnzBlvnSG
gaVQRgQLFD9sMDJLVMSktBopBF/41CL8Xt0DwyapFfp2OhIbJzEy4f1Gc+NP1+LcNENDEkmM79aP
dlES30LBsS24pl8muIUWgDowCN8UoAdWPebEiZdSxfxxSAEQASSubloX3iB+yhmg7nE0Gsww8j/H
9vHctQ1HwhQhoy4DLFo1xLOQhi4i2sTir/Rg88dYPHpLwNH8OHhJ11mFEg1xcO1vXcUGyK1C0Bh3
eyq8vm1TnEAK3eVGB1SAqVId8slUwmboIke9sMYLIJpCKLpNeAmoOWTd3yPlk/VndamsSKKSu4XJ
PuNFGz48yuys4g9IHktCs9Z/w1YpIldSwrZpKsYXEl4oIThEOkU4ga44EBWYtZnQZQTl+C4NkGFQ
lom8oC036zAUJCQeyaChHKQQHPl0gwF8Ptf1wVs4Kv7CQaDo2VcQwVEKtxijUKshb1ycD0LarHYW
dwK5buyn3K1nLrjEiCnttsiTI/Z/dtilxjcQGT5EbAw79v1CxO7ItACxibBziny4UOzjBN0OflFr
+XABzGmALXzfZSiRDk3ZfOkeqSpRNf3mObMM+JqSeB0tnEqAMX+IXWzpSdq3cqHJC5iGX6czxmTe
MMFEpQzXsCtCvkYLArsAodJ8A3FLr6zm9KMCl17fLVDzbuWDNIviQ0z4JlLUNbolTnJHOed6Hs3Z
qMPFGdrU0QmGKSrDpqMxP85Y/bRivApeVtpOCUnSPNhZK/VMx2U1k1Zjh/Ai4Yxus8E0ID64TScJ
4kOCYOsJQ7hBhAXBNU/Mgbg7VbciU7ObpvrCzPZUtCQc5IUMf030vFySJ+8h76WJLtcm/PvhNJCv
zTuJnJJjSzTxmKQRQbC4kF3P4qi3/1jJ2QerTVJFK35J4SKpBwgcJDP20JMOUW4JeES78OQZ6maG
RO47nbHGmUvO5bsbUuidX8fPCt86MMCfpKFlGHrSxRAL26abli/swfjp5mfWSerdsH/Cp4psxOZf
QgUX8WTNKa8RpfqKMwk1Km5Atqur5x+AMnqPp6l4Re04fDCe9Jvu646sjNUILsfD1mh0XxFMquKf
146hHGXdZqVJI2ZQnMK6Jm9+2Z4e21si5P8XSc57l6Tf1F99HlVFmqYZhX1fQBO8Q0AWalujy9pE
8VxL0jklyAheBPX2MtnPR4Rs/d2s2kyDrncxsyr8v4dA26wjpxG/yRScz4KzWbHQv3lmV1X9vcq7
VyN2myJEiaVx7f57AVlh/x0Uzp4yTtA+055Y5Ixx/YG0IztHCjJ8DwIIypM0BpqZuBCFWPicW5BW
sHemvfT++cdzO9J1S1KIpWs7Jb60OeVdV1s0dQiN2TaRqBqGT4OH5A/+eyEKh0ocR6BiFxJBlHVw
2pbw1/x25Eq0wZjIlRwr5b2Kc1097DTldpPMpgBBgwM7Tk8gYKBNya0reC4rVs+3FMbWUYt38Gkx
MzzV6HNyDODiK/yY9YlMuM3TJxVUfFM3cNDCikapPvBqiwvRsUSr+h2WScRvJm229OrwzIYXQRmq
hkfGzZKwV1DsdH4FF1A0IsPflfMmuLKPu+/OUU8i8whA4rBbIqmsQn0JtxXacYTUMhV/r081jL7/
XFM74x1rgwKlLGsA8lXTgkEIPu9XANPbswOFTpryZL7cnbOX5AGxGej05Ast8C5wbeWaqnx14zSM
Vnu9TNinDUwSjbKnPf+4rGGEcfbp7K2N7dxPii9pvkFV5/UN0GCmHH3mgDhqlc+MtUqPLnf6VLpm
yDqgav5MNgXdORCjMEe7wYVCS5ug/YzJs2LvoMHrTZOJ/u8ADRvJQ3JnDcwZm0nS1D6TTeO1XMIq
T6WSkuCzCtBES8Tm0Bp1Hn27UIRw8s5W4SPPaFF32pVPBsm2ckhBRJcUP6Ofse0LUlngFfHYFKNU
6fAaRKSCMQYzTLx8ITfceK7+8TG9NfBO7UzL7OoO0aUUaTzX2G/Pvhh9TD3uo9jS1z3nCJ1lDSbh
Em4XQuEp2QMVIMfi8h/Ah67Sk+5JXf4d4C7aw2KZtFgeV/8p4X8i0HAooSk3iojhdu7bLth7RHxL
eQXLou6ADgOZ/0i3em9AzBGnYzGh+X2Xxf1thr2IYGmzhWU96bCmSL24fK9DLYDqS6Hh8sIRX0nj
wMfopkeNHkbp1maN5gkTsLYe9lhJ5uQt4SL9II6xFiAuEpXz/Djdqw07J4jgnZkWs9CiqSU8wJwo
ule4R5Fgq8UAYP9Xsh5qTE5/4/GwAaNi+aEibm71qLWrafNxbUp7Dkgpg3P8tCc0PusRCpbvFdbD
kjcx+2wp+1tADrcR14Vm80opPfPTc8Lw+XJ0VkhH78ZVqr313BeM+0anWtlfvZQB1pLhx4C9baZz
sySUTOQj7mgKij2IKOrXXJDnsqRqoMo1vhGcfUqOcHAy7tXCvFMcKmlV1GQ6KKDq0XnDsQKjT3i0
UCpAgybL1O9AenoasbR1xkphtL7EwlTDhjiN8JC05V/riaU1HQwx0RTSHZwvh63ByZwNnzWqHMWc
CfU/8wuavYFa48Gp26OLLYuAOl6VMPQAB1p0StWTciz5ACNOShqef3INL9fmVCtmINiBBMxLabfS
sta+5TrUDLzCZFsuptVzvb/d7jj288q5T9Vsx7H9Jin56RQC4DZH9Rr2Eoa1bddhDlvWszmq5v7y
EaZO6jbr2Sk7MH8ypSDcdrK3QF82HOlcgKOOUqfm9IT+6exYzJ7oFxc+5drBhZAVqBocQbzJjLNB
t0Zidw2UoEYqkzEuuGxld3gTrYZzfW19ImwYxBLU4bhQnx7oc+9Qn6aQqZVodGVGKGINDPfiMs2H
pIT2bXIjfPuKrwQLRmOLC9uzMl6Qsmm7YtZ90JDmqXwiMUXNxnhscgTVCPD8TqcopYyLYcx9YXwy
JDbUWmXE9IE89CbgVOA3QuxeWBhiPkPwKIKmrI4VjjRr/EVXV7t/WTVIMw5trycwPxiuklRW27Er
qAEcuUTe7iDYFSkOFh0pUTlhsngggxObQWMsbdjaxz2RgY0fQbRotmIqqyshvWpWRVlntP9cGn1u
bdWEKMpt3V6wfgsXKwC8Bu0ZzaLUV3u6feIG5Kt8NC9Vuv/zSfZwUEjsbg84JAtQSO4AEUdlEG35
QDLzs9k6wASkl9+rJy8dIExV8OLDl9q6xFDFbC1ShR60vDXkrmlQHbTbx195QUjjg48gLvGfRXE6
LPfVCP/0OJxCpjBOv6jnZb6LSdysZ5VieI1UrpTP61e7i0r+vHBNfY/1oq/EroZ0ZZYbszY/Vu8T
o3ZqoC1ph2VB+OJqxFmYnpzMCiqE8IT6b7ZZaPkTJkEC6zgonw3O0D/2oppAGidQWYTVWu1VQ7aE
AkLoA9nCbO/HPSLQalWHjoIw7G5pB2fERfV+TpG3PY1F7Pjbikxd0hCTAySn3XAYmAJTmEhI6KmI
sggZ2d/DYNuQJlj0PA5v3uT1srul87Fx++CN+5K9jVtBVhykwfJhyk/zrFP/9MTZtgpvvG1mbeHq
D5+uDfFLnS9s2RUsIhYMh2UfrH6VQFuRIVzBMmNcXvxiDaRMuGZ2jdjK/y5XHAAqL0zTmiGwK1QL
Cr1TZy9J+Edpdufu5VyOcKndPgWSMw884OXk00PvrxFfcoIPO7UlFYRI/wHBPciVBRpbmiOmr7AL
9RHvyHmg0e/eOO5oylev+EC6l5QLAyTIG0xpNaZ6w44/19fexTwZH2pWgm0GUZc5FDSfX99FDIar
ulaOe+RaQTaWV23MvRec002K6Z64NzI5VW0lbgLb/UxDwSmeHV7Opg6I9hbONdkmYwGzR9jtISWB
5NBmCKLzUP8OM/hwShC6NcbqXJ1tFUoxCk+wj40WvpGpFdmh0dn675PICm8kWA8jN1y5gJxtRugu
1ZqR43tTHcv5LCgaQQCvHe3F/qri18Z8zk3HLwbXYWwtWtbN7V9ezP3/x3jZqFJpn9pPanI5BTeD
881pgmQKe5wkJIyu/C6vuKX05RlYZtahejtMxjQ33spyGGHQI5iLhM3cQPou/+JrGENnjZdMY1bw
KTDnzSgb0KBlUAZzVl7YVucexO+EX4OwBhgjoQRu3R9mBTbcoO0YIuzoeO9zLViyleNoMBjBkftY
yZqOES2Jtl8h228fo1tUYEVHVDo+pKwZwIsBsBo2SnGnOjHtdHWcQCBN6720gngBNBgVGndFEosG
LDuFNCAtN7bhjiVw3FHaqSGeB3dadSXTKuHIT4eB4VMqiLbO22uhq+n4u4diDlXA1VbpyUYBkyLA
ZNsf4cotVPTbTxBlsewG2kNkaqhkUkLUzNvbKn9aj84PCngolGcc3iwR9GcC0Pq6/GjCbRYWIQll
xPo0BQvftKxfPTI4YWU82DSHiHF+3vhV5lFl3mQTDd0Pb5E2FcWlNy77MglvYqi0Cc3KU4wULYZh
XqbqMav0NWbWYqPIHu76JnZmUgVIURBJ6UuVdpeg+foAvvWgP32Sv9PwIMq4Aka2BgeGJmzpv61s
ko1MCAaMwUFkZBPNQxI18z5vLHPbk3ocAyLdQh8Hibcfzk3JUWh+1SGP5RhaC3TYSp1NRdo0dbpk
SAoZNMBHwg2ih0Qjux37f5lLlWY1hUvHyMQSd6RjDtQvkQsfGM6dxylZyCltgEeaPEXcBBT7PZn0
XuTbJ2jrTBUIeOZVVubPSL0NYavF+vZTCulw2BjiIE6Ev6CDNnWcPWd2ZW7k8BcvlblCGnMDv4W0
8yeV5i/5cTwRX9aFHVMiGET41jx7daI7qgwZkUuBAYYOIfpvzPjX1tmquIvZDONOTijR0CS33T6R
2q9f+Yd0rfN6In/fOOQni4wiYaUZDR5Kj+PvreiZ9p+hhMoMvqnfLhixdTErQleIaovRDbGDPyFz
aaHlG11qg8OzU2UV9LwZSaYcRPc6W8P0xy+OYp2fueojLK5opRQFoxR8uydwFOrgksqjJrpAhE5+
Bl10Su72otMV5nXJcoVNQQPUhiZmjWeQTXKwbrTcnTEklIgzZLbvSQ47P6pm/6pNmeMLTs3FcqM2
deBkDVWi0LxLYidAqJxUwmK0E4SQBd299bHIPVCfIWejdpkpt5N6wIBNErl+u9evTbe4QJZhw67I
k21HxpMp0SscmGQ1wgZwgPlmiE2rbpaewFmp6pEZ4zE2A5cd564yfUes+FRE3aGDoI0MFpzBT9wd
6WA2bDnzcgQ0K5wLBEvokWtKY7SW9D2A0Ld9/MMA7kYbTPZzpsCqFr+61uRI4itd/rrr41cedA0J
QIEao2If4NY3w7qN7bcY8XQ+AdUXVNUPy9dooaN1Ypzi6TOJwIgLkHgQbtiakRlH2JzVzbvTQ6ae
OPIEZPXILaxAvoPKMPPWOmrl7f475mCvuciFBqLWqZIZLV7ulFjbBWG6sIQ5GHlW9aS28C9sEO06
mE46VYltvXOQG3Jy0eDUWzQR/3jHJy5dplhSqFXLlYAgBHLymmBC4pscIi2PRIW6gRV8A96K+i8F
gnT6BlYRCnYnN1frQqix8qfIYeovQCqBM3C9Q028iTE452azjPQKdXblMB6eJuByz4wV8DXQCcJ4
DGnRIJHypgO9WWkuxKxN3U44N3i2/Bv3d86Oz0ITZJtwzQkmVLuxNjaBDHSESIVJ3HjYxbcFvAdy
erS3ji6JcJgHmB2Fmu9FY7ahDJ+on8V9dKIk6EZ6RQ87ntTFC/ukCcYNL2GwCm30J//RXT3Ia/Kl
e+5/dpGn0Lfj138YSTklxjuChKrCh1cgCL4Kjg02D2u2cHUcSeVAzwuDeNsX9WRic53Ix5APlkSF
gJG08b0ffTME5N4UFVi4FfVs/ul5m8wvsO+C91OVtALUntcd+TkCHT1TiDjKIhVq70IYoNnBiOGp
z6kl2uphkWnxTvSZWe+G4lE3udbi8s1ssB8Z+njl40p2VFc+jJXYsmKqnpaVr9al3CZ6iKk85Okq
2178wdP/6T16X7IsZBcCzz1CHXdKwMWH+HJZkpJ4BHFpQRUvDo4Uy+aJ8jVb94tjRlumfwtOTxx3
aPLnfX51pRttEr89rQwpR/pR2YEvln0TjiU7PPETfuO4Km6/FZwTC1+VlApmWsycfJorm3lhcVOe
RWvXgVmEi8gcdmR8I+zGu4+Fxavy0BDM+aLq6+ByU4aoNI/lMBXTwBY+QQqgNUvOSccUANM2uP26
oiKSbGoG9KGh/xN8M6F92Lpz4cMgFgRfduts31lifUqQy/zVDx0ohYXEaHspWroT0AyLtOysIwuc
MZ+uXfkdh5L5CPFRR74MBVo1wbJ7TLLzT0+tEweg157jVVSnm1qDkDDMNzZi17lhJ7trSRf7+QM+
mnTY5+DCfKye/EySEmfYQE2zfpeLt/ypucMTyb2nOzZP8D8Ji5LMaSpb80xY2f4J94wcqHOd9x7u
Anazn3LIt3CX9ymkwcRf7CVw7sTHPXtwan2T/xK+QgwASuV/56l7XWocCA0XgW8jsf9MB9K6o+7+
e1IniDAP1umSrHMgiZxFyiDTrGBv5CnA38rDwe8dIvwZznf4yBWlIxuxuiblhN0oOsdcIf5aR0mE
26eJfx5XK73nShm4cNjjof+YGZI3MT7hiJCaNkOFQrr62lnLqcqnQh2hHK2uc0UBK//xitmIYIEH
8WaJ6hMu22g2mkqhhwrWwAflYtPp11lRt/3xpfhMjpDaBPPSCcpRmay6Mav9CLULM9YpPigEZSmP
Ck/j0Vth+yXQEAt9A2roKLU6rRgJFCAZk+BGGhqUwdRHu8+91dOieVcHkDfGkDENSzIRNTmKudEE
KMhgqTgL8Lm4VmkxqnPnWv8YePLWaxIO2zUMNgGCtX2swfc6/dfIdwReO1E5fbrPqth4xqarXA3n
mmnCEyP0k9Na422owK7rMUQsivioaWCm7wu5Y/F9DgKd9TmIIkKACNrg4AC9LhBA3N85KWV2teK0
2pPa5rIQ2AbkBZnFuqsnMWkj0n32+U3wxi2w/G0t8D8ehcwx5XncZ5+e8tO+tqrkQo5zs+bWB66g
vvUdpdHwS0wdlGRuWYYg2Plw1FUk0GOQL/F8NEwnsUEWJlEqcbQ7LsjRHVfWRoLq8eYNdTWPq12D
RIZfrAB01ssk9pn8c4yBh+KL6FbGHCcRb4uU1iHeFXEc7alUkDTdyDYe7eelqPuQZJHOXd+IlvuJ
MVP+EoQDgVhdtGMYMmx2LmLjdBVyC8cROGJ6aFUPaL3r5Rokj2JRs6lW7/DLG5aGTRLDfzaTdYQu
JpC0GPJFRda2O89vSmv4HfjCYMrngV4E6Ydib5yqadDL/4GwRfMAXBUGgy0eHkUIC/9WP7k8+Hjw
Oh4dul89LcasdfEiLykzqswNfEBSP7408HQ1kr5iEKQoDiDJtk0TXlg+V8NifDe10YnPBOPP2iMl
kEB/8pab3J+JMzSfoU1lZVfcXbJy30e8m2UoZLRYxwRnMWnHvDEW9FowbW6BstZeVkNoG3bXhojY
9fMzZ2F1rnXZ2cXK5ePypYZRNuUfThHA9/0pFVCpQe5Jsowwg+IpjZ8Uc9lQP/QnzfixMJn14n5T
WEwApuIfPY3K7NpwWXPfpQMU/ZC5oExP/sl4CoZAWq1u0nFmcbwyFsBR3sIlZtEWlgdBrOno3UXV
MVHC6qHVbzDGYtt9Inn2Yjo5Yea49fQBVHUxobeMuGZw8d8PR+puVNQ5mHY5WaFRNaWdG3o5zI5I
2EE9NhLzTBeGF5ZmsbDjcqxMWzgh3qTM+JIVtQbOnIifT8oBZjLJ0jL1X7W3fUfO5qTVd7TtrjjU
ihgrCIFFTEa7LpOAK6g36Ex2PiFCFZh66ogDdSKlZeowh//DtWnGEkYNkcsY6c1ZFTXapNwn52Cb
s8/hXLnCAV5ukDUm6vOH9yV70V9cCva/0U/n+aeGFi5tsthVRiH8RK5+Ph5IVHL7uw+e6retFvCz
vZ2+GlwhzSrfNdMInLsJxbP2TxjHPiAaGonE7ahal0wtYRwu3Hu+fen9hTUCCzzL+V0Hq5vGwr/l
zQcLYOogUJlA1LoCMFlIX6YF/qFmX/xyocP3IVuUDH+63cTGE1p9dUEUim+KGaFRZ/cLVp46XgHC
tFuHqG/xOgyW6pzRZ+CzfaEcZmPEoHaNsBa+JLxgtgSjQK99GnsoIEpFLFI9UzGh4QhGLdDdR+8b
/6JrFNQEAUDW3Hyj044KwvYJiMhLcDX8BTAR92ak7NpN0fhOEOZHXjaMJdundWc2pTV1D48q2+xN
PvMaRUTKDLuC8hvrTPNf4ZPf6I5aqtgkLvK4T032uTJ7VISsftNEI7XJcgSEvLUPzBySf7lCx4Dk
fgSzlJqfm5Aist1LOxljEecB7iigDckwP7U+8/CXuK3zn8p9A+eIGk9+ETAnxsB+vKcv1hAZSE27
kHJ+Q+C75HwKm25v6KRupkD2IhJK8MUhWx9pVvUgU7/IEM4DP3q/hR2c+pAzEF2+RUwGc2ZL98T0
6Y2YUzDtkIsVqgdFY8+SocYyzm+OglsmAeLiRrSH733vrU3Rtq2MmBxZiugJlYpL4E3AyA5xjLRM
zrIzeDbPRAoS0WeQwVDoL0VCJ1Cob3Vc1RNUqcpshezhDMJTx5N1XGAyGpfUUvAqXBYV+DR0e9f2
sdxVLQdMUB2YceMpGeguyrSQID/Pwpzsw75G/hMBkftRNWtpajnXvXthhhBfNzDWS4bm0Jig3aR1
00YmsfCqTOPNCwMuNrNzedupuw+c1zcdEkjYaAFOJK45FXz73a/2MXYShSwGn2T4rCW0zfxZMfFB
Hs/54aTlio5e7pC1F7P4aOBCLq7b3rd3NQZdSHI4p8ePggckCby5ZvY6E32NHAU4FYRq9uKz6cIM
BF8L7PoglWwfyeyBTp6I9a3gzth3NzJOJkaFsrDknvH+b05Cz0IS819R4ex4cJIVbzxYoY8gyu68
K69NLw7pv9HLa4jwxgIO/6Y9VPcaTwXCZjKswAJ+NeGVus/YO6WUxO434pwbydSTcyNTxIeGNcsO
XLx3udPMxv99DNx0dPT+KDb4HHdn9KOLuLD/R8dSvwB4FB+7mO3dUioO+C2xD7e0MdCKXkZqNN3/
8sKkQZ/rQ/XF3aS/doltlnxFup39klmvMZ8mnyuLx+TveVDM0NXBdY8slD/44Qx6raGPutoJRWr2
lVXwpwX64iDOdZI2KmW1UdyzbzRQ8e/aGXkHfpFozwwL+Q2QFO8U/QhhbKLN9XuVU5g0nf6GEFYP
zwYORfvNVSLKIUh4NtFvJl+QWOWBMMAEW9WzyNco1ae0amZsWCaVf3WN/yTiAbMpjYlXDB56uzOF
HJ1BaYBwYaPaKtlAar+W1I9nFZ0oST8O9+udb+wIP7s3u0d8ydT7DguO60jWPJJE3Eclj5aod4Y/
JMBj/vEEwvooNvi2Aju2mSkeSQghFUskFzqxl4SoGyTUbvHCvjooM/Lce0wEm9WaE3BE9Ym1AUDQ
B3G0LCsMf1g76lC3CldtdIB/p58vGFO+S875tkzV45ZGHcQfaK6fq35g0hvu9OPXUd1aVNRfTIxS
K/XIoUDUXkHCno2bKaHUk0NecbjXojTWwIHcWdg2UBKrFk2+2YzhN9rsRXUhqog0+y0+IL6c+JyY
u3trRhPGp7NVqTTAr0azYKFHRk8Vo6zl5BFNzHRgMroe+YGwTZwl3G1boLu/tqaRLsGXaBPrOpTd
s+F/BgP18mL5cVAfbByNcDNGiXJLGtYC4eta36k+4wRx6DPlQmq0kBXAa7LFOp/DvltIQ2X5tTKu
ZBVLIEaBBgGRt9sZxwn0jLdLybbdZ6AUC9QowX1yurbFIPQzBKX0TQb33a9ekoD9gU37dwWCGgHN
R5KoPovsOhAGAX7fSQ3yTlLl3ZLBJlMsUC92WCys8N8jbhhS/TbIAZ6NiFKBDBRiCfh/19LcrC8g
YbMCPHGz8l6iFeysQ5DAjxMHO0p8znPYJh8ZyEsk6VvD8epvTBQoHBPrvN81Fw38xFK8SXGabR5H
vjvmicmkt6FCorpaQ3XdTwy+ASDQCVf8Xv3hQjVYpX+D994oqfecxcjAOhsTgYnDH2v/mpp+59mZ
TsQSxhsc49MMk7M3HG7xTP2tsM+EG7c82LIU8N2UPKyeUwSj10CdY1e5g+lNNMUmEVAZUBVcpo58
ULZqNE5MkYf0APCpmpXWDJxk9ayiykSqRkS43HLH+JvEmlrwSNj71wV4RgDMWXIAxLPQBiSH70Ak
z/w86Ll/taJDaoSeNppffz4TQ6730+Uc6nfQgyT6UBOwdpqzLWTF+W7y8oUGP5h/JuoQLhuA00tZ
1TqNy4Xz7HYXFgD2V0EHJAnrvjr1+PGOh3uZLP9JnjFyMikSOSqTU/Bp5kxSMmdCATLP3+fFQCxZ
QFh7DxtL7ws+DqJZiGBtfdxlsh7DOSXAT7IDvL3w4Qu/wOOf3Q6P58Sa5Oef5/FTxG2P011KW/AX
nIKyfESNv6lbVlQQf38DNt2NE0isShFZCWngQCmxSp93QFJbnChoA2pSb4mnUrtH/DwPnPKAa+Et
jyak+CqJBXR5cVBjFYy4YJm6VRujJYU7fyr39URRe0+3doq4KPgKDrdDxkzlsZ05l6R77OckbhVm
l+MYM32WxIFTixPDoAxg/ENJIlD8unrcfPuqpYFj
`pragma protect end_protected
