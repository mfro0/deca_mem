// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
13Mj9sIHASmB1Lc98Nx/OksgvnWu6PFu419cL8C2+YoFKPWZdYl/IspMHGIrxtoI7ZHXwECx1ddU
XRdCOJY4LZVwi/Kr9v8AlYmtRTHUCXN0Yr+lWVC/fEanO9C6MYhfn3Y/L3PEY/mRzKM27KpSpVFn
4M4EWpNRwY9RSn+FyKUqmgGWAXY6omjE8l0ad4sktWo/7zEWFN+/FIo4vgSdsvNilWDmMF6W1Xz5
NWq7erT9hJh+wd7hznoZ38tSIHxD5gWZFCgHyqOHY14dx1GfP6W2fd+9tvukj9X7r8fRzjsFCIl1
npKwsGu2Vz73hP9g6WZP5MJ6rlQINbzoHfnceQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11088)
HEXPJAC4uBo6ImjHawpQhgE+LVgBB5luVG6qYE8JajT84eG6Fw6pMfjWvCiRzNFJTXExXGzPCjNH
DmyhQN857nJQ4b1CgSLLyRgnsuRB7nhaASoKhSUXm9esbTrTAMxAEs6vE4IUtJ28JbHAuFzv9kcj
RyRwjYXsdFUBuKgmcHOoKwmg638WCWQoe6K7ahBlqdOdVGz7AawQ3TJvTJgUmL3FI6onILFGfG4b
wMx/HCYqcUoc8IMEkxXF/KuXR/qA3MyhgE50zfhKSd+q3Bu7UzNWNGxl7y/yvQVhoru7lwAeOrip
tR1XGkHcruKYmA5ZZHNHs19+L/ZJFe2lzg5Wzz+K0apn11UO+7QzEwDmYZZef4kL2OKS8Vu0Qpei
JQcT4W50IMPo/XkBery+0rz1ZRRobcpXsjo7uRg2AThHfBW8vKtbyu5xg+g1FQEv3JIKIZFMSShE
9GpCH07zyhJ3tK2te6E3IfSpDjqtyNUK5Eu1LEhn4HeZBbL5Dft9+/xP3n9R5QUgiuClfCmW0YIK
0ux+mHwA6zufuArR1PfTni8wQcA6C2L6ims76c1CTwkuhN83cPPftRL2k+a7uWuroVu+ApTtNcZK
DsqwtN+Pnh/zcqFCwV96fNxErPEBXB52j1SaYri2nWSCVeP47VYPqtO2f2o3/CSqE/+aKudkHRH2
Bkn9O8VWzVs3lCv0o/NuDo5H0WGKYz+ohOHO+LKeKry7/D7AkNCfI5CqgnmKLsHExaGrkkGXZz+n
Y3UleaibxN+VKBlXqxzIGB9tGtk/eaoPDQAUJsV9DYpx5I2ivTiD+8ukkwSzWeF10h2kmRQPSJwT
2Ah1zGnMR6qZC28KkCR6mbcrA2Yy0TRMIqxZ+Ja8Vu4GpNSbP6gWCJf6jKTsXybgRYlhvVYhjQrp
vvsRZfBrVjSK9MI+O+OkA3mDdirgtQkXZQazo0G9yQuh9TfcsXs1XVaFeAbqr3iEXLJpBeFldaVG
6hhXRsPAEdQ7zuhJ9DFSGcuAXZmllMUhHOZsOUI4waJHcr2dTi9iq6e4pXtz675O43IlSs0/Y3vT
bzK6lh+f3Z8EQRscV9TbqwkpmnC/EXunwCpx44B5vZ40H1/PrIT0mmlaSfO0uVcFsz+gGM0Ng8VE
3n1JefheaTra6xh5vk4/0yV+d/4TXFKXj1ACIH3Q3L9NRyESlDF4xAas/a/atRxMZl0YZ4Tn2fvK
vg4Osl6Z+7bQpHLfluVCxY25IxhAxaYwJ75a2junUOQJUfzk0jKlB0LYPk8GDtooczy49HtMUnSS
HliCekQ6/sCbeqkJAXPONCcEK0rPDuzLXjMN6Q4menrYle4zxPOW37RD1xFl1C7a86AgC4UZ+25C
QTcFMAHPJRViUlJw2nCs4IdYDwDp0Abv1gMRfNFYNPu2xZfYw1G51fuynXMRZhsvbt/w4w+ti2Ne
PFZ6JO7ROmg/NfpQAauk/WJyK1d1MiuwM64wsmat//wVDZkixPUFp49+Op9/rDYWWLKGNSf/a6XA
t4QFNtXlg8kYXM9jMgZsXdO6ajmOXBMPJEqgxe7gRx0fuPeGXbhuJfeLDlDxNw2MY4IpCaLks0Kl
TteI0VJMhgQ/eE9BUCGZvTw3xKO4t/CAwB8MObTbM97n/8RTFCPEWkyt5QIuJd7+iKMVrl8MI5Hh
8LEIsibU+H3QYPiAFJmUFpdGi3Gnl40k4JVqLUvJzH0xeTgGhQd749SwvIRgTzY6hDXNdej1/XCt
LToI6tp/ANDkYzLx0XDfznWcP26WuvtTGUkvOGg/d1abHnV1HbWS8PckpddBzbyrEQRHCh2MVnXM
Hizy3SO3KjzcmzjQ8Epb6vY3JZPj6mGbui5a3WbrvYTRbrqhsxCzDoFEzwfNrn/NIRXOGK9Nmuup
6ouT0A8kbU3mD+MvtPzl3VgVdn1vSsZ82fWuuDBmTwnko1xtZcMuRxaE+sBUWWEDIuTBWjMORusO
w6bxonnod6/plOv0iJ9iprkoNrFjvuEauN5RbxtsPxe2XZ9LNxKSkutHWZbWPycG3tCJnZBYF7QX
APxNpuIIFABNTHbmAHRM0VYp2va7LMSteBjB0x0V86p/2hq2ReFOPbkQM5kH7k+A3y2zjfOrlLSr
tniadZhF9H6JRA8V0drjjXOSVkVPrWTo4T9p5PUZnJIUKu187Bgh0ise/aZ1UFpLC5V2Im/H7N9G
8dGT0Sn479MDq0VVFWxpN75mWleFJnOBWi0jb9j7kiQUBKepqA5Cpv17Qp0gNuw8nelntliqCj3S
4RBHTHVzIWYKsIH8jCuw/m5MViipvMVUdZk26SnhQlPpdhUr0nQaXo28qvqh4iOxktFkOkgAQY2h
DpRqUYyRsERmBIYnNh5X7lTfp5ocIdvx73XkSGkxPtn2rK7nhqFxlcPBB6ChMSoBY2Qo73fuQ6sQ
olUkIUrcX0RnmHx00kcEnGspD9dVXsPhUfJro6V39zY4yaFE76pw/8Sp5KXFoWsH+GBIiy4MpWpk
wMaX5YLtr0gAhQ4uPhI0nO9uqkS7/mLl18v3e5K/6jhcbiL9xL2XGWKENvIRfSxw2O+CbQvY6pr0
DKgpnFDwt3efqE3xI7jTO7aPmh1D8Li3PfRCLirGp/SMMU4IvDJOscqqaJaQMwcieuaWLjcJmBD3
5ySr1k14DpiP5zQiGs1kX6hPZ8s+MUur+bZZuTqnVo0yTs709dbeDreq3mrgFszZDNWGKBqsv5xK
vfpFvsUxFbGNf9uVtDmMG8sOQ5nedlqAZ9/4e+X7Y7gI4uN77aKLIMCBrv2nAqp+xxQSUX5toq+k
xyPE4mhk31feTsqCjvkVMF0Fb/1JxIfshvScRCQi67+Qe4lhT7ece9WK1We41mxytftF4XX0sMX/
iLHfkvxni88KUG/dTXqFLpmazN1ZxOgWJBvYjiivuvf+IPydVSFoQlZ9E5ABIp6PwQTS3Han74Lp
wrLNYYvG+kMsxoawibuNyljwlwcRqZoP08mzC5fTazdY5I6dq6a27wX4actPcX958JiGWylcEA5G
JCck7rQqO6jWMMR3v7QwIXVeH/fUGKrwbcogXPPXNFSXLJTwmaTApPbN3eVlqDe/s8akLU98+pKw
To0q3W8BzbAF9IDOlA7AVTcA2NKUDSYV7BegR8Qu4Fh4B3kiVN7HZieUTtDIH1iXwME8V5CnTB3+
nkvSyE/K7rVRe4XulSQiB9+OXTPMqxd2cyuoq8R9DR5G+tF1S2PQTuP6t6QljNaQ1gbcjJa+7jP6
XFw61cDK/JXAgyup+tP5FBMxcX2kcF5GEu2iWNLIT3DqmOVEoJajlKnyAE1sxGdfUqv6rHSXGbnN
rHxSjU/cnzGBNGJ4JVXgNYk7Mfnxc8UfzPC2c0YqGcvdkEei6sscKXN4UEUKGbtP5/7V5bUvLaWf
ekcamhPI7of9KjN5N6qHdrdATHQ6i2HRBSPk5SJmX9f99ybOlCA1Ezi++P+4FIbNk0VmcNT8xYFs
3BgmEJRlbXf0BwpmuoASnsWrXAxuM4E/R9rbOos/9wgGv+ZJXSXE9/ywQ8bLcmN/GDwM+4kc6DZp
XYW5gP+gG9lCJlh9kBe0i3+d1b4sNWQXggf6hMuAEU2sBajPwh93WyN07izisT3jCmQ1CWT9R0MN
vPhixK6xJNcim6uXEreCWg6aOtGwsBMmKnGBgLLA14iDh6+avpv4nJVCY7L6LwZh2Pt+vkSdjlRb
X1ajelDN+YqEHGkm2VFBgOlgFF3RpXcPRLytm3tJGN46hGRRM/4jKqfsXWJFp0TUiEFjfN9j8mmA
dmjvhd58dhXmmBIyldun5WxSa0N7RdGQHiyy9NSVY8YMMvw5SxptECsRdEopKDCje63aQVmYLQ1y
zMGjGOxHfmyTOuArbUH4f+gt+zu8oKZwNgfypxgp2h1rzypzrs0wEurswIDeso77gSpOzMLqiVGF
JSnxJrettmkYFbZre5sISgvSVAndEMWiC44oX6M8J2YpgJVdajzy44+uaxEP5RSFq+eLnNNGJa5i
EXb4NRXznKeUHMaLmDbnBqwKA/ec5phqla5/XAgl0rx+AG/zt2ukqj7Il/sHm4OmN9ftv3Hf7IeO
M935B4fPbvMuqQ5eEit0nBXg+uD/NNXYYbRitadeD3jBxILY25gn/2Z8VdyvlO0K0cgTDOPsczV1
rX8USU9yoT3nY4s46pQfnGcf6zdO4UF/FbHqRdA6sYMH+ObwUEPfA69cUxYtz8o4aC6mb/v/6KUT
9/8NBxerPVGpCx2121OrqTuzQi9n/FcOnai4+KIWLjsJ5r125yUzuX+rCAeGs3pg33GMvByLgqui
5ISdIqvDTsV+W/ngHyKfTD7vQLImMCkYNmCDBghDZIZXxM+dz8QCDjeOeFWUP5Bu942+Abc+1Xny
csHxqA18EZFtYceJJ4rMBjIuGjynyNMswntIaevi06qJtZDOxRK2grQhGp462WFCdoeTRmGw6MoI
Zspt14tz6EouiyqKaLBcl/3FJ0R15dCY9sEpuv1nsoq1nrW3mLMvHJo333Ik3y4dBKSBZMMq05d3
qPa0Cv922Xil3TwsvjspYNPsZcvtjYbrSWQPOK2QXRs5h7EeaPyook5zgACnAV8swygobi+3BbmS
+S9dJWhU9Wv6Z+//HnTMaFnJQk+ysEpXR/wOMKQeyUmIwE8frgPTQEyrHMuStDEGafEB92/BzmSX
4W3c2go/C/udQbtC9KQCXISfcIC17/RMUQIMFZM/hCMMVjL/RMcGn8M2/0Y8klA67yUo3ufRqFwG
9xqDm2KYMLsjbRDufZ7cyxBO5b5BnpkcFftALr+ToKe3ueedxpVgOMCmvnPl0CQBeF6nMR9qg4RP
YRFbNOIV23jjo0QQOKwFQj8B4IgvoufX+m2DNQQSuhsSjd1XdaCJ7da+a2zR0Oxv0JsnM4djvUSB
qVFMUx83n5ObA7gZuXG+hVUUuBBIuX3d+rdDeomRZYzI7Das1V/rY0x18ndhLsSjjP0xAxZM8Uyt
QxBhLXqGWbYI3L5zqt6YEGpiHSXZ6mwiQT8132w/hy9bstRA2gnHdxeZ0FUOFJnGfESFIwo8yoJg
os1Xq43idT8esrQF8mAScV3Q4H5b6JwdEtMlMmt7+0m8mlCy2ALMqlybtr2hOryD2zuhEpdJ9/iG
pkZBzsuPRsz7Itoyi1SnapfUi+dfPBugSDopQfcKz3lyUbrvUioOC4w7vzLG7RlLzT8qbg9XrNa5
AnZkhDUqK5B8Ng/7zA4z1JdACZRX5YGJJBM2xtTnNIHvgkwfGuA8k38UWV9vscHuQcaZKhPuPkqR
mH1/BAOhmptrVcj59ZZ9Ah66sfofoDTHfyiah5ikTXvMiW6LTFTv5F3dMck/7nRQuQKtkgfo6PSm
+J/4F58AtKYcIZ+O0DiDCMnKGkBde8hi7X5kdjWkUc/x++4lVYXPmXtvylMdzDq8Sb9sLWInkSKE
k/xePN815d5FNCEypE3F8BkdGofXKbDxU4ubYZhxl887OeKKGUW9wi7Qo7brCDtlJFQdAPkZJgb0
WI8e/vVqQF3jX/DVsCGgvPhepqtYQFwwyKMboH+s6F/YMPFq5IeTuEqSj+xTA2RezyzOC37LVI1O
um1Lr04QAi+obMR59W2DlR92mZofxGQ57WUTKQJh22v/pqZS/TNX0XfCtELV1FiJjNB4X031OGh7
bzRUk+TQVJ5GbVmUzsUe/XbUsFKBnn3iCRoysdzvTAVeQGRQRFqsdYEhVlf5NBCqacy3C1Xvfrbr
KnnO6er8iTSrwMXvlV3UYLUq44Q8REwoaBIlO8Yk8kYQu9of7fvnzaqe1cdeSmIKsmD//J59xyN/
DdKjZW9faMhydTfzXrmZ433Dku2hiiUrvLvFrM8Z0OM2izfbgpAFp01Oing0DtThR9j9m9X9l6jQ
P+ttK49E3IFavdwE0/Q0xoIkxMvh8kneUECcYij5ivwzAvSpe0dGHEl7NxvA02EzFYmTU0qTt1u+
5gkhHs/fzTrkWK0StDZXiW34WnKbMHigNPSVnkWwX+TRJcKYfhYkorwYkD62G7SnqVLedQHS0CVi
PJCrUCuPXLue9h/GLdMwDfI7AAqdw8l/NEICig0iQBfCVtPrCpXEB+akFp4QtzbgNfnQ3l61mNcc
gYzqjSd4QR2ChOPAzohpN1hNjjJX1IpPjTcrDChKd3IWIcjtzljylOttxM9uATJOnKZR13OYl4Od
L61T2cAmSjc+WfVribMQIVDDWEL1IDrAa1mRSATySqeZDpxl+JELGMW2oiFjwkNgZKL+NSUb8sDv
OsI5qY6xHnvoDuWsoM+5LJkoSGSWgPlSxVihVrwQsO5sMNBCAhKNhA7laPv8jpWy2ADNp6KvOKVu
eKq5W1rrOpaZ7B9voZygRBm5n86L5vAfGaqvbqLPDo1MsuuVn5ul/VVeta3gQT/lBdYhR7p1jaI2
sirNykquhK2klJpY86N8AtbqLz9FOLoZ+FY2RLUbR1+MEoMgWbQJ7mt5D/9KtvVnLyjDgt01LSyx
UlTRtOlI/U5JAR+HgCLkbS4muApkgch6qVB94TeKYJ4vJuhqrq56DZbNto6RH/d4YuIEMSQRlu0A
UhiicRlansAUrJRASbgpxA2aw72oJ9Qmhz2demWcR5NHdT93E4DZLSxDdBNvxB11V+ocioq/a+QL
/3AWOjuNHrcjko1KRYYcQLK9TFzC3xT5P9vOk3UvsuIceE8f5c3K6nXbmSqoPcDMpCxIBSVjAMG7
ZEJ9wTItyqO1nqUdL1GLelqP/cjmyOHr2XDg49sSFm4ZafJfjVVQTekF/4qdmPq550ND11O9g2Xc
87TcYoQMl03n7snCfaJIlNpZypdEFKtBtCbjh1zIoUrWl2BohIFjhO/w9aoPQZ1iNE2t1SPhV1qH
W4o4kr0wuuUT269HzS0X9ubofvx9j2D7A2OAt/8tCXQkDaBXWpcWY0ZrVUJZFK+sq47zbrxHeClL
XMSRcE+1Puk3d2TlUFgCWVxxdEXJS1Y+ClUkNA1LU+JA44ZQLND/b8b4PkqcxJUWvr7THlBBbZwu
K23iWVtQPAMIdN54ltCrxgsUhrpDYqmWWYqpmlC16muXz9M0suA3PlIti5G9hmPYure0jH8Dp74b
piw42YLpF/Y9A6rd6DdHPqAXOsMIJFHcgb9zLkrZ9l+vUvFIVkH21JeFhy5XaH/kMmA4Gu1pIe1u
1YtwzJc0Fgg5UvWU/YkUgBwxe6QgcdKDGCCeywW7fI+7xPSyLBN0fh/J7qcT1gldyPI4mGYyduDu
zKVncCfUOqIFPcGgLLV29julvWvsoBiybbIKW4HADAt94CBdvD8vwbIAv/YOz8ABv63cE7F9rY9Y
XJWGJIy68IQEc2ZlA1EoO+0RNIKAHJp7TE14UeYx7oN5B+StihZmQgwykUm1EXz+7pXp1nK7onq8
QhDM2crz0XOgfP1Eqy+HbBtwBNm7vP6eUG+Gyvf21pxRPZc0wg6dRUMUcX3dqihlA9mgFi5Mha37
5LQnNcmkCiBgQEfNGdwbARTb+1LUwT/ZirSpo6uVji3TLnXi4uxqTTVIpkLBlLpkenVVWVYnghON
+JdnsZz0t/Dl22lu34oJaddR1uu5eGk+3ZIqm5JyT+gHuidANEHt2bVSaIE8kHBf/S5fX6WVyPhv
oXOZo2TVn50id5WDpcANjthhbFDd8p5t2Ww0GgmgQ7gU3gk7RS+hvnvUig7SaoflJsaQASrTd8jB
x2TmMc7MSlLaXnhLMl86WHXiRDGTS1829dVPtYHUfUJquY4I9y+glPzcu5qVLPqX8DS94ucCIZqG
PJrrYybDt5bV5qiIDHWxc2sasGW38iudc3FTHuC+kgDmr46yF3Pc4IRQdX7PByli0r3tc+olu8ZU
gCpTEeZZpNuZCf12nICUYqSXgzp6VUwMyGvB2rsOalt5ba4IQcL6mQh/uZ/FNnBAW+j2UUM7fPZq
DuZARSVHSvKkDpUOHVQ68voBk7agvLxYSMG2wdL3rr6M/Lp3bFL97XDvjFf2iXy4JxJkBv762Btm
BDterBBuIgqajmSO/1cBNu6s3Ra+ZBNThy1dp2mSfVK+6QwFW/YVkGzEXyxRuUDk/BqXIp2qTgsf
TgGKRPP7ZMFlAGpsaGApYmDmNBwKlIbjr95FIEPkPycFw0srxGNXHsGmHnk649fb0TN0Ma7YcKK7
kdAqoGiyHn+Giwnp9A3EJnO6q/WPNRFp3bdw4nGj4+L1TyojvilpF3O+1AdnRvDSklTI/OoKfvt8
ccAEKmKE5TyqcG4XQnUdYL2GqVZ+PJ5lx5cGwYFhPtlcWbRbnrQ4m9EqgZCxWnxYT6598KRbDyYX
6F9KoVBI8uj47tkJfVlMTW36vImrB0hQhwsZqiFDBgAUtA/CdbL3p+5N0MhkMY5DKcCurE6uX1AI
f/JuiO57eTiuqSENXVpf+4XW/o6FLTSXt2Bu1TNNYc63i1bvsS9lLWd6YLshj3mK3CWpGTEb1hL8
Hbp+BFOhGUDqt7Vf8eMWEkyxvco9nEX7+MzWJBwTdzvlkJ5nQXx24WjGNaN60NgC23H082W7FNjR
6IsZyJr2YR6XUXMNc2NDs3RRFufAhCA8fxK0MneiuUhYQdEUHx3pzy2/PQVNfdudjVw6tGx2PL+h
hqaGB/A3PYoPgOcW9q3TjlwfZjdXbW0jvDZ6gvNPM85lcDGOgKagtMHVU7E6dORqf9FwgRrs9y1i
uFC4rfyOaRV4QdS6LTEEgogljDjSnd2eiG3ytmooW6ZRW/HhhEbeJhocRpiZl/1RltyQzzvfMCFy
g7kg5GDqpO1Bn/dUvU83XRwNYVC2e4T1if+1yOmHY6fFqZC1Sln/kl+14VbYvBHj84fxshG/1OBX
qFq3IzFSk/SPiZK086RbbFft1+K41eMqOPZ10bsZPmn5WI5Fyxqe51sSCPEOcD1jqrMtjHfXuual
mjcn/JQ5BFdL9e25bfR2eF+tFXv70fH/l9scYSJzRknJFIwGcLrW6+BIuM8/QHASd+7VPgCLc/T4
TW3Ve/fG59zBHvs93SeUnVWn58BKmF8wIk5TzW/nvakSnq1vP/32qJIMOut0+c0td6X7iAroLXgl
98A66scsxilojwSlVzKGXCo2/ghidQW7vztCe32VPq0hV8iMMaMFyMFvH2/dz3eeBGBUn9kwwjui
USkgNr+mWM8XSkXln2e3ZsJS1e7ANxKGxBaLcy/FBmS2Bdxapwr+O8WVpFd4PHKI1nmYWmJSYNgU
zuVBkSfcckhN7J5xoOzxWaGWQ7eGxo/2u9Nj282fvRPOld8n1994p/8ZRySToKRkOTnPt7iZ8s/B
RIqA+ND5nObubkQ4jm4g0kV3NgSCagXTvm/jdzzRbv08vS/K0MCKCsmjidATWQxgFybNPhLJSmxP
DJQqzBOVDRzAHZKcetz8DOP5IQGljHIG/4cjFfN4HhWz0rBpl0xSm9ps4B2UHN6Qhz6d2UYNXouN
iwbNqQOPL2tKN1eXVGdpTtIooSM+pRmg7DOefPheW3XBnucj7fAwCO13Zu2BjbCYCguMNjtc1jeX
9G0dR2HSPwdMZZ3+2mEc9qOqupLWVgBFSPZWI36Z2YuDnst34pIaxRg4qOn2nbaZ4M7+4WW9J4Lk
J6DpNrX7Holn6vlFin/M8ucTU5xyJ7RV7/RBK7pwtKoyzNmjEgcPJmCI+ECzu51dS4cNaM1u8Hof
MuOdodEjnflWSZwMwUITEiXSjVQVQry4dvSYHaKOMYjwruEl6jBnjEBgmYXMMjBfrez9pI6D1RE+
073AAlAr3kox8HRBkN9yp7DPhzKRmhK5QKSF+KM+u+WY7nHmel5G6chKvr83rQW5kAlP6hHM5exh
I1RgZmGvzGLFq+WOcFNGPTkMC+6lJX/9cL0j3RoAbkR0/XdIF/kgvylsatUPqx+dVEDTZX1tLoEu
876Kb4Sm2BKGADt8McdiiT+LZJHxsZv7TcFmy0Qs3ZqaZ63J3HDMBAhCdZSrp7iRG5XuuYLG2GAm
NxjdZY8TfNMbWLVYT/jKvBp6JL5tTngs+EDLsjjdnQSQ/3XmdEe0xWdwxpYPp/ufDYR/mXb1KZkE
7WNj7o/4nnSlfHMaCbkT1Jr+TaQbt0X8x7wo5dCKwogxhmJD1+waRcOc7cw+4rodXs9UMsgjxMEG
hEl08xHARP3oHxN0OkjeGxzMgH1dN7ZR5AXhWiSTLoBqVGLcLdCfmtVtc2yNxNaV8YztO8hp/mD7
Y2/R4wY0YicznHSDOtxfw/NeQowPCvZfLwXbDkacYkX6M2fHwRTwr4nGeRnjUd2GCVS8vQYY+p5B
NsUcI38NWlcCmpkYxEZ3PtT0CsbnETqLjzalrZ47S/UiGO53ihm/ODdsHNDEws9/DEQ24SJQGHaZ
ZUnG8oIu5eCiE5zVVb9GxJLwBNSUCG8KlE6vhqMzwSnW8j+RU6Kqv7lKJeqZwL/mv+Al+C0dxVBI
nYudDYG9uDKiVfFekmfWJKOLWwlbNHuyTlM/8RXgfbj6W5sMwGnaEVJRCzl/zvu+bYFNDSElvH/7
h/cboNflVhMFeyCpa2nxWMPEGDfZwQGwRWjIjY2AHx5Qcfw3HnPZgra5QNuBKZDyIMWz7Lu+59tT
zOcSG8rjCZV1QHh67FVeQiW4ES8LJMTTJpxaioQG2B0ctoj5aLLRPnPl4nO6QY0TBgVaEsAEFpt6
iQHi2v43z/yOnh2QFqy2idt0BUasiNgOAVnLARKmYlefPJUpyoiAZs2Ri33dgCPusn526xHVZi4F
oHK/KU9KVzWtQG/KGrNVU/gSxbM7vkQvYWd9xIlv6TbqeqvMnJp0K1puUc5AOtVl79Pr629uCBfr
hJRcq2+6KweUEJisJRatjiIEzj5uLcw7XmA80BcUfSbus6equTXWyZUt2v3jtcUPKdwlMyJtSCuk
8OQUiD+d3BGz6boBx4Fu8EqrXoZJgdVpu9+gbRqXMNcXvll+eoCyh4DS7hw1jD8QpXMJGPfcwkx6
FYnVZ4c3TJ0qzsMPUhEGfpqyWikQ1wltY5XE3mmDFyAleH31Ht3LlZk6VFqQZFkNQbo97wgDFJ8k
gIcqO/nhQcDW1YcQAdmled6poq4SevT+QT+3sQnhww4udBZz9N9mTA/Gxqfc9o9V72DAUghznPky
lerc2ySfjczscx60zMUah4ENodnuuyXRJH92PLSUOr/YldUWHDGZZL6PuDY7HxVeBoEPDUdVhRP+
jEWaJwoNjpK6FAAECd89MlhsBdncKaVcqdEh0VSDU0mOQ9EROmEJbf9WSLIF79M+3bxDp5sOy9EZ
Y5T3whUOySiaC2j2A+aBskmhzfx7w0s7kO1960OrbSuVClOPg4IO3NVON66MLRCtdyyQ22IJcyLS
gMy8i/WuPwkNMKDpcqSBFPeKBKbYRHg16DyyzPfO9fioKRApDGTjHEXpLhQSCSeTAiIbAcszN8Yz
N4ZpoS6a5SdtRSqNzYmubNAAimibg8b06BxI4DvscyuEJXroBePEwVekIQvPi3iFExWrKfxlfm7s
Z4J23FAtpZ8VTk+bY66ye4H8iBAx3EenmcX3DEMLH6GQHF65Psk1CWIzQkhTsf6Kdc1vlANQHeNO
Vxxs11qHIOMrJOxczcCFzJ2MgX5lyCuOpO+RRt1Pl2Q8FC2xc5EF8uV35FHXEkx/aUTDvXA3CNKs
OEgnJjBD3QaI0Q6lya1g8We3Qf5BygvuRYegqrJZcz9u3+VfLae16kPKUm6TZz58y0+XmAE3QMg6
+ZFrFf3huv3KO8117KDdoPG2XXLdbkdO3JYTTorq5m82vgoYnFsId5Z/9AEi2h9LmdQ7VKMmsKns
uBrWL5EyXCRXwbzVK+XPExidyB2f2DMbBrY53Ox5queWWG/1gtYerLXLVJ3x5+xTvJJYgC9ZRAG7
v3FnUSBj4RcPV4P+WlwnZf67TKRw1gVK9uvINe//mvMwlp11D5O8icwWKi3Mouvdfa8Y2i+fbmtq
ZFWH0QZnrY91YpQkahYHf5xFY1FzV2XmDdncv2Pdw8cZ5fzofO2BOTYWf4j3gmNLFZkTwT0b3+EQ
TFlpExbU7e1OEQjZDbv6IcjzG3dwYKUs+ophxfQ0Ik+NOKuYPdVIeQpifNVRPGhr5StfXeZa1Ig+
jW13VBM4pMnDea8/HE1p08TKgs++wt8CFqwEES7RDS2M4x/2Nt4u5lDPHKPAy4kY9lmYXp/VTpot
+iJK9uvmXPv9eojHZjDQ5cyndmqs0ny3ZFRA5Bt1WJiKQOsDZRaz4CLmEPgAGwwdZ4nKoJCKOVWN
DAD3BjxBFwEAc/TaSqQvE0yjwPHMrmUOa/LsbL6CXyABN/3Nyts9+SFj0t7UOvgSKSatJ9pfaTvZ
8y7mjYbDJ5sJTzKb12EfWmPehkldbIq8KgemU/BS9HJ5gXHy9r++/yAnkFRy6EifwvRVbbZIyvSI
BvEyPoRweIGt6m3uCnHPbuIpZ/74Wg1Jgd/YaIK8xeFuSnk/661WRvJzEhXmqSzd5lCjF16jg4f7
8NlOhTjV1XsrEl8K4/Gm2l6gA7Rp9ZbBOV0r7+tfZu0kjOZusIPnc4geViZIXgEFv4OQJHnC7Oei
IM+ixaAy90jX3gRnWEA6jtyVoWDHvZogXI54aElswiKzoGjxyzsyFC+qjQuSjR0YOQxfSHKs8Gow
HY/hj8FkV9KsSJeIoSIdFue9SbFXkFjzEtr2dUTTbfLGCXj5AMIl17sWzGmUmCC2LEW4+rQRmKoS
D9SIFZe3PjXnTPa2DHAtanQBFFg5XXzBfwY7Ezx1ewOGgtlG4gRZu05MLzdTFbdz1PDpOtTWC2kq
XM83Y1iRG2uOragydmSCuRsBTasTRsnPAxii+j9tWfzP0JxT0D8YC6FzZiJszUyUV0dtLSXgHWpI
RbF6WZECpA+QXWjgAHh3QhVkYE7zzqKZtzKYT9TAY9O2IqRbP5Gd77SQOjHrhbKxdbtKnbisp26v
xntxqJ6soejGgjCn76f3K8C22uy5Dgbi7vL27EOIu2mth79S9Vkw6YaOZ5CyuqI57Bp6CqJYJwrs
QMC6gfg1XoT7QswkNIPiAUWdqJyu5VvYxAbp1m7FuLUzrMFUX+Ykw5ziqMYCZVd79lBEWotwRlXV
jVOb1FnFZGQBw+BmC95/FWmeoxVdm/hL6Ud8K2g/Fh8Bzmzwqx2rexnMpUq9hjCoJA3Qs6sxAs8Y
WlFM5iXQMxLbuFLbJVFWpURvA6//9umibz0Y9RpdcPBPdyjecu7L5w8jcj2Vk4hhVf7/ZVkPsHJm
V1L/OHlslPMOediwJROORlrjzxuJgD3yDjlNhtPg2839bJpQwu/dDkmii8exD84GsaMGVg9n1wSE
BLrhFdAdQFG+6rmN6KggkJ6JxAF5nLzQyimMgn/GEBJu0oHdVadsbeQvr00V94ObWG+3nRJ+vsU3
0FJK9LWT3hiaYpRyiPYrcOZ3G1y/t9K9NUaTL4xOR9rxASSGRnZHAiAWfmxy6gUA/Yg/HrYZqMKr
4/fFFr60YAqvtK/u/HcXrEY5jBTykIVj2MLKGji8Wl4UhpKdRC0y86ifywvmfr1RxNevB1RLnyxO
KsOswt7ayslKVmG9cDuxxG3/WROQfYIXfj2y89myOoakhjueAWLGS+Z4rRkIn8MyKL5H3XuPgjf+
wH8Y9uv2OST0nv4FvN/F49kEN/dD0+T5byGTKusKZ19pLaT9jfr2syVA7dmI84kt0EqBQ7SXBsv9
sixHiHOjuslr30jNymCzPsEnh/DUGesWmu0+9FX28ku+HOegzPy78/K0q3C0roBMReVT5t7GDpwQ
IXeWIB0SEa/oSUXkgE6+VZGm3FW2kRd+75FEgIbvqRxqR3tepcoV/BjMDGNFI21Of4JYx31S0ioN
QWy7nD00jEjpD8JaBDOdTzhwAQtWBqdEwjqMEwkPLI/feDm7MR5+W+UGVE+a98tyli6Zos0dZQ6F
nmWJknUuqvVA8NjBBBzr9bsr5W6NoSYg/xETWlirP4PU5Gi/98+2HVfZC8lSG6F/N7rDvC1EYQ+0
U0Np0XsOyerfHNtxGc8NsvC2X0CFH9Qv1aOR26v5/LCUGmAXMF6Y3oOBkmzPkOboBuG4xL+w48cN
fyXDpGJTTK2Bb/MtcBVkZ/xipmF70Teka3NVVsth2e0F7CIGkHlXlUe3UcbTWQcmvYun7iCqKzvY
7Yqoqsm0BaN5M5PmYpNfp0Lmj71k9sNG4xtS6lKKpjjWx0HK9b6RnOfWB2lDoyTTeH+RdNmc67Ud
I5+vra3V/wBstyOcTufh23o6S+0FO17KOz+HfqrVM5CGLmam0basoxcBGV2j2YD62W/I0T7CXyfb
lG/E5C+8zsI6CPg0e0/+OsOgzP3G5JKVWkFunNVmHbCFGfa7V3dibkYi5i9iL3CJt7h7TvtLhNsk
9oq4AtMtijskLsjd9v+z0TILMFjJi22bOYHU3NrJ93oJJWHXj5LW5A4hgHJeq/5sxkNVvUpS5X6K
KjDdDgkG0PbAFwDsQ9y06qLaunR/f2kBait38j1fBFOTG8VxwCDQiS3tpLjnLagIAWdO4Y3uWebv
2K4FRo8v0H12R5yuBhVT14kPS7XpQz3tBoLtF7ElxCqh9X3+jT+gwdfeorxyLRzoxynuiVgnjLz3
LRCSUwhVz37J1wUBS7TPNqLbkbXAAIgCx1fC3gGoBZcmmWm+6YWreKSbYWFv4WEtTFfGGZg/lNlj
DFvIPyc0gx5whvBobj+pTEVdsflSy5Jrz8Stj5ug
`pragma protect end_protected
