// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:13 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mFZHyM3oXtfqns6hd9yS9LwoUXPXy2oUIA1Y5tRH/ifwiqb8rMh9hQQ6FDVuY+me
w/Mn5Aes1NPNERsF4NmuZcJ07oOMSnpYq9yunRcGI+wKtikx7ZRW+0Ie7OHYiofr
1A9aW5P1wbCdUgoD+1Inr1NyOJqVgjSygzAO/MPYPLI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11184)
r/6wLqB8st48fuqIujKV694kuTtJw7bfZDKIRdZbumjBjdV+995+PxtfCUyrUgnZ
JKa9ozVREquodTZUR3TnyzNI3QHlcYr8iuHUYkKI4orCVUfTDqpkC1GK78byyFZw
EOpq4rRsp5zr72I9o5m3gjvuQSeojL3+ymB86e4+pLMWMN4g1fiM1QQ6pXh8CEU5
mD8GlF+xeC5j0FQLWpQ48abxzgKA9TMt7KIyoQqxS0D4VxTPplKOpoYAYNuSSefN
IZE2tx3R14dCg4CUfNCX5oCBLAEi1Y3NBs+FQajfV1z3pA9C0Ld/ofCeZjtSbU+F
AViWxhnSctdlSz/aRG08vVeJRg5Nd/uFqeZCQfH3jBcubulFsfMSdXPzocyaS4tx
TeK7UNLCTxtgeTjAvKU5+p7i9xJ8QD1jHqAqYmNpUkcYfVTTRmNJskmnYVDgppj2
rBQQxgN6B6FEce12zT2TC4j0qZAxSfbWQkK3jeFElPl0KSrcYI1G+fUghZPxbez7
JUcjIsGN6Wg6U1zOobn/HCVXwm/bvPA8m/pA6YuJAAHa2oiNQsCjfCUicvmuvsj5
+4pv3CtgNoTtBgaPV8iKv3KoHueI8we/po7nEfFvmEyo2M2TzmjYhbSpmAqnwCRv
qkSe2YFTvP5cigdCn7xQFgQW+yNP1/QFKCKbAWRb3W6OpB4Et1ehQC+KKbz2l8Jj
wxJ8q40O3eoNcWxKnFmfVJM7EPbTe5kEcp0oV/z4ywc9y338USVQckYe9HyIEEWs
alZFlJ9JNX4ZQglJyBoLmQ4ZKtmeBecR1DyPuigRWA5dWMmUCNOfsefXNqlD7Ti1
od4bFz0GoQdEr1VEiaRmIN5Au8oxkEXQfWbC1udxVJLiniicnpy08MkXCJqN0XBP
KhJNpXOeLxkv8ibFzDgDT7CnZYEcfN64ZRFePYo75/5n++hEVXovJpkFeFoC+sLv
Vmk7vYPBYWMk7qZqQK/+qCJHEydmuuiV8h1f0yjhOg+ygAM+Q6bMXTjivmus4ri2
93Rz07TCNmRl5FmRo5kAkZarLrZ5rd9cHitDEpd/nKhy0vN8RewaVxhxd6gZYG10
TVR3K+zmEq5HUdyVB8hikhNKV78nf6iXm+mW/meZ/sXTwWNOMKZ+Q3VJYO7tmJwA
iWMIHNu185kvMEQ/mlKCNI98aL6DfywF+Q+e4tFwDVFXeqEmtWyqkWz8w93xvrM8
+lgp8lHCXenHBYLdFDLDIXxRyg97bVvucP/xIjx2WpftWycpOYRreOmXQDusVUYQ
ncHfDJkFFkBwJuNql3TzU6PgSvX6fY+Hmog8eNgosoRjBxww7COBmdOM4QAnki0p
zHv9T4k32UZ/tU8FekDvs4P1P7OPGzB9/bv4kPsSOshyfZXCbWDnMhxHYpl1yr3h
FuSown7jfd1V4jUofyyCRJNYjNkoMTJq1r2tTykjDcWGuqczv64H6rOlZPdobQCn
q+lz8KjOon5MPudtDX+03zi9dz1oD7v8nsYKeIxsyLwhMTlon2bdnw4/yOtzepEx
dbcFsSSdLkT3rGjBArLyhQs3lcomGxECuul2FvAH6kW2kVrX/ducuHybZkYVhm16
YqGAJNqpBncOvxGrU6q3FtJFOOKwdf5oX1NJ0OJ11p5eascqmVnCHI0giR3gp2rc
O8J3dgyJXHqSUO9M/d7aOZa1g14VA7RFcJ3ybwRyH1mM8Nu1I5DTvPwOodP21kX9
5GUa6DfTIFMHq4kL8euDcNkccywOidY0T5mdMo6aL+oQKjX0s32BcwdS/WDd+Ceu
G9U1nZojKO7OjXZxJBbL06/5Y7ykwIMaWTDui0e1movT9fCfA5mTSquEmRNSASmo
eLj7YZqKiWCl+2UfwmY3eQ0FlGchqSuJlKN+7PS7Vrpm0x6gWKiiRxU5C/3nnwXk
b/jTpCpFrCLEBEUXyNIcM6T1HIObJ37RQ4oQFSsSAYfKQmcLpIs+S5tVBloUrNPn
J5B+7U2IPs+3LFSKizWAB99015qSlIKh9r60o1YRUhxHASJIcPE2KZ0XC5Bk5AO/
L2q9jG6+99lKOdK+twp3Ibis8tOL5BLBLctX/trFC7/puThMIbGP1NzcbHFsbMkN
9fkB+g1IqKb8f7sCjBVqjpTMHkJO+RuU/NHb8Y5Uwbdj661Nhkba6jmHgxnecd8y
HL4lQHyaLRvbYr1EdQMuEDCPMVI9bFfoZDM0/VvMQ0GLXj6mbuEJ4DibTvStEz37
/qvHEyz7uZPyx1hu6FZpG5zdy1ilwXSyMCNvkXgf5KTQLuu3QY3vG/3pcMo77Uei
9gdFvsrryjNT0/WKAdejPqSi8mbBVaDJ40EGmMw68ncnRVAW8CUHPiTErHCL912z
KgCpfFQ4vmzCdqDcmOHIXvBlxaEsrdzVsvIT2JfHJlNpth2vbrFYEg24pjyestK9
QPNcV0A/d84t6MNd43qYwTsR7mUasCmOVindqy79vpTXJHjzbrQoZiRLf2wEhgR/
tjBC2wfSUFtAYIbWp34nH7N0WnxJ/wCeJ3uUTIzKQNSW9yYPT6WXF7x/uoQTmBvR
SBwssRxOCCi+SXHZM4FxvP6G7+HKi5fBfWuV/i3iCyulANNnEZsQNEg13rSBw/qU
jkeuCkMi8ZuOFCpfwhbtApbqy4tRVrv0ncyWXAO+cR+otkGX0unjFvyuaPOnoDwv
4tndpguWjIfy11JB+B9UBTulppTzSvs0ZDyQDdSc9rQfsEfbCne+oxIgWU9hS7Au
XueXo3txIs0rlSwDJNEHG8Q9EK/hlvkf1m5LYnMH/4jsCvODWC5+dJ/2qhbCqsXS
cbmv6Z9uqrPxdEKHn94xjQm5xWbddRnXhqDng4Io3gwvPRJp+THJcDMsmjvA3e6e
3nYVfFHTNzvc5LFRN6s0gbuIWpaBSiJw8pdcwwqOwgYqleXR/CcHZoBFkbnoXQNM
Dd0I/K6PJTSIPw1gC06ndhkz+20YJ9ntoEfaNp65wQ0vWJSxySXAhT1Sa6kyZufR
cU9JvS4nf7MTBNiVSE7PK+AjkiLD0TWqiSSMlpy5SMO0jdize3XsNrdky4UTp1VM
8jI/OnFyscNFcyUl2n7iR3xOd8LTcttvxi9kFFTQV2ycXdYM/wz4h2qTzjHIIAMm
mRvLMks9BhtxANvIZdXl/Au11blqSDFtSFc1HZt0LKfznUmcnsD3q8pUiFDGpv26
qlfq03l0G9QFeYBlhSm3UofO3Paa6nvngfrBT1O3KIQtPKVHefP0ml0xKzvvp53b
4bNV8oJsbzQsK9cUMPMCnKdTLZiTCQd5OMS56dpqAeLj3ykMgtfP2pECh6KoGw2z
gv7HAuJNsnKjxClbrRmE9b7SnQHhjbHTVBTat+XM4Lv7DrA49H2BI2SNaM0w/9Qn
AHaJYq9/x4BKvnVW54tWgWOW52cXGFnkq9wLbCVDWbNRddp6ov3DGPMMmHG1Q2DG
JVVjr7Cy5Lv9pZpZCp8BSXSTmp24BLtnNz/vvgd2bU966XlZL48RL24iO75WTSdt
7JQKwuJrdY5XdBLjiiioqSKuTc+qi/Vn7y6Au4q+30gfswY6bUFAsB2w5nik1Kx8
zPr4sFGYlCKp3G0wc3tbie9rNbozn69Cg78ZRz6l1ufILqgLDd+Tp3jMI5J7qcL4
f75lqkd77B3cE/ZVYNRp2S9rPq8Se6I0rCjzjIPNgLTVuSy6IVUeprURAx98H0Nq
hWytsEMRZK4iP9CGkrvYB3SwrQMT6zYkEx2YFk13J/WDczUB0FMSOw9DwYnTe8ii
9d9Q8Z11dPNgo0l7GeCbwhA417O1G4YxIV0V1JHhG1x6Menl1hJ8gpuRlmmmEkwW
ZGKtTGAXwODbtUEtytfyjQqzWxBg834wFolweCCUYveBXMpy/KBj+3xsRwjG9Q3A
0iV53RCAookVqEkuuDrL2iHPa63lT0hbA+/S3HDXD0mPitytwhwYwZeLl+VA+66r
EYdIHqpUYMYOqRmNrSejRYGinZFWi2zgYOYR5jiaftNfpDaNTWkT5t/5bpH42Sn3
8iwMjH+2bpDK2/CKYyE+RGJHDhSl6A5rf3Y07Ygo6mbimyMASHSa4XcEmWAa3Cnz
jrPUATk2/ZIYIa0Vdv73urKiY6MPv3ipBJVP1r88DO/yb8pR8gpgp2uVQnXEITXm
CIK19jH4Fnaw0kp7vVXg2Vjzs2BuLUW/Kd1XVt5xDvZN4wQRFEEgZPuVkECEeKgG
lbWGxfj7R38NBSXyoLEMpTSjq71ERqqKzH2l11/ZOsjwV9QBhfkntYU6oA4Q9RJ1
79sLgPeMVGysra6Z5eDEciQdnSzas7QRbxKuIXcW0FvnJNBqr5GRnn1cbk3tlDLa
2sr4mjJnSMRPd7dQr87fYvqwDkPYqgtHH+A+FLOwDsY5plv1FLqssg8Z9hKHI45k
VEANZADADG7i64LBllSnoQnA9J7ZfgmwFXU+6P83F5XOj/7aTCTsF6jAwai5gZQc
VxxRyFBINeyweIZp2clkj2ZdLA16YaDnJ+ql2BAMiXmIoRzkAB3wa7d8KShDZck2
xfzvnHpLSBMiONQJeWqFDr7bMxMhuWgB+I/rBkAgezhcVEA+AzgG0mIkrJTMDX2L
uZNYi2/Zi+Xktg8ktSREVDP358+ewwNRYeOMEn9Z+WkN4kfedE2w1gJISmcjtTwS
caTw7RtrX4rjMLQFUHH/3bHnMSXi7D8tb+XZnFc9vG64IBnW4tqpzDdqVkLLAOAu
YIGOeB1R+eybG+LcYGhqaQZzWnMhOkBkXEOE+qBojsWK7B/uC0U6xO4vcyQYrqM9
8hI0RX9VLOo57ir8cN7qmgici6ao4gCtmEL9L4hkxNLtOSlk9scYwoz/NjPPGUKA
CSIV4RElAq9sY2mNHQRwaGFnlze9uKc6XQ7dO/V3ENAWi3e8CzA57EETXMxAvRlj
b+OLzocrCs+1jQf3vZqqn36twsoXhp3rtIBxTBzQcEQuGTG7G2dG33Eymioyd1wn
Bl0QUjR7a35S1Pg2T8KDE11MT0BHUYta+LanN1DbBl+BX5mqoL7cfPMIjuTPnwjn
Dvqqq/0C43CEWbuAePeZ+1gUKflxGoxtVk/DlGt5tEKFfScfgUmzCIAuF0bYdfyJ
hx6ePDA/PxU1cSQscMknSaGVMkax5hcFbqeEKb1nSABr3/GabHaRzm2CdiI6wWV2
SYV5Ff2x1I9lGFv1LLaNmfj4+P6fEQAb8egpVgUhP3xegZevNZiXhU02nOhorNJ2
c4qu9Qsc4tAvs8Cl9QuGKbL+Qvja7pisIQn4YTWcOyz1x5i5nmJRiHqdII5dfLkC
AgQMHW88K2No20v9YRyfFABF4MWoK618XGxKaHrXu1oku6KdmzYFlC+Py+B86s8a
8E0FaPEXnovCVZvLmgxWTiU3b6OgkD7o0WJXODquLqCwNu3hVtXKZF76uF0UjJqA
/xy/1njoO4gxo9KlJ7coQjUARTvC4S3iIsZlxMhuMpHNau5Je/49ZBnB57b1ou1c
VRHzNPrl1iWBx+DOfak2ZvcLKvfR+lw3nxofXzHJH/02u0Y+ZdGQ+930j1dkJwh6
sGnCafnTDKzt9vGO/Hel0tl6E6M7fdKb2L3N1qPpW71Pr8gRHFlixaYHqgPbLGEN
vNHM+PO6NO7qtv3zSLZSkahhHCqT9DbfvtQ3MzGGxDKk9eqHCXZHmwHdL269a0JV
EiIqT3IQn7THnatf58cH/XduSESPmXWD8YKuqvG9KZ/GVGpTC5cTvOBSsjnUb+R/
o7UyBtZl3N/4jtkUYVdpF7aD9SN6lktexeYbpOvsAmH86bqzOq/givgALm3xcQBw
JBYlRMcm+7uR2a9nEeS2FW5c1QKEx2YaRoOcTg18L3V8TlgQ4n9+NXk76Ii5NOrm
wtFlCsny1qrEPrDReZhDsZlqpEs8AQ68dM2rzW587qXLZJ2tlhIPQ+9ij0BXjNbV
UUYRcuGEbHaiif/D1gwTF5nvgsQE0mY7Sxay/NPakC39qdboIhwI7jZTbxGl0Eiz
lfbzm9Fla8llBqAYVkeVzOSorksx6aPaVJULHhLL45nzVKpoRIR/qy4SYVXykr19
9aWJjatinFcdaTXY/5FQEm8Pz7th+m67GBd3nKwGP+feYmIn654FyxHGyMm423Ei
L4xals1qP8QhHV0I9eWN6nhj6gJEhUdfcy4Fgr9Z1Fu5/17cGZOqfTE6Uqn8GluI
VFpJHJLUcqGa8HuKbVDuJvszbBa8Th16kTpqzNBTpFV5rKApoPfXNTJ3U9O0mQu5
ARO2phtgaeO9TL8f0pTQIjiR3o4KV7/hOh52YYSL7Jlp+ezaQt0mAss+G5zPQQlV
K06NhXIhHgd/qH7+0bthxbzyqzaRjQr7MZnOd/UoDo2a376asotsvJUK1ue38e2D
y2NuF65VMtfGHg2MhuFwvmONiyZRTqHFzWSrqiUxLvdzpXJbux6k1SBFbP89bvI1
zJ6VQ1fHKuFVFyNnb9VAJPmsIxt2EU5RT2o4TeF4XH0UNQQ3OMdepW4B6QzZDny3
LtpfgB8U8eRXuGF8Ycki9zJYDM/tcqbfskj06jVgbLZ+dasN1kjUsPkYVrpxuNzZ
Ll+nhJGJE3neETD4t2gRKutmYAWK2NAAdtczLVOIjkcdvmHVmYHKjl9dXZzbv2X/
tdDFpND1eMQ/OR43M7dINw9MrhN1gOLMKYiZSN6PsUcNwECGpvzei+BqaaFE7MB6
UiY2JK+/bAMERgjKJ7eLppaLyjNQoHnFpL4cCMgA04fb7kfVDTeKZRApWfL/obP/
BDVdH1NR9UBYel/hYkDEh485iySDmB96+OiJsR56CKT+9HSV8eq2Kjni96qkxAS/
ppl3L4xCvVhyd8pHjNRn/yMevdFyQB7bnaS7QiMUKbxvZxJWBTHDt4E3Tc2eJuBI
Whr/d8u9uWexhkiVcYIe7KEKupOzbFklaT3x13h2izsYMWocu0T9/eIsjxP0hM57
k5wighLrmhb3Af+NZyCzx7p8psGjCPaBqpyVvB/XjiAU6p/YDAvUFNhNwoRth4pz
Wf/08HnoBB/WvOQhAvx7rgqozYnZfs8l1JMTO9/L5kT3g7UpOpZIFQmxYv/fN8fA
n5b6v0FLCsclEemxIoO3oqaFFLgIJxr+Igs3+MjKOUIjXJ+ICSL1CxlSNYQBGZm0
wSFQBZZqMtjL0lXCivDSnjsw8Enh3sgQSLwf4ZcjhSIlOC5gWjSJn515qZEmyG2z
N9YJoVxzgHz/X7mPmwYH93NuYjas+Q8cp4TYYQb46KfSvSKRAIBfWAEeYqZwqSjG
4GJaZlUZjJ+Sw+cJ7DRk60XjtLgN7cvHUcll8wvh6jUpNMLZKf31L+n5q8pS0yRt
QYIQLPRoom+UvF+QmFn29mZRLQ+ORkrZjX1pTxLYsakQfS9tiLdVHE3IM/6uCSZe
uNDhCUcZtkHn/F4fhRAjmEGeRIiRvojT05pmwgH0iCwRgb1LHcs0xXVU1qsgBx7w
xnzQIVlLIL1T60+zTAjDUavCwn8FGKvePq+vRI2kKLc5FlcP/zUwb5u11ZFElIKI
pB9v2WzsxN3HWmMM0trbphX2Qnen21cub3+pkDFyIx4DX0jAc0LPHo3KH7oMJm50
tHfFCLUsi98Fo4NRQCOPRTwqW6q2NB99ImEz2dxHt85rWwC1EV5JPwCyOjnxuZ5D
kz6PvtvQRK2nUlX+HSv9IkwSDYRP6+0F2aowI2MEEp7Iv9yAhNMq6xJYdk6YAUFw
qbc+igVxNdXNKomwCHMlftHVEGtWdmAy1b+1rWN/qBaWeuzsUP7I9DKTDKbIC077
RmIK2r0+aX/Ka7m2GAAPbiGgNqXuQAvYy1w2f86brthZEtWnreQcBLk1uUyb2xiX
AV40bNVDs16LiEspXQQoK/yhG+6ZqTXLPgc75F+ZFz6JChCrKW4uZBLmDuZrOssg
b8YljbkZTZospUB4/c0utVy+/cCuQ77tV83vTllCNbU9KpWoq0nRT1cmQUEaRcJB
5voHkOXnOEYVo4N72lkbdVw7Y0N2uoTISRqKHh1Y8E+Mw2oU67BvDvvqhJIQ9he0
w5Sb17hL/eHCveKNXfHybhgFmgPi1gPlyU7poz553JfSY4lOBpbwtg1GZPT01n7r
pw2O1cxd8txHw0ISVtrsjP9c0t7a/2jSxRnaENTPpY6owyEohS93AegzjpeRj58x
ey2tC3170Gy5hix0zV6XDASU1SEwPekV3fTIym7NugNpipcM/aRbZtcpzmz2oeHY
uAEBi2I5rEX2zP8b9EB4OhAQ3QhGlFqmzF5ZMCVpFGC1Eiz7bM6xUYITlS97e4hm
vwEzbPipfKOcVGF4BvZ50MhzIRpvtuqkpPiaVgdCjBS3XWMu+R9fIRi/71WbtX7b
bTGbdLPUcbrnemSr5DfBsSyfGflXF0q/rLfjXxMd/5P+LiSmwLxCRaApcjQmu6hR
6xK9Uw96zKTJdVajhgKC0eWvKgOg1yLt+EjKYI/HtzcpRm8eNkZz3uB4HKSEsgx5
/FyrVoDasznfUxDMKd3md48wzAV2UAcw2rBAPWvBaQnOyKCZY63glwmLIp6R990T
ADdCPbshGcEFQfH6aXj0Jw/FeOvXDcuVhF9k20w0T+0FHOBiXf1PFP5WSfc1VsQh
vZdU+9Ut+BOxMxemmaOd0zWzYBgIA8TisOnziQc5U1T/m9GUxLtSo9XbvHsh/b0B
2BQzKKckgDuqfinyWuVH8iBg+N8MYNy/i4bkotoVhBDb3cSl/+axLP5Lx3Wen+j7
zbFd6yVmEREuDLKILP2b0vGQQSIiBD2rYynuwjN4LC20itERucD3WOGdm8jwtY36
TZCWOgh6cyRY+dRm6XcHBWiGkC3oqQgHdzojslH1XHiLvi8UIJpmsN7x5/MZsbL0
6eRn4yRJ1tPcjg257/qPG39FnYPRsJT7Fswt7HZa+qvIEEnwabCRciUVSYjl72SH
o+QqufqlbSLj/yuYY3aJX7w1Ol3Eh9xUgngyE7VvTyuWLRNVBQoBZyjY/26pbgOa
ZB+bANNO7mGaf+ZvX9HE/FIcNoeS5/xYTc9wcE+Fdqh/8IercuLp/itrx54wUjhh
0QWV78XwM0O++KwXqhj1pBa/D2dvA7nVz3BH41jS8l6WtUC3QeCTflpzEhoVZjX+
wCGPE2qkiHnKTeYjrKXLck88iyOIcmb2MLROwGbUPdzUN0hUtzjNQvuybCcrakrK
z3M6n+cOkxoWPxVBPQ/ATx7evgK4tyvdf27vwugPUGRRyVRsG4OXEOKSBzE8ORuB
i9jzEMuNm3veA+1TUDBoy0p6sMy5Mp3KxdxmJiuOoAs3KBJiuZyAXppaNAgaQcDH
qOptOvyL98kyIfOpSDGDNfqpGTVsslGAMeq8NgIDTMq6AydnqZ3DrRulrMAVSq60
Z4sdC2altvOziLgQ3/PVgRvpkS0s/8UnMrlE2l1YMjPPpmjafBYjJVhdSbENt0+b
VpAXXBembOmvu7eQKGnxraz750ZxkhCLsqy31kORF3s1TUV3rwiKfPpQIWuyC80I
feQKDaOnLOftVZXKXAq2Sl5kOtSHrxhcLM82mLrMZDW/ufl+ttwtkRDlOBQ6ki9R
+Nwo7SBDAOJ8I6uEcS6qdrh9bvy2+G1u+OHlDuSTvTIgI4AQeOhKeWilOu/+7XuB
2BFN+XFDeJ4BWTuj2sCLsr1wb7oBaG99XJ0u3+dWrHZVlwI822DHHWdge03mg/Xb
NaLTlMVO7mqwgsoxpouhpfeMcnor0WpakuL4L671xWM0q4znsmsQttPK7PEbtGLE
ke+AZamN8T7nO1AbcBVxaGHdv+6URbTwX2X/xObRx/Xo5J9hHlWckBmWBLN7JMES
V11V/L8RHg91+Lu3ay5rxeAXGX/yi4/febeiUV6M5HNtpKWlv8OqSeffnD5VZWJT
FopeRhOIPrZrH74UhHkVedcfmDP8zG8ccSHM0CNSKW6KErtm5GvHGD2/0uhGOeq9
oQY28gXBiPDdexyoFfz7e94U+kNQMWGBSRL/zgsOkqbG5KmFew6v8kxzK/VpuDfm
PGW6EbwPqcShz7xO3+u3id13YtDnoIe5f1OleD/JtYlrZbkf1XDK5Z4OXMjNLInH
R7xrpLMVcMa03HOM94/3pu0esRcmnxiXW2oKTtiqHTIJTCAaPXIVlAP3ckqvHON2
12vzV6SEDRykFNvIhSgMO/583TZV5fgRy02ufHSwLumECVQbSRV8CsXQ5uOMtBuG
STLl3jAV4I9AuXJta/fvE4r7gaUB1GDwhjJU02d2Gf0evVMXjgYCcLvWY6mDVrI0
C9CuTSBWP8rP+/V9Ze11pBKZzwT9y5dKFEjF3wfbAUfXkPPUzGUjOwiai42fQZgM
lZt3sJRLFMcL2szqY5WUdpljFLB8gRcWFsMhh54oTuUUbkoz2AqX5EGS2IbTU0Zh
cfk02K6FNM19LW7T3v06EPOKqE+O1bmRBaGAN/9gya6VP/KGLKmwqdzjCdETIjru
mu9E7j7Flccu+UNU2r3V8aAJOuDXn265lvK/HKPDh6o9KFglrlPaKhM31jOZPDR9
syC5OWhijktHxZJSx6992OUmhLP27IumcvR9FJLLGJ+gwTZ+unA9MYy3MZZQ3EVL
8VvPTdRysHuxxB2G6oeJwlfpXCH6HE8eaLW4okPpLlWEvLGA1jMgECNZ47fH6gVT
6O8tzdbep9qKROzJpCBYk/4sNU66PfumFEHODiiBxwxo9gViJ931dms/lRQAQ6Sl
2WTj0km8kAoyMMikN/JxqX6orLxec9cTLQjByMv9ZQbEMeMuBplMLMHjha85NEhd
r5sCXu/TurRgGyPVj3cS5RPn9jb52Mx9qqhkmZP6cSWai7F5/U1fJC8HvVZ5ibF2
rh8WeAomEMf21Rnn9edd58qUO4hK+JkgSXjhVDYEJyamXUnCRqqr6ge64QHFski2
HKJ9mgSqNaTioogp4CkV0eFBFkH82ttewWHDXhgjPJlLC4KNHAxgshjM0Zxff+AU
5cnXaW9E0By/Iw6PEMqWiXyGsRqyRUDlWFsGSCYfnzRJxgIRSl9wCv6fpt6xvtis
qNED/pM0XoSqcfAjRxCaF1+49F6KbsjEh5XLHgBPYFSstvjJHBoFkqJqJwyJXZ4e
oSOTmbZqAgzraUB9VHdMAm5TbZqTLeFWwo0ePxf1dL6X+jQKOHwkuNx/zpQe/Ta5
1X9Lxxx6tdNxor9ryLWU5HKFk39RkJVX2unvLtmU67xUq5v40aLZuVG+mn4Txfur
/pOvnUhVhb185BVpFfzAjd/IxIvtxzKSWZ3Jje1CVgA9jcr4KLFS/hFpK/4K77Cq
0ymVwpr8ylugfkXZBXhEF61XZ59uUE4uoeROSgrTvn6avEJC5rduANXW9/RsOkhq
lSg+nfpRvhwT7VDfAHKPyjUP3nkTM+q+QwFyxSOYs07RccKLbcGUSJ5CVoWyW+y1
gBSiv8c4jXEpc8MrZFI4OBTFyEuvJi//gSANI4PtXQcOghPUFjoOgWtQhBAVOCub
tuZGaKLb43od/2dAiED9Hej+C3+O1LIBOq4YewVbOQ6NjzQ+khIKdi5eJiX0Seyt
mIJFoJ+pxSfHsRoCjuFREeb7/RfSlgOCCw60una8e6RlEx7uRpzOXd0hp+GT8SjA
PSTCf84TiM4eNnz+J+IRX+D7buZvv01nDJPFWvbUg6czb5/byygnms2oFz8DX8x2
gopRMUyW5fX+MDwa7PFZHgJZ937R6XVTCqlOPlqE3woW/Zazoh26V214Q8r4u4eg
6Owl9NTEPvev8YGSwlCs7vtoil2Ydz60IGX4Uv6KNSUTGhMrudLotdyGiBDDKOGs
bSEdYamvISqoubBFlFBFeUV0CClw6Pty7/3PqNEcUfya0VMy89EpqCHjFZOpPaBn
CFohpQoBFhtEyhZNmiHr/Bui6nrMydYZgvMuohOIFZUGNR1kFXyPlzGZ47DZ1CYV
WLgmZomawEWo+YR/Y2U6mxqI4OHKG57qXt/C95XrH8xC4V5m8ikdOo2Na/9lfBxC
HZBL7rnKJQ/pC1x2g5uEsTDeZw3yTfnQQFbuuO2tFI5hiqbogMoNL6/7dDLHZC5C
zppUSndbRS5UBR7dUHtH/eT3lefhCUNNlN2ianXav5lKKgHjJUd4U7fZgpEvx5Y3
Ko94rfz1PfRueJA8U7lMc6QOxgUQpl/196CfHgBgrB2wOu1Pc3CKF9P+OLXIcGkk
PC+OfU0Zyjy4nELY+43hPK/N2E5TII2aKHowUlPwrf0DytOH6zEVfwrmBmbfYvLE
C++2BFg07hXBoPLwwM2eCQJDUKkPJKvwD/nWDkm0zWG2ZJ/vJcQxnLPiOqyRsIQg
/otWDsWDhRDsqbqelvMB0ubU97zPANuLU7Ten2vm7P3jD3t8zU+GTAMdxEvZor7H
7xnwqL4Mma1NSNQgpmGP5cERQzOhmOrXZ47Ku4gQLscivah43B2CPEORZf1QwAv2
04pj77TIJe7ReyYnvZweOFEakLbJfEsQcbdPMBOGYeKS4GyTbH6oe4jUXycZjIox
mkQe+EZwCxV1GmBKB8+cAwu/h5cns8Hqxf+DXC5JryFflRJdEzQVXo/fvcb/DdPy
X9lbM6mbUcNti1Yz7F4BKXpB51o6Wrx4Jj0mAYJLN3GCarUhLkq243FONznVwkB9
9eGVkRBkjE8Svb+EUG6S7fdu2g6co5OdUBNo7ZtgAaE3SrJDKbqD1kL1AM/8dyqk
SzOXu8CViHZ+YjWydpnQjAfulDLc36rp8pZCNx1wmCUaui161DUzkll5ElwCK+yw
6mKLsCAVYUunQ4Gqw10qmfV8aVVrIOcvJfXKpnSrGfRvkGOxHwrZtgZ0+LZgzpAI
1DQlRm0QRRC03u7ofiy1omJaI1IgdnGejBAB+k9T40ECHdJaY8HiqgEbZeY43Vv4
xuTCAmjrQl//zc673Jw+XVdaAzyqxkCdFhRth6tKI4KJEeuz4qV5/isxlDNKMIUb
oW+A2eSyT9lP0kTYsZaXmfKHRUgkbB8sh63/CASLBuO7UBQKlysjUfxykOyGg6ER
2S6WHZGxDvVjl0HORwE0Z/GdhAFKi6fafnXRbvNQ7Ys4Zc2t2xE8S6u8KLx6C6wO
QDTldrbSf5JBqWV8jYfJNJDKbeobERs1W6mMqu5T/ApIdoRpCRggqFkQl20fHUNi
JZwfGx9dOErgQM6YnGKAIdrGhU3yEvxx1+Oyy2I4xaN1SM22zuQPGQB5QUo8jRBn
22pVCSPfs3BNuGDNAzaUNxavjpBJYoUJgYfINK0kih5eGINW+nE1yHur43wZGuRF
n3J5SYtg3mEPegi/3nFD78tCkTtpyCTe8ufbgg+XQbgsSiPXI9S/KN6/mvqgsOKf
GNFlBi0Pto/ieBjH4mkyEY/V2T3mFj70YxQuNU722/UjrgYYNDf5w03A952FQG0Q
IQely4YrCWk25O6BSvS/PtaR+mnw+5+vYtINlZcTr85YcW8nYPF6AmDfn61oz4SY
6GlYLQzDgvnVaguFpd1bQLIdufgrElbOBoau321Wxa5yv08EMOZlH+PHUXr7SZpF
AgHhf1YI4FeH//GaF1iNjQM1qyiv0KaJlvYwVlEP+/uwdOP/034rpzvKj9ujcfaM
dkoQw6g5A2zVTuWuRZAvKAG20BogIVY0ev2j5epPfW/1whpv8inSWRcnWKRweWKF
iGfQD1TW/AHhdTYN4XlYuL3BqShwcq7YTXHEfO15Xb5r0oUHqtrR8UsZtBUZPYVD
DOpziM7tUIApBYouw/YqSlC/p8QiLy1Wahqf3Zmmof7+eGn77k4XmOqVLO0PgDrL
+Wv0MVPEOfO1oI3H0vtPPpiX54UDYXgfuiKWrBI2sn4Ru/oPs/eEO7s1UAFWfx+P
Om5MGGoVrKkD42aqBGXuqg9Vn0nRqgA7djdFNtc0pEino4WJ2pkb5AIKwdTHqZRf
dXZYRMmErrhLTIqS33gg4hW7DoGhH2Ns4rp7Mj+vwHRR7IVVKd+0UCKeVoT0j2J0
921w/kg3lMb8faQ8VNf/V4SIaZygip71lO/F5Urze6WfnfL/5eGttOJH2ihBhbFJ
N4B31gxV0mvorsV7OTRGnTFEIt53RqvYLvpaGEMHfMmi7e0+10d+8IO8bJ4Wt4p5
kh9BDLmoCelpgHJNiZKzj5DVyfHxt009X2knJdotHNadIHRqcDszIcfZPH4KuoXx
i1EuW1OUsCRd+QcwFGczYuH70rQG1qA/tX0T1TezHWo6Ts+usw6AKcqO77KvHlGg
MZLTKguDYxdJWIxbIvwj5xEH74SHrbTidqIcmrGo11GXYEMq4e4ilYs2/mN1/Njm
S3rUGXDmOtOQ6zBhJsMsNWNUEk3Dql/owDJlu2xJrdxJ/gHq7f14clPRnbTDXe8v
6az4eedNN558oFQweSyKEc8gV3GrXrNRhQupnFW2soXs0yLJNc6bG6+auozKaM74
nhWuHhWY5sUdBeL2umdKh6ehiaWk1O9tt7qvPZHV/7aWpZmesYBn+K//HYbVb49R
CkIwGyoQOFCFlBsGpMZCoTp2zRW2wP5RHXjwxMnEUKS5KI1eSpt3cYh38+B7yYAb
Ouq51wfGS/c/FnozoWCl5KT0S8vz/PBaJXgSVj5DhO5Mq4dzFu5vjFNm0UfE806w
zIynuykIjgtM5XBtWXJHG0crmyyQgp3JZmG7jTzKnht4FQbI+inY2WXA70Q+PkVA
30oJPTWYyzamJugJXTVsvzpJ7P7wLf+j91m9X53Sur1wjKX0cI2+nzJZKMjEOVLF
HgPoz4AhlWOYyEjtjYuKDGM3FSwDoF8kyRLiU7hYBGEk/+llxb05RnG1kRXwuBXB
nFe2CvktqCTr2h9hXrNQJhqK8+xdSmOJHKwZmrmHEqq84gHK3eMhfnXNh2BC0oWx
`pragma protect end_protected
