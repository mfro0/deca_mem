// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 09:10:25 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mpHWwDptuZpRwQ/A1PBueyUZKg/a8ooAtJXJ0eSsCJwpOt6yeC6HPHw3jAS1cCpo
xgDiewbKBet+xmKC9+6Onc5wmXEU06gHASZBR4O/kNne35L+0I7FRE9R2RjSuVPV
aY/0E+eHWF3msTaLGWokT8OUe25ZcXxZcivI0qSsSDU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11184)
1ziFLh5/Zv1LPWMliYm6nwWXaxf1HjupEe88hKcisg42j1BGEzZnb4+bYStLmIYk
/1pnOtHOdDtWHY9ek5ctaa0M6E6/VwqFxlKsrcmclrPqpYgEH4eQyDJtUtVE/MrH
JIG4bFaaxlMl5SQ5Ap3A7Lo1XHeFOjW4YCfW1iiEXKXBF+8tPFMNzhbib8EOenZl
sSJaWcJV9k0ncr2UOY+fU0IeSyY2Y3rT2TJigW7Fr5UuA7UnGRBQoBTAFZBPvLvR
Hc0qXx/iytU9dJVPWfbwfBSr7thZAKVC07MDiksFjxOYsShY9H+QaNjf+BJtS9Zo
qCorPgQXrLh2oSQXe/5HT0ZFmBb5d74ggEMwEiDJW3pjJZlcwcJzTgYdLz/Twgrz
VLUTIOvuLYbnrqphZWAqafnxwbfrzcPqdrNawXemE98UT69pTe0nWeGqZRpA0kUM
vJVtLgosOSwPzltkPj15fsU421evOLaBhARk9fDC6bi7GH3H+mIA2/ppiOSQd9rm
NeHJDavK3m3UvqDhfcajAoppAwt5qDu+HPXqt+lUd5XAHEmohvctsORoPaR8KBZS
P2APkF7n9MhJPGVMdWy0pDIb4GjnQjBA68eYEp6JRSruKeQ/QIDXX0Z6wsZ7h7eV
qg7+lvw2jgkhWcXH+6H/aVvZSBWhG2oD0EOLH8Gzaw9lxs7UBh0ZBDK3c+mHi1y0
/u9qPiLJGw72X0p2/s2rCvwtKfCUCMHIGUVURQdCrXmmAd9n2VB/dnIKZ04W0/bi
DR4OyIumEgyQvkEeK6PxvJx/1rYOBoofXYEpUuPiKvG/VsFTlGT955+DY2R51nRz
pOxYFdmTIy3eitoGmdzxVkzOcK3EdfXrpQ6reBNKfHWfZlMsLUwFslE6ao0iozhz
9KpA+octzJKM1Hbikwiq6oWD4CBNRp+blnaLJZSTXbHHwdtJOOfn4lRKjKAPyoYs
b3VpSqL2GzZVuM+xH6NVVic0kelDUbjB8/4wpm9pox0+QNFi+I3sLxSIOSzgrAAa
fGWJfIj/k/+N98/GvwW7T/Yrj2A+xw8S57PUJ8lcDCphHy69CoRNvYAx8pmaYANM
Vh43mr4gMdAWRpMf77J8tcOsH8GtPRchTfz6LWeVLXggFiAOVYFTcsNleLpWgIYz
loXW+vLlkUvmhIANXDdE5FZx4VhBoGstgNYs/WEej+aYMkUYdSS5zBgbsxyS8u2I
kuY5CL9SKfAVln2dl5GvKn7VddFjrX6nrRnnGDOX5w1xrltv/L0Hkf9Z7lX5EzCv
84wnUgnlnm2ZlLYBQnNL0EJDhx3jlp1gRyHwcWQxu87BUaw/d0df7GNii1k2hu3b
84BXv4Ixq3SWYyTtRK3D533Sgats/YEo/d03R8HhXKLMDK/ue2mkjNDi8KA7DrNW
4WIrzD89suvb5YK6Hli5ENIiQSSS1rxRnE7hiZQdU4VrSsS6+07jMJvxY7aqJw72
b3F9M2LCaXjscDBIuyqozFLWdAW0cGvZwHkTQBvDbfML4Um8kN2IVpPku0toCoek
SEOtsl0M1Pb8kAWdCO1EUl2uJLGsvpAmT5y7zQldDwlahG4zt/GOMuLgKZlNyEPG
uGyKvMUspoSsR7PTKJnjUZY6WR5PoQCgYlTOxQYAWLdoXFBgEyhJ2IvPGg85yIHo
aT7NsSJ3r+cpfIvZg5vfzwHvLhfiYf15KjGT8Qi3vc2fM0p/oPcgne5BNuqzQtAp
afjzf8i/5dFW2213lw7cl1Q7u8BDEL3GPiFNUUw+YnTSHGJsS5T08BOgGoa0jHfu
gb0YyAN8ncmwGqrziVpIub812DH+wysPF7Mv4QK2tuJDtcYkzc4yxuqjQVsOIDwJ
bzQa2JBuKrNRbyjNMqpE3uFyOJpszHjZ9LaU3LCA3NpAzoIagjbMyvH6LXOBkE5x
F9ucKGahzX/BvU7We/wiG3XLhVZrm5TAxLsVrz2Rh/mvnRvKuzTF/1w2rT8mFf5I
s9VjorWpHHZVGYYTtPyGX3dTSlJxODi0dZS45LnGswv8J+BBlImrp33+IlNiTpCG
mgTK6LNwO53VepnA3CNZ41wKdBiQ9PPa7jYGan6pa1K5wqGpnn9XOitkBcDfqXTM
dZEMlalCh7OyBKFwDQwdveaKTX5Bs0aJQjk12AtI3CZUJvS/olJSXo9fpVfPJrfe
IeTuDow8WavJjPpI9ACUdm5zCbKOOnzuGrt6sy9SEReTJwAAc8ZqmhwOMJ2Neu6T
FH4njoh0qOiTQLPpl/ITXU5ss3VV9kGqJHSPEvTESBaCUFQ6hYvUo0HsVK+1PpFB
DMg0KKmaqfA7nRgQL9PDZ66j8inq1x66oAe2wjMYwW8I+7Zb794r91xAfzDCfu3b
BF3YdOADAet4pd1KradZqgt4F0oakuykLWfDgVJWegqonyDgGN1p+/dWvs3pO3RG
3PKaYPYZCDa79PD1dWhuyWu6tfr/GG5t/tY0p+IhxjxSjgCXEturUaZ9+ynrcjyK
nfcj7UQPwysH009BXiTkrjaFsRh6Sd5IlK6ETuQ4gQoT3n/sYqgHpDoVZpY1gdQr
hO6hpWm0y0bYUR+yH7KbNqk1aUVDOdvDlif25nDYO63S4Z6f6zy87ADNvuzqjnxr
JjBIEGx6uiBu/s7OgdIZ+y0HeQDMKUqiKzBxKGcYXOehfJ18cI/VAS4DPn+Qzwxw
xFNhH7/sor2jl5sfBI4eOj3f95zat0SSNmQPFs2cCxZe/Lrz/getFUA9/++conZt
1XTeNYYFhEn9Utr/vmocpfeAbVvSvRVcT0xK1e8z7gcDC+b0YVxjdmx2V6mqL7uR
k+sHryYVggnUwwBG6WrwYd/QNPdZUg2WzqoNKUVyq31FmO0VdQFLLOmraF6PZ9xW
3knC6H8HSa7+VGitBRr16LxQomNvhIUn//vsk0Yb/T0QbOnIeWH/TqEDcLbnzmh1
X7QtHwQo53ieXP10DBrjANzwhoXXLOTN2h5V73fi1Zx9JG4HQMNlTyUODqxdhORp
M41YSnGHxUmeRHS4a3r18Q1uLIC1yIkN+ZoriVjq5tAuuyuR+PmU0qS9IV6H2z86
eGJ8dObo6c1s8m/OfaeFybmi4NQigqALgsaHoBGAgbRyvSeJrSxJA7Epm+hRbLWV
UAqxGvAZ3w2exTnkBCSvtLpqtXFFCbuMspFVJtwldV8DWZM7LaPA3vys+B57KNuv
K2ktRS2qi6z9VPqZ/xEjnoawVa1Uc+9pSFV+WqeJr5jMocwNONZjykRSZ3H3mfIY
q0p9qD8F2VaYkjuxNJmv0Suf+vy/vTkvOxXfoHDwGao5wqzl3F9lUgdWsbj1FWg/
hXyy9ojmcV/KkEkTo7bEYI0w9SiiboDL1kadg7c1S2okdDP9xQL7jC1+8J5XULw1
QZEZ7krjFDv3JQBPQlq40Lj/ehHu2qpWbv20VbrCyCnQ1upBVYo5/wrIXatfT8rI
20GDguF/Sniq2uzpDJ7Gwa1nYSRTBzNZ0twVtXyIOHDA7evCVIafx/BRgQKsbvB9
POG8rO1ekUlg2fGbeK/sFw0QXd7+NLxFvjgxY9HK4oa3juN7Og8uFoifjV7mZ3mN
0os3BAbir85X+5bSaG8VHtiWTwMr4yJ/m6IUQXfpd1P8uqp3KDxkognhNCQVy+YX
kcDdqhHRFgLYT21XEaHFDuJ6ujhbX0LtqPNmZOB/xbb3glrfnisydL8JybmAjEve
uVcmWIKNTxuEAGbhqwsSeQwKATyY5sBhRGYnoKsoiwtTvn8ppu8+txltRrY36cPe
ApxFJCANWAWnir/GA3KHdNA70nz/W37I460j4lvaScQPUpeFdtLu2XE5K6+O7hVK
WZjrz4ATWRWHTCSlRKOc32MYFMJ5Yr7U9nEPlfEQ/X/+woQn+Be0zRg/0p5h4EUh
QznldWuhcpAMgwFb0hJWd5PCIfgQGr+8dhlQIFFVvm28WI0CYQuNdi0w8Sq/e5Ji
DPKvcqRfVoi9bF9pMHKGGAVG9/+Uf22+8k0IbwmVIRxhbSrJmgiIrB4yWaHWRsKM
PHj8ogVKjka8LXT+B+wQnTzCrNCVl8KGBbUBqAjk+p7BTe1eFFf87FputxxJSqSe
2DqVti4PqRd5Gc8bl4WXRguZy4CiU0rqRZjLGqDSZlMgwoEM1p/6rb0Ej8Bsv9Rc
c7jFBAD/sl13Nfyew1+NlJ3rmpd1AQ1tyw+aGp78L1sCJlVex7If6DFDv2ZmzY6h
MO8wzN99pjCdV+V42ptyuxJq+otydDeAurz7mduwlfPw7JXq8gqhtdsK8BAt+tAL
G/gYl7drzE1qZrlU5RH0E648YU7WGgRTGVAh4MyYA3eKtIAorXF8DL0E6djktMsd
1CcVEUHhEm344oFOrwQzTmhN8VJxajoFJezxaMEu91f2Mk73P4gY/zVmsn6Rv7cE
3IqSR1t3D4JEkC20nUKelcVw1PJ2w3I4RuiPxFUNOtABQiTi73vY6a3mOBko4xmo
8gRf7e4UFOZEflsaw5s+Xpa8JsCecBfDEHdzfvKyc88lQF6uweQZ40lZ6eFud3nk
d95f2B75FGxzqaCK60Cq3fzhUzXpA388lYvAk6WPszVuw3BoWYCIfa41vwgYEg0I
b9xKUrYxKaBUmr/GGOggGtXx2/Bdya8Sh4lO/dn3LeshmLzxhuDFBXWsmgvtdZKw
KwKJy1V5iFH1GfBmZ66b51Y1u/u9zAnXWVT60m92eaMFTs7sp4BqTwrdDGxawesC
3AsJuDC8H77i/9uanZo2ai4zB1H+iZ5BZFVw8C6zb+2ncGhLyedfoIvbOhtoUW5p
tgSsVigSuwDw0jyQ+zPgPHPvheC6j9WPZtdxr1SL7Oe0TBY28pSFM18rFrsHmbGG
kYGZr4M7e5/mJMmg0zoBQjsEnH/xCpZj5MUAaBF3yml+cOHcLl0xacvUQTB3teiy
BWYGZCvW7NHKdcVTC1Ss+aC+qKOwrmt/uUsOgHITaYFvNvCH50dROWY/7Mr+zotL
9ursOM8jrkCcZwicGtU7LesoFJfPOWWdBmq9zBrVo8ifsCfi/PH98/+/nt+++/XP
tU4rBTaGn2cLZ7s+LcXGW/wgvE8bk10W9lrAgdVpS+gRi7Dm9i7ovedGXYLcz1z/
mtRa9IL36Y6+esBcZYvLNOVOnuC/XFlH5DSX2+mX/xg/T5mOJKmN8nDXtrjaj/DT
uYbVrm+7qyaXJvE6N3kn0A85Eft/u4emv+M7LsGtoNOCAFcfppK2nJ7eHai5YbiG
48DD2lh+UrDJMJ+TWMX3MOcUqqaHViAZeViGu4MOqR+rggq20IWAlRDOFDBoFIwG
hQlT/sM1s+WEyo47vnTb22XoSZLHW3vCLy9R1jjCt3fOJEsKv2sNh+Ab/q3RSSYi
ebhx39Fd+BUCyZC/I52Sinskv6u+l7ggNd3YUrf2TU4cRV95zpfy7muNHiY2Z5DY
xa01eHePoMT69dxRfHK+58NH+3oQKMMYv88228J1RCNbywi9ggN1G75XOGZ5OaJQ
wAVMVQ3cQQk9Z++pOu7Y/fkE3w/a3h0DzwkT39yyaj1wXc04Ye9nbKizcfM0VCr5
x+NNjtOdx65IeqpGo5VTe2exTiaVONd/GhLMDrWQ/8XoAvx9jClNd4UeghmpABMO
Ek+zP59UQWyM818pcZqMhiGr+kndJ8HUTdqdsFTWBARGKvpq001cjaA0xx2ERwuu
hV186odEaFneahilNmQSjTLg8SDrbh9id2qNneaxwhOVZkzcURdhFlTzLTAOFIiB
mM5Bu2LxXrEwyIGFeQkDv2jm/2kKXwAed5w6+iBWrazRC0fl9+YgqqK7yNAcPF5b
dT/QJJxOhKzrYw098UJVFIccD125f0soS+KmIgVUWZWr6Hkz9CXNtcOFwvz63te9
+j47trs8BRLQmZRfCKAe9Wphfdj4cvqUqqjHpbVyKqAFeDnPDzD9wv6FOgpqgE1N
bivoRZDI7MetiYWpb4Ra4WJSJS5g/a33R5Sj1H4pD9DfJDbz4B/IzaGBtwdloEDL
7HpDTFnv/g24xbYEjucx85j3972E9pJPCRL+bbvfLAnkF/VXM77qyERiXz3VID4z
wfHFlqneoOZUfHrVVm9STOkkO/35divruCtIi63UjA1sNc+hgEmqwzxuCzvfikXX
byiTngpeNQVH/4i0CrX+b89rNgr1TLugejX0SyjyxZb0IFa3pDjQ+WcDraLKWTOc
msXmEzgYBe1eDERHn1rj+CItDy+LhmhlalxughxQPXoCs2NjUFoGbylHIsQA+8u7
c8CJQUcEQIhNOfGe/b+aaJ87eTIxYjeStDYs6e6MIvjF7xEfmCk1Tl8hARn+jAl0
HLy7m69VulMoUs0KwlxgHJsdFiqk8bSNRMb0BBGmc1UNjwcHiuD8QNNk0BZDJ7P4
05vOuN6fznkXIUmxQPLUR7Dvv5yUJVdEu0GEI81Ob89m6kLb6oJ11lfI88lD3SxJ
enGzal2JbnLh0KgRtOY3tB2j5IVBfUlnrIVHTd79eOGd5mJ9XxSFO9h6dSfwIXVe
Se2Ri4tvLgyOhEklx3Hf2KQLjhp0EPpylX1IMdljdYf0YzVuwJrbhxratEuH7a6A
SBS7kLBOLojyLVWusQA7tZcJ8QwjsSjvDKwiWw9BXYNWd+hKEf8yYMfhrlIHh7A3
VIpF+6FytcpZKbsgkj5yQ9/qbYlAbKNwsA6Sem05X1a56BfX+qITB8608lX5bUjc
erbYwZHinK3PugLU74rIbomolBeXJSzFyGqM+TTYmvtFaoAna6Utkajc59gaRyAO
VHckSVRLUfXo2uDiqO/DFjXFY+LRmL5TlZcjmzbEhjLM7qdfsL/NUqsOhdqD997/
9UrwclfhFUkW75YL9YHhJ61EsLTbHoUWHPOBJ+JGF4Ul/EYpRU9ZoK4NnTePH4Tu
FxMX2XV1wEed712hUlHxJxftx6aLdDJI5kIMZ9sAYrr+E6g0S1q6sVYEjFQaSkmc
ENIw021DX+wWiR0YTxh27ELTmf029WG2/cpThy/QemnAnABHIX6Vr4nWiHvYJWrR
A/1kKD+2WwhQfq+G5IuETT5XPuYjSr33YGj9Znkv5NM9uQhArPQn1wBPsxuGG/EC
Un60Hsy8eEjHuekWUMJ8F83hiyadaOR7YH7S6ScHeZzTPeGo+dBAvlbG1aXxhVBU
cwT1zWDp8szl4jZ25ArN+wkeYxXCGZqoZu40ISPoTSYUtJv6a967lfxxraQiZJIL
qVEmIYr0yiqVAOup0vX5r803m72n7Di7hEjkvD9ayOuEpzaBYcS5jboGDSAmQP9G
36hCE58TOw7jrZzhwzS3qKwq/dGBNNvd9eBvXA86pxncI+dbOJ9dh9epQyNI4vU2
LkBRwGL1csp3Ob5FEqRf6LRKbTcgtluSgt510IJJQjvZvsvim5Ju5LspZ/tUvQiX
bN4WKNw9//FgUYRDrA1JvmzMOuUW5ZUbqcxhaZE/fTAdFlMytDI1l9gvCqrRx1TL
ofmnrvjIOwmGBL4EwxtBRjlYBVCxP+VzKocmeeDjNdeM0EXm63n8mQBttyGnhrBU
Mv9oWGovIREQI8kMnXYmkqY6x03LLQwp5yBL86iXrtqdUTrADMtGxK594Jkaz9Js
BiUvvfp2DZXlBqygSTYm8Pzsc2JShb8MBFmCGf+glzPRQ7BWX4RrWC/2Wszz4f0W
Je8ikxnoTLmCoyjUcvqQmU6hzHxJdd4m8mu0HmwaZrIheceqXTYFJQwrszjDkZVE
mvZIKfT3cTsQLUJLstJF+TI6+We7qvo+J8mj3VF/khO/UEH7/8ST5Nm2GJsLlin1
qh+sG+z+PFCMjvZArzujW2ctsRY5LduS/3xp9U8rSqK74N2yN9VsrvjYqU29jJqT
2JLPwFjwHB8+/TK8MjkxMcFqlRbX/wLosv6MoXNsAeLgg3XUAqt6qoxDQYGRmdzw
njH0ozOmnUN7bTPvPvQcIS5jplcejdh93W3MWpbo48rL09rPiKqevJsMAWnLn9o5
KTR0T1ZTuejyV16qmd/yW8IryWceL/QXxCwrsE0wE53IlpJpkDKgFZWqQkwuqmsX
0mTrkuc5qNmtcs0Yyx9mkHbm9jksxpaqzW2jQOfM7iwooRy97b3T00cUjOQvWsi3
q2UEkaY9akMPNjOxCtyTz14MmgWhbv0gigDRD6AA5e5eeSbmUiicVfee+GSZxC5F
EopF8vKAkmEVYumhHoCCy+Wa0IiVWfL3SStt5BQictEK8CAGhLnZezsHCQuUIGR/
+FO1HnaHuTMuG6ef8nmgGRN14+LeC5ZeguSp7PWVjXzD1wKxNhl3pwDd+cYzqhoq
k9JtRVG0egR2KBE9jGw84cazt4nL3lV063WBSgIivAmkpM1WziFxt8X+Leywe+7/
K4/dVCQYISqY/mtWjeteCHoJpSzC46F3fhmKH8N/rdeWfZ1y2vzTlk+lckNgcFHj
Szf3rRgLZVqFxTfLL6t/8cJT6irkH/fLBrBg9GF+Vd7RLERT/whS5jlqRsbn3pKS
onKV6duci8Y18aLCBzgk8ZXPiFoZbPSLSVUS6fpIYvvWXmwzfOH+gIYGp1b6c+uj
PXJa7aFTGpWlnfRDGjdsdnE4DS9hlnlM4uVtFgdMvinv9pOotXGbTGweG2QqMaKA
2KmaglUSxZB7fTu4kHUEj9ypBrhx/HhU8q3yftosgnYJy1wlWzpXhvdRiHNEM4nf
DFndvB0UjdyNwlyM1OMDqcVNOZDsLGFqNjTEDgEAaGcVImcMEbjVsdLrB4bvv+MI
d44gq3g5srIX2YhGGWeR5bfMJez5zVeeft9kvK3o5gdrnRQ/O2e+jLDduc2ATYAS
mDxNAfw/bY+Hx+QARfJbKfXL72W34Tub2L9U7wFKBXnulc/MBwmSFzsxfXbtD1SJ
xSuAecFUm+Bhz25Uve0TEzSaWKRHgCfj6l9lL8jZtzJrWyIhz9GLwsSwyII1hIk4
YUlyu1+7sv3VammQhryZFE16MhWMD0F4LLTwGaejGhgjSJBUBz2A9jzQS2exjpR9
7BkhXrqB9CHJ3CKgJCPD3W6IuvD9Q940KQIv8hzyY+Z1rEottCgbc1dzKvxkXhK8
Enw+LbrZHCo/CuxTC6uavn32lRcRMuvpzSyHWwNx7jqbXjhyt5nQ7yPouM0YQzve
TIBLDXyN/Yu/Zveobj8SDgX0WnLkmYaMAIXxjNMz+ywm9CTi4XGBQHUatzTr7xgJ
flpFnzwVagCOIXovvOmYZUFZjoUGE3JuLWxSQXAxHQn41bOh5enkwLQvC2fPvlQv
mspCemCc/5nYwl6vjHCdgPI18fpm2FPkDpEt0CT249QiUNiQg/AVNwmgSJX3qNf/
wdKi1jOA941FMhF6xyi1GrjQB47XEIImHxYdAjaC8MALZ/WDj/uGbv3cmPiDgsEF
L5S81hS+myEYdgBnT5vcKuXKxpE7goAp216LJvSTK08IMhhiDK+hYQSpUXkptvW/
4CuMhYbcKU54U0HhhV29mA0gjGcgFqLjpgbvJILw8Om+q7kS12ejsHXyjpRGYH66
ewF9wosJlS7OyXODYUhL89+jde+T5CVbnQPG3yZ5OX3f46jNntljzbwFLvPys4Aj
WHKbTp8mBKLlEYuDTC9lB6aqI1zeCGzp+UXoxhVLsXj9/pDtLDvtZJOF42iac0dD
JAyWF1UINXcJf5xIs3OZDPhEjv6yIPIZGDwcDTGFUPkdsIOs2NXEYT+iiIKnk6yV
jLQKAqcp5bzp7eFlxiAzaz14eTwqMGHACi2eojTal/PcuEDFA3oE3/Y1tWQ0DBJN
8GrvX9xbP2dCwQVZfv+BFzm7wChOxMyKGq4zXMLC1J9V8kunDUab7Ld0YQsPao/w
CkjyXo1FkxIbzdDxHHOT4WrvlYYqPiFE8eERGZ0B0cjsnR3Dag01JLS54wtNKuk/
wgJGKMJ4abvvcHAsz9QKUhFbFe/75x4lQS6HDiQUa8UUJ21c8iEqDEG3OaZsltTr
HSwvjixcAvT5O/M/nTqZCiOLD4kn/QnUBxuzaLXytKftKPXsjEr1V7DcwDapre/C
nsqRT5AK0dcizyfqiex6g1lHPTYl1KfGE/d6BbVHsdl5uw2nw4Nn3nR3r1O93yIe
+6pWhLNMevcpWxhBe/cDDjiz6USmNe2bP95uhAIy0FyIHjk+rSr4uq9rJMwnielE
wxm4blRcG3SXSDv/xpzWDINFE/JvnE0NLSoh5TP2iqOQ+5A/MzLH9Ws5Zy4p02bz
Ga0112aChS5tZK+12sFOGiuWqAbXOqhjagAAZEguKfYhQ90sYlbjSv5Way+mFm56
DISGPMStLIpIBW74dfD9jc8BSJ7K90CdvMieyTZNOGNqpugkd/VVkH1UKyIKbFlg
HFXf1eh7yCa3A+1UB2N4OYWpwG4/ySjyBSe9sioIbxjFodQdnk/vGoTQ9mFwUC2D
3BvId4CILH2fdcNN5wKzLF/ZCQp54mM2nJgBW9cbXEKDcBW24Xm3KREVHpzr/soj
R2p+Lha5Ti79VQjmWgDua0mvgr+NMfoKcqBvwZgKcAt3nsiy4tn8arovEELvvuGX
n3mRMYpFSPoeatfjpqOztpGNLIkZ4Me2qu2laI9Ddoek+TIXmEMgCn9anQvV8YoF
5LyxWruzKfmrUnDZg5fKySE9q7wiH8bcREdze4nVpytdontJie0hMSwJnzdIStU3
rQgSU5LFH8nBAtaekucfz2p7Qtm3O+IFgBWBcJbF8/pW6nX2dmVPqvT2vYw70BTz
a7YI8DMX4JTmT3ILNIwVREY2hwnWZAkoa+uo6l75wzqBtqrA5QApwQhGerzCTf40
6fj6c2uqXDCpxFTjkfY240da38KfMCgLOJslJSS47TZDI0IHBdj9KHAWE3bSm8A1
QilkeOF4Pfl4t+lT1jOyPSuTRC48lnCWRQ8jmTYSRLB4xmVNaGewOW8GiHNT8kHc
6/0Lyegfi60D2aLWsIwW/EFcCdfKAC8E3bbT86KeAZzJXLzJ2ycsTd/Tf1Ikf7N4
1VZhCnBNmMxR9WJsNOUZ9xtvbpuVfZJXdmiQMUJK/5onwr39Hz3c8BezKV+8Hqsl
B8HaDJFaQs0phYQEAc/tO0bGLKbUhi7zY96FvsCKfRIrDIo52rf41r8QiBAe9iFE
AsP6aVD6vAI2cTWOwB3ZLhM7aaO56NITOSSNvb7focG0R9ZQhZxZSuPrEoy8l/LG
j7vF8HwhDmzTYGaalXvYq7AR+IzH3qSI9g1fPdrsuCiXZuXvDth3T1FUw31YHwNA
jq/XfQIW0Kw7SRII0XW2DenNoU46H2yTdnZuTNxg+Aa0TlEOmwsWOW5YFwb8Qfzn
yn9QQQnYDxZ7WI23EFn3tSWl6hFzWvKjnrShCRmd+PLCFL7cZPWMRQmdky5m/DEC
8yV/OvxOJESRPV3UUVvSm7ShzvUGWFDN+sNRC1GdO1HKuf0VL4AnoUKAMIVnjoCn
buScLsN9l0qhRBI+PLiv/rZBSP2OBH3psnUfYxcDwduc4XoywP2Kk/m8TNLqwRMq
wLyiGY/0DzDfGfkW65DCVG5SmT4KtQiniKYoSHCNgX0pCmOcy/k+19L7blrqBaHm
RnlhWABzhDIjy5ut0TNbeac777WWhrD4qjenZT5WLbtnmVKz6RZhVQ2mho6yk/1E
2OtY3XdtoENggfayevt9tNTJs0OnO1JlFQslg3F0aJXNaGksZ9JaFc69LNUrDKgM
/JiTigdcKmA2pwbOV41nMx/Fmm9Ux12SZwyxipaKo+7nev9V1+k50rNuL6mu6Jmg
3d2X9GKht+1qtpYTxnFcK7DEkA5YuftRKCQ7xxMom9x/GLHsONRJqCkuv8/Nw01J
aX231wfWHxDaP8eojCymyGLkj/LhHQ9P8DV0eQHTvOUbuow8QEFA4ASCMo7Ji59q
xnxoGeyJDN0ObfZ0JvcncYR9IPykOpgwjgHhg9pDG9yheCYHPaR4g1nwqY91FNM2
dazUeJOYD747v7gk7nqWZ+qqjjkKcrBEs6ZClGxQIX1GtFIJZZxo57b6Y5hqRTgg
wbZQjuF0pxasko97M1Z2qsWIU2uMFM9RtGFTS1I0eDynM7QjpNh6GyzMB27P4iMP
4NNcMSE5N/bu2En+HVgTGIIQIBnr2+YVBJCHX/iuXtNmHt6qP+m6y7YsLVeTVjf/
REr9pt2fMzwARCbS48S73yx47AenSvvBsBdb/q0YlzKVkusOqk2X3G3GeIPsMH6f
u00DO8wVKGyCJriCvh0GhrMfzUpBQMuWPYNLC2qHNVI5fY0qBEwUDmakdpazdjDo
TbWvfcUrynBCBeiAjZy3ur8FIVTvnEnqv618R9ZMRVLS0KbK2YwtbuneFKspahDI
YmDxLrhD+9ZNZGmRIiIhS1jxaBZJ0GGppiJL0o75DM6T2n7hPfpp2dHVBk+fF2hv
gC3nKUZuMrF6CEtVrgStsRRCdZQ6zjaPwmhQIHPCbgups6/sWAeAj5r5SC+2WHmX
AfHkTWn/Csxlnq2oKL3c5M6qhAvclJrQeLTLPwNhhoZ38Q29jjw8ZEmm+npQ0n6D
Li2Zli2iOJY6yv7pRiwjyIkgixH2xDX3+PjlBfc4hZ0c4zYZw6/qzFejjHtkECnx
to2OR2mmlRa+fgjPkJcSn1OmGamsVNrf9bvDjoFBV/eLOq04EswTfhwhWHMyZsM8
9jat0AEae22zUu7ejGrjLcl6RGglXoUEZjRUvfmRjTNo6rlktKgRpWA/E/A3ZjaL
/m5umTYeVLvZtpygLdYgIr0GgwjsdcIZNH7dr8TRR1XZmWk/yGL4cuwcHkuQj7/t
P+KfcivSW5416/Ux5vrxZhrQGeuJmALTjzBUUfi4M3ptHA+0fMyej0U9uN6isvnR
pYM5JuQrQ+54iBgYhYW2Nn3B152/HHbTLuRimW6hLxkBq3y7YuxtiFqyVpURWSLl
smcBMVOkUrFgEz0Xr5mjkv8OHxwxVQH3vltUxoqUtD5ATmO6ax4ENy2kEQSmsvpQ
KHJgP+uQdchZmZa1/gQkCV3LKdQuh2tl8Gv1UpK6THFvphPZfAZxiygZRjhLoQw+
mY5/l0N6f1AakaFC7GDIYbxNdW8qAz3TkcL+7IuDJwRqAY1tHTQkOgofDwykkuXL
cY0cIDhoGyJhYzAwUgC8dZ0ynjEM7qInvhCFfPLJzSv6MDloT6yU0LLoDEbTEfvd
YnRAyK0sWmMDS4qUhRTX7wCu1672cFG/Afrb6ljypMGnNeu9uo1usYnqyNM4cAaN
0iSoRdn+rIta8UEwAdtO9uQGWuXt8zUgjbYDgdkT8Kf3E/O7HGAQM4Eu3+HWEf7S
RwW5izVfpMvkqc0LdaNPDfC4ooD9pkTRpo56HtJJOcwByFREIdKrS+3A2y7fdkJZ
MOAoup0vjJQGe29Ngwklha3vxFLfXxXkjRqBhMmyq1DSjGMYY/wufcDlkAq9HqOu
OlRfp05DLqLi/rPWr0pJjPwdmKO+2gWTPANejOo0aL2krbgeQN1vLciAUHjX4EFO
Bes/adLo1DGR5AeJIDXyDZrj0IiJ8wW85czNvnJe61PpnzLBkI8DdOKJwFuyeNei
gS1K5y4pu+yEEnXJ7bdjpaoOKmEnf/Okb6uVR0RQMslIv49KFLGWTLHlqAcK+Iy2
H1xNnYEMuBHxZVw1rANZJkwHgoRTD0D3y8FeLHi9gVEHtlJlKtkKc5K+wLbJzZfT
Cj9fpn8fejg8Pps9m6hOtMoDDfkzbEUuFReLxg1ACuiyWT09e0S2IeipT4qkV1WV
caq8EYqRLRuumrEd9bfIl4q5Xfe+quyWewqanyHRDNvT4VSsW4RVwrqUmEx6k9x9
nRzpI/qCb0ZgGYJyqHVxYgK89nn0z94mpgrAmrRnrTpjHlacnq0WZ9WIhvw0uhbn
/FAPyeR3qMq+6eTaHPXscbryftGYDIRbvWeNY7DyorQJKSZ2YMHMnirHkRf/X6Bc
GQabRc9xAYklR10qFqvPHien1Wfv3xv0QhFws4Ci2jLOox+/oF57bA8iAkubFP9C
8cmk0x7xa/3q6V9bhqy7fe87jaNwOv4SXXvq1iBWRyBcNYOKQSAZEIIs22aWzNuA
GxNKwES1BBbOYqKU2sHWuzIzg6iGtVxsaWH+cX/hCGx3ShMO9SDIJ9/91lI1x4ZY
fXyPlanIwZEyakyJdTpwyi9zkeyL58EXf4svgpNASBPokzFiNKklkRojQ37hEA/b
Uu7BThEMk2GQDEibbxZjh3TXm/EI3/QObXyE0zR+YV1MZRpprqHNFyMtw9ugDVgV
3yEUZMC0tVvLkLW34m2A7GAOMk4iCYnX2HOmeZ+1UUjO9HaeyvMk7Ro6IdCsliqI
xp6nn9ozoqxoC5kUWl4IKfvwGif0cUDPEAhhncLFKS5+yoL8COpr5icM61V1EB6M
8oSEZlj9FkJVEMqFIYnpJ0bgz1X+357w/T+FNlwwo4Dilqixi0SuSMdi6GOrwI/3
cp415SfYRRCoz229KDn85tzHG/lW+qpNAXaiFtLCm8gUAxxKAk1m7H6rcL1B921E
4EQGTp7IVvBcBbUoM+qZtdxGmzXHN0pRYA15SFGV5YDiz4TXczaMyNAbkouUOCoq
0MDp4ekSJAhyi/8M74U6l9JhBuI8ssAXEmfo0vA5B/MzzsTsbtXXTE28Y6QfTuXD
LEgEkgCv5Rj5L04azja7mRClj4GzA7YAW98k1HEv6rxNywi2zJCYhcPlubFga2M3
e7XqbYhLTuHo29npZqSyo2c4ZoCm7kZ8fvyAMOs6x4LfkIvW6AD8vhGGxSwhh86q
kemY3yDO41B4QdzKoQtzbv+wA5wR1ppNpss3RVtVP+vzbjDTZBgRBmFDLKVeC7qK
vGWN/+NKcJJ2HPQEzEc0qKkNCBjfdghs1nNJeHcowvA94JjrS5dR+vEK+lkGpc9n
`pragma protect end_protected
