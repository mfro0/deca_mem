// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:50 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OTzCl/H6MSNh0LSTjrcVIU93H+2Q2hireOjFLWmdshovXv4BkkaM+jfOlF+PYNbW
Nl9iZDu7lrt1DC1qqEk1e11Kux/a3XAlqKS0hb5IacchSc/JhNLxDtoYhLcwwk+8
8Evsd/CwNvSZeym7yRc7I8lV5nRsElXvTq0gxxjEfdw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57904)
wr4ikYhLC4v51C7QAhW0payM1P5AKrGsaDHGouj9Gcb13/1o9MRqj4OAAqGZv853
w4/AExb4hgtGW8NKlZbVdeJaTCzRCzUyw4yIEKlCQMag9kylylGP3OVufvFOFWdg
CaIfjcO+WZ5JxObl950ef3Vts04G+vjVLjhX9rOMGT63XcsurXeRMZASENA46FvM
h5V3twTNAMoSDEFPBa/x0COTQ2YjRJb40/JWdkeF+5tLokjURIex5jOIXN6Q2ACT
Mt6CVm2v5bBgmGyotzBIqGzZlKY4UyUhAw+vy/iEoBhYlGlDsfmBAey3s6AtCm4h
+kCd2886Bj1CWSmTHldZkq0A9SyJ04y+Qz2tFry5ZcA/Gunc2QCO5xtJR5yCv+im
7GGkrtd/liyEBQBm8P3rCHeco4FiQoMHkQ/DWJB2WpWoYH7VJKf8RKNjyTyfrNlB
Yj9yyz7QrYxj+KMA3SKuiBzveOMQt9ykdmNDQYHq8dPiFl6gXPR3Ztdgr/a3EgxV
m2olMGG5nJ5HlDxUhsBECpmXpVszqTJ1Vu4U/Vg8S29gijkWowcggdZ/W5K23AL0
9tmhRGhOoUW61Cii52voumn15JcbmRKz30iBZAqLzwBbFDQMARo/E9GTJpa/uV+d
Ls4M/xuTMgbhDHx1Snn1gfjrtKTq5rcuXUHjIqvh3Tziwc/3TkpTG8RyEkgQ2oOc
zNwz3wtcDVc0YwJt7rve9kcaxi4CZ0l7zZ6mHcCNuGzH6PVNT2pTz72xrpoXcgKy
CjVjn+/H+aD7PwFGh0uw9ZL07gBAsfsH43D97akU+yJA6rTcO+xPHuaR8KrysWBA
OBtlTfr34hDZWwCMmt2L1zKDl9KIH4Nr4k+sv6HnAAL4I0b+ApucPVpCWiHmsWdx
b0DTlHmXI0e8StjuWzBO8TNVfFB2C2FTRDBsRSFmh7SoxJVymuW2nHSOIaMKuC30
N/JRBkV4ajT8hpYalZj+Dlkcesn+sTPIdV00uoV9QBcyjXvpDXIYnXWPODn6++44
mLL3lkJ/sETzEeojQj57Ot0f7/L4N5zuqpAG1rHaOKPGo9ZuiIthJupoZuiR8bKt
ySvHUHTcUQbPbwWuluQbzhPm8CxzDNFNtPNeRZlpjzBiT5/STvajObQEi0Y0p1Xh
t01xL7sXTyO8sE9GiHtJaDrNXrAABB0xgGX3dfj8mNcLSrQKmP3YsGXoF+u3KfbB
vHh5v0iuDLBKn7YIBpyzybJ9i2Z0fl1pYEwbahUjUgaTObPkBhhCeeYqkCDVAweY
xM1B7sR53DlK+402vw8X8lBuWj+UZ7Ia+HRTk+mvQWDsn1AeyTLfKXUAr2zmyxdI
8oAVGce4ztES3lvMPihhqVmq1XL7AgFXDhubBzndXtfkte2O+26tRt1tyRvs74UX
/xlPwsr5HOOTs0ezRvyESM35JGK9RwYNSN1NhVZ8Li55jzyA0iRLGn1W7HNk4gpM
vK44VBqZgasMKgTA5BfNO0VCQ1KbFe1FWeH3kUIES5jU/N+tITzkr1HewhmCb1nh
BG239GNLm3AfvxGe6amjkdoi9zorGKo/DGE1glxNByD4iCp82B+ISWF2MPNEDNYU
MLJxd287ThaDmTEOlr2/Q17qzmA+fpVX3iXzukYy9jQihzssC7hrowJ/9hbhxyKc
l/q/WQ1oHSjNNtZnwpgVnyBTlo7JNjRJoYhbWrJzXim0rAoNdsmmTiAoqEwOmnVU
o9NlHaVzlY6EvPBk0IPfms7ItK/gZ9BdCy1oVwU9MHYfXcAFzkgbtOwbBG1/KpOE
MsGIKqlyYCO8lI0j5BWfz6A14k8euWyykGVQs9qbASRpGJpttWq5gnT92Wu0Sh6Y
ZUaZLHAlbUjtd1jFHIWOYLRx9UQ6bXgCQEGP9+2NFJdHqoeHuH9k35N2Ae8BWdEI
SYH26S/Tz/V+vxGaE0moOWQmsYQSaD8QZJIMq7Qjw4JCCZLIWGGIY2bo+nuhOIfq
te42BLIX0bEB8hIthGZMxn3K3a31OlLOYbdqbhDBzqiBtgiXO/Hda8Z1vXmrLtzl
VAxiJuWXNE7WI9kgy6vWAN9lLHaG/q5IsyaFf9dw90lA0pnh0h/Ki55aiZuJo8MT
6GEC36+y+Yn0e6hDjbt+LGftXksNJDwhBEAId+LldXBc+KJTIh/3YI4gSf4lH+TD
cZzhqQyUlq15FrXOEmnunZ+VKkM5SFtasrUvcq2h4VEw7qoM/8a0X8u9yHLeOmCa
GX92ADyrmpFitj7Q0VheB/Dqx+QmEIK+YDdYlcu+XuwJUhynFOyAAwqNEoSFfFhm
8+ooO5ei7nO9fE1TDJrWSkI7fOBQ7ImhOkU83GpnB0dOrVq/Q7X+R0Sq+ucFyVEz
ZMhlciF3b6lboUqvjqZB46aFuXiCtWM76MAd2ykiYI02pMM5bt0c0eDHcVwPIFIZ
1dF6WfIPPfY9SgIeWEF2o74ZtBEx/dy9y6l6ZWuhSsXfB7LPWD7Urn6qZON6nY1R
8/t6ytAEgYo7TcsSxhfiPc6X/35/0+d63UItu+aXAuw6U9jPxcL84QV8Vu2GEJRT
+clQkOhXsC2A+Sy3M1FeJrG8LlymBiFBCI3I65EeM0Yy1LcGhS7377GsaZbroZPj
QooAe2mDRi0lETi4wgWYDDdt6u32CdiquHdey9naVHwzb0v+YJfYIZKATRNlQ9I+
1IJbfNmSZBHuzwwxa6nDsyj0TW+lk52OBrxl3BaU33dwfJ6v1YkwJaA6KFGWuv+y
lahHGWxFGupEkTEnBN/3oHcP/HXwpYpLiRGCC+aZDyqaAC0KbnfwzuN2gREHHUCP
sfauqayYsK3TTZev4SQqxfBDSMlSyA7bQ5q4FUj54WY890Wsqs9ElbZhLPNteKqU
ECq6pbOVTm41PknidKOwdx+YSQRbWvvxIWUvfr4kKGqEJs43Gg/pAoDiRcUiUq3o
7qILd4J55VVzulNOyTOuk5DFLbCjRHq919X/Kz+b6tlmSTfsRTy3Ez6/hsDtBFtf
onEzxsm2o/a3/Kkrob24WjImYAd6OEVkf8lrM4+t+Q5vj/N+DdLhTgYJVMtRotqt
s0+31+o5PDGuQ//8WGqO/LhNsHAI5KaG6bu8WIV6fRpAR6gjI0GLlpNcRRAuGa7t
KsB4zHmEiIwCtjEZEuP1UStLx/6CWjVLfict0Oa92rozh/ngy0as2HDMk6+X2/Hw
KpneOUDqdaxFjkWsBPYCxWP406fzn3+6NzEH82i9/3naz2G2TeXPYFLedux//Dix
WmspqsNVzvO7STQfTciBbweHSy4WxSurfkH4AzGpJE6SDfzdObLv/DbmtZdkWDfL
S1ywoLy10iQUggA7Q9EbLjFeQypP2CIZkFh3qrh9Zqp4JfxGJjJme6ilTLZLF91A
xVktMZiYviiBzMm81az3WfJCNsLesLSr2IWb0Y1hFMY2vFTtA3DDAfGOXgAYElCu
T21e++tWxzgLCEj18vUWHHO+CD8dA+7b4sueAtLtqJQXQF6dA/uDImbzFiKREXMz
qb0eDlrov6LsrGw+UH+yXnuzG/IZ2m195MHjZamrrO4hVOqdrPJLYvANEofNlXBC
zphGhyoULNuHLGBV/Ieno3BlLvcfNFO8jyk2HYFRkGhpq7v/RK97DwOE5mcfTbrF
d8QasAqrUiufxUGmcOJstZ8dq+UCL8RNLcdKJC4N6837tDSoTaPyPcNdox+aQsBg
H8bsupEZfzGmogjoAsuZgJny5Tm835/8xmyvgay5BGJAPcmkqVWwuC9JcMqlUCka
+3a6j3/IEw8hZdv2PVRzYxc0VYjronGnSXLz55jAYDCL0q2JgGlth+OVMHz9gonW
yEDIl60IM/sx7IPv5BfsXSbe7/IgsnJi3qolBPJTF7xMOecFpGwh1EBHtMLKWpyU
l+xyJvzGDMbdPwNQpXAkj3L1s1XqsHIULXwvQsaRHpMri4aVRg1HuXYSpd1ZxE/F
GZyUaUjlXN0kiHTwha6lrZN5ePhW8kD5BUoMH8CK+HF/hY+TRY3M65KmaLsmQ+8K
Huot4sqiYDvGmt8Og/UFbLXULTpswwXNa+6ll7Yjy2sFeDpr92AjDexXuRXA5JBg
v5yylcvOTL5RPH/pcutT2m9VOmyHg9mxnyrTHcCAGPqUT+wD0Q6QBiD+Ukb7Z3iN
Z4QPucKzLZLSuLHAJfXCJ9c3y81gZfiKHprylOptcmXJsWUhDXb6V2ZVOHrhZcM4
sJsTZRESwTciUki5Tjuu/7yKg+SNR1RtW9QIX9oOq4/u0Ivhz5M207TODa31/YBN
5ZB2QgUQ2nh0U463qpv0Jr6Z6XUMedSOqZewNjQ8NGoV/Xm/SJgPG+jdtBeDS54l
Za6tkZ2PZI9DN8QL7aOtcbDFkni+nfHtYHdbyMF3hu6x0+zgxoShIRbsuxR120rY
l3T5X3eAsd8pPHjK+TQcfgFuzANm6zhdcpyBvQNLPtzTOHohyWb8ey2aeHFTE/AU
jFUWasFiQ1ulr1tJpEsnq2fwRvS1jBqU1INhjVwqxrzjdaud4r74vbxpSmrvwhb6
jFhZIie4wYpNIa2feelC3KLUpVg50uyL8SXfqt5o4DF8o4rzbGiOaOf35X7/ARP9
vkzMWhaxMJjK1uwY2D/XV6j85pnvDL8OPcBBlYJ0T2vPEF9DD7uhqTzNmn3QMNqi
N676dOucgFrUTDnujPXAIb+iqn22/XaWF05xH0i26bmQDArBNIE4E6oQJm+/aZ4x
Odp50vZyL1IHCeqwTwMCp0q6zYRWO9eYxee/QGAgbdVZ557vo9YU1WmCMbM0tNxq
ukBK5yX6sAZH2HjRNf4e7mAhnDMdYR58o3q2s0ETmfPxua0XyhuOWN7Qwr7yggW7
mCIR7uqefgV8OAbqTnhTZu21H4MfBIx+kSAvDNb3Xjj6pgQCvInvWzv/Q6SIxzn8
EQMYGb6RlKIXvJnOqQgAzlQcPLcVNvFLIHbgDgKbJvCpARWer9U6Xxiu4stQlIXV
Zx23rAy1jeA5yUSbPtJ+YXJTizf6qKXggEFvobo1bb3pFy6oYIl34IWKqeT2nIk3
gsDrY4epvbkOjxzt7U40Ce4MM/1TCskxNP4NsoDFVvT07cg68PbP0v/2t2aQeQfg
oY3f+mqMWReWkD3w+wzDjNc/fAnVf8cKjMaSxiSFNJOojqWnnSUiFl4++Do2CmOj
opXaLAhHvKFhKDMyUXKmruU5zL5gzAhXJars0C6rbXqc16L2WtOB0XOauo/n/KuZ
w0T5uerNGQj72AqdOJTQNOWnHlp0mteTg0IU6WrzIuSgTHmxJo5DQGxnFoafvFB0
qoHpkytIAc5EcfnT+gd4dIyYc+oARfxZgOq6/xz+oYFedWIYoenacibFbPPEAGg8
YUp1mosFChjCuez10FKdL7ILTSB9eqBxmZtQIejGEw9NdRcDnZfiZE25MCDdkSti
WZQKZipUQocTUPTWLGg0rc6RH60ZL5m0uw0j/45FuXnhADBLpFp0MHtcUocTmbJf
P6Eo2gN3RlBQiTxJ0tv/fNz4MSdBbR9BLCxVzr9LBGXnrUnGHnycF7XBrGq/ONgo
dzdKXzS6zv8i0UOv4bxKsJdJb79Nk+OQghUun6o+YzN0wKIrW+i+FrTSntqhSrHw
pZOrYbpLBdE0B4dsQY1ZftwcCKXZWkYXiXeOz2fI5lxXppv+csxPcECQyCw0xRAQ
sFpSeqLjSvYESIKHa2/243P8eUrqrMk8yayDcn7npWfeGJrtx5Gq1JTBq1/GqZ0q
RiLz4e3Q/zbjoBmxJjliCGiGpaol4h52z6IGdmrgi7sNAxpcC1SAou/z5nlOZc04
kEbBE34Ab8Rd+CO7GEkSOpgO23uG9q4mvZBepwVCnQgBSyrg5JKys8F1utAzEf0w
G47Z/1/5CyNn0oiles5akb+iRqocKp3m37hzYZrAH60EXl2qn3fs1FiLaBm+vpyi
+ARFKbcBIICR4uUPpeIt662cXiUXhdmb9lVwnqbPMAGilnYZxilSek4b35FUtl0o
CmA4EfdP0PxuyhEuluzukTce0Uyg9dgjWwxF5v8BAeoxHgIA2DWcGC3rUt7ad5wu
0JrJSqwZKvxbRW9LTPo+YKhe+Z1lpJSWxbI3Sp0XOj9ZNZTVDVlIe5/YFblvEZ3h
6Uf65+NLciWi8xbMEpF1AuuKUzma7QsGvGFlk96oN9vqRIpckpxU/e2NRmVQAIHO
qdfcIfRNiSaMBDsd3J12urhpxw7GwK1SPKV5u90pt+yG+9AVxJC2v8+JTMwZ2KHE
AFTa6iJBX1B8WJlCcqD3guS4wMgKpY/OuUbaErLgAZIPijEfZrmz7pD6KLY/vW0t
95jh605LoKmfpmS+54umUo1WYPIqu7OoCV3efaX+Xb3iuLptZ2i/fBA2tLJeyEDf
jozSCmeMzffw80JObAdSTKAcbWN2tXrxbJS5vu5ubQ9191/37aF/5sAZnLVAVtfn
g3WEv3JzI7d9zZwKMDpuTmebaaBEDTy/6ZSq2H9GHJdPkxRfyvbifoPEwhWeWc6g
v/W4Hy+DukRDQJ3x2Mp6b0EuzucQmBDELEDEGc/yEBXHtvIbQI4UxNKtkBXVf7zD
pjBxgJug/m3/+MEdCMn4gysYcMdGFvhwzhMkBBrR+e8p3aOSCLOcGvff1IaL0CJT
NJZJP3tzEDPcjuq/i7KXzmOrFaKhJIeUL28GD6yOcI9yrzyA6C+Ac2c2GOzYxYhi
pvG/1jBOePQonK9YB9Wr3bVeQzXreERwpCbywyYVr/4z94+PW1zyHsEH6NZftFHO
TMkp4mrD++BZct9cj3O4nAKqGXYU7VIhCMZnjmbZ77WvPs2hjkvT72oE2GX8+1FE
89Iyw46qY4Fgv2yW2Fkh3LfbewECjke2+/D/PdU04uQH1NPpFQUZ5VndDeipVGi9
uyxd8/F9d5rgq428Xx6l5AhVY5d8L8mUkkdE4nZNLPiKtmVTt9KFb0SEvqcdsLk7
vGCjtk/VNuqJhXondrg828itWgGSLblK1j8Z9PcU318SwCDeEvF8McN6PsczzqKk
dh6gVj6oF08CQEqC0/hSK6eUfAniRnFblVPT/krAv4uJlaQXvjDbRWyU6DSExheE
iPH7KKmwLnqsCRkpBi1hxNgEbwmt2bZmMU7GSj++5jBrrSzPovirGCm1SUS2bvGx
v6btXmcyhIVbwl3pHWbJVFBilNx9I7fovDyv0QdilQwgkzQ4cNQ0IBX9DovyH5KN
1zdcxBHcoLwVCCSP4if9TVFKp0r8qLBF6pTCTVB3xf4aGCvpDth5VCKugPfmZ7hf
V6C6W3kuaLZwLC8n/oKB9ettUOmdrZ20z2jRkHKbWjNUvGh/+/ZZr+iem76V7RYi
WG8szwvUq3F9CP+nWa488sRWb4/FxE0VoaasBaKiho9DTGopGtlCAbB4KM5CIqif
r9OIZGsoU5h9aKtZQ5J6I7GWGNUNRqDHClyx8GnfN0v/NlGk99vy/c1LNsB53X63
D580KQDPwarGOMWl5uZM05ciOEtInIO0xGytYwc1iguaa6DwxVoD3CK72cWxsi/j
q4hFJjEziaApC7AQeaXp5Eaf+orDUua/0VWt8kNp4M/gT6MRneEbJkeuMhTZQDzf
m8wX7lyq25eyAUPjFD5EoxIge9hb7MV5AzfejZ/+PwmqCNOLFn462V1Mwy44sbWm
/uOUThmLgVWNMr8mf1x29jguiTxSMdYtzf5ddFR8k8/9g0y/vJWVhQa0cIG8JmXC
H9m62Imo7ipvSXb5E7MZBctdvjSmqOAyLdeD1R8FiLoHD9flzRBChosuzh3he9/n
HfdDj146rntaLca6V4CMaJz6DU8sZi/kuSKGSV+SCCcJHJzOPy51APjl2/8fyGfZ
UkXAPDV9NC/Dd1+Cbf6IwjNIOWSkxdMrc/RAS/Wo8OW1BZ+n4+skcC2KteQW8pSw
3UhQbyftR0av89WhNNPtglsp98FaW0PtCYDQpvKbvxTf1nLFQnkdg3SNTPXFmIMt
Y5YEgueB27cYJ8r73xbDD+0uBZXgg0b0FBoRlEsnsX4vUa1sOZsUCAAQkOAciSoN
g+prJ4wkeoAe8zG27aZETGsqEOBspTlT5F2TytBRNQGth1VrH20gA95J9WLVhTFW
K7yuOlFMACHn/23rRO162PzhGl7UYZqdcm8Zdpnt1xMIa74M/sIq2sBHdHYJ4667
UTwI40LVega36s49sFFGiEwO3OMTNHsxD3eS9EA0J0cOq9diUPceuVzzX4xnng54
Id5lTvlCCgRrHLu2qmwYKCPOd1LzjOSs6pQnlJlVMYMRtVuFEMch1+pSPTPBseQr
VLwO4fR91mgh+j9HlELFs4MYASlzglnTMyaGFd4YhncrtxiQrWL6Rg1vc+tqVjBn
EomhRDQkwUJD+dkn7i1meaXVijAENeqB4m5GPpq91cQELZlX65chdP7NDWwkk43Z
CtH5syDDYI5qd3A4BH7acTKwNzaeWnXihn16JFDv5A4YJP5L0Fp1BeHFfoaed3Kn
MKFkTbTsZh7dXrCPUHIXRfJ+FFueMq4Q1PEP+BUxeUsZ5hLa5dLsA5nDSQeIizh5
0fJCRhXD917C0n52ROyYHa917lPrMLThQLhoVEHFjz63ufJSErqm225qMLsgi5j4
v1WNbzAhBM8eYw8P7sFocuDeHEuu+jijlg958RBJH0/xKf0Z2ZBbIBsUDJFhHCAS
ZcELXX32TTgSYj33a8HUR56/c++9Y7ThelJGFS/JkTtfNn0naOtb91fWrUG7JBoO
ShNtBO2y49nr1bs2L8ZVqYGatBna/fvbMZEyqumwf8AtY+KEBrLUkIILMWEuNRFI
iKtLgB6yApp55vomR/uDAMXo9SkEXfpIQxqklvJ0leHRocborL1ONvM28PmR7RAA
eFJh3prb/VC4uLY2xxyxttRjHxZdGrawmWfuclJKhe7cgEvJfUNt5Q+T3IL8oIWr
ryn5e7zjPGsrB6FV2Yq5109BueCFE3dT9QxKQLiCXllM7qiQ7SwHTovAmpNsomyR
kZwhztcCKVZVlWqhQzZO6LFDM/pQIk4uOwpC2ym1FrvaRkB6i5fe9TU7aeuSVzNR
PNw84jQim+de21kdH7PVHkaGsSg+/1DcJ7RzzrqDY401YD36ute5K0tNUuou0hWv
dwqZpd7iwoXm8QYwYBhCG9maIoPbCcc5zc0BYswZhO5tCg1mMFQB/nmFgjWxK2yA
nXhe5+HMHBKgQuWzC2XdnstHEMAHBEc7eDvP2H1FerzCUUgdZeL1gAosRJMjUDmp
0C1uPDIMmgnaik/9n77Wz8YW5g6VEyYbvzTTW+H8D2Hh+FEjnvUQ75dUyTyTLS4r
0fw9iEx2NrLs71r5mapDbmqV+oB5bJcq9Y5C6umX58U1xkYJaIN9UzCKWEYEaN1O
vUBOn9lHy/5fYYAcqPddjTb7t1KeCRtMigvGNC+ozhlpxuQ/KHi5m7YDtNt5g94h
e2cKnlnVps6sWSPY7iPlHMqaalqwUSaD1wy44+0qLwZdC1iQJeOA5eilQ3Bdte4X
gS4Ai8T7mn5wf48+OVyZukIibOGw1J8zRlzvGV+w70gqc90CU5JuFyBNHye07iFa
B2jzHvMfWw0eDM1XFZNOb6SXcmTOiaexVImNhRfZTVrgWsPSvbklNj8Qw2QzhJ+j
yKtsUBnNSgK/YHPVSdl24Qd7UIYhQY2c0xPFP37Ud4f0jXQPPwoGquoGFp+Ao6sW
tpqL0ziQ6ZSefZNLjkSOp76U6vD0M/Puya76w3Hod4YgCR/L6TCJdKm9HOvl0RpV
eFzQuWradGNouxlgmWpXUMhQ1lDiiR9yfs9J8k/BMLnOSY0vFfl37E3mR/d2BA1R
cgnBEEuTHZ0lNUXY+RhJ1FtrOGShdCFUXTVaN/wX5n39nL/F668pOshDqlq5t7VH
HWlI8FIvJQ34b2CmQcX2BGwwI36wmkBFq3GuOLjXoogwnKbZjpDfyHSqdkcydSjD
/O0bufo1RUp/ZO4jOP2DttgvC0294GScSUD1r7OHfXGsT8fu0jxwQGVsT0XWOyCb
PxaoxdOJJFbAF99pU99kjO63i16S1Uh1ndUllFqR3seSD2H+xiCn1zaWio54yCfw
aYPESm6CyIrbBQI8pDFbtOUHydOHXPyjpsTbgSZZPYOe4ptQLjQxQRpTLVSyscKZ
HE3MCaZ4XaxOzVwjmEPiHWg9kixEdoOjxzp/P/O8TO5WCib4a6KdhfeXl8G+//en
uBgLqfgNMdXBnaZXecXMAsFr765YIV08sw4sSkX8ireQEp70R/rBtZETmyJ8u476
55ORyxe1um3HCxZfOwdbJFJT2Q7tRzqEOSNgp1JvwUO+wGxqiFCfLr0ZMhTRgjAQ
umUKGjtPurODfGQuXt70s0rGHQbOLsqdh7GHnSrzVZI9s07iDmNmjGaaQ2NywsJE
IVSRY1RSRxjEUCl8s0au5AEzvXUdCFMgOP2pyEiEINsAAWrq8ifuwXnommAY8bz+
Qs9iafQbHMhM0NOZSnq8z1cHla2HdpXU+4urY4vOh1LaXcz7de414lyH45xr7jnK
Tane8FMvRMQln8HnQoBOtsQKCnAFX8Fe6lMPzCUDIV/Er0M/JGgAb7JEsmLOTdBL
heFkhe5fVaTwHnRionp2Rn3gCIoYpOez48xzqmOIHnM9UWvZn9IqjyD1t4YbMcyP
+jEsKU1u85SeiFp6+iKtHp4dMOHayz1SkPULEE3Qf3sSIPyCwCYNizwKzvEbAFc5
VFOIhVKQyZ/k0Cnj0hSBeHDcUS9RFiYKRUvksR2RtyhWVCHKO+svnmHaIUsDf9xB
NY914wdzI+7VPzQMPzQ7L5VM2RTkNmotyZTE/AlGT5mRD+mAH1sysGJJuSqYuNs+
f/jTTxCg5W9iXIJQTxKCyZs1x9hjw53spzO8dtG9KBijre7UjuxZiB5QDIw7vd8i
cqn8jMMshP+0wrDhBFjTC2v+sBZkeIwKI79xkV4mhjHa1/nWCkfVmXt1ZphntYvm
soJJSGAKrIWchV4rSWTV8D3bG+nSqL88npMMU6fuEsJVs0unMh5WjyMRj1E2FeZ1
claXg82p6YorblKUM5ezGsaOPj5ob4+P4CkWxxsQykVw+PiFdlgsFkKEuslD9F7p
4IjH8tFquD1yQDva9je4rzrbnOioFUB0DZIL7zGN2AOdpbEa4254lDcKrL6eNAEj
r9mFzpQvlsoEXwUOIN9h4aGOaKMQVJn8CLIAMDGdSp5ff4agUpjRmSbmonKUmWWc
Dv6/pzMTB5TGWEjm3XtwUZslUR2Dog2SqSEgIptJgWEOEZb4hHOG5vA1wceXNwMq
R2RXcdG7O16yFVHblCypA4h9nQIRv07ZlK4IOisSkfiZlwMA139WlD2BfeeyVI1I
CZaoYQ1BWg77qijBSq5/a+scaYTRVpX6PbDtnXjQ0WpeZJOqSE8DvLSN297b9rcI
6fVPsYvTyK9bnZcY/k8F5s0XQshDrQUKfQlzgRoxmwlF16ogJkC61b/IgvhqqEes
hume0y6WpA2VK/wJTQDgWIdh4nOUuML1YjNKL2pGXONFE4gaLLAcvOfX7A8il0dd
5U22S0f6R++iExJ8FV+CrNFnx4hG02b2+8gO1RhRYnDL8Z+08GjTodGziNloEJZW
BicaGaDD1YFT/IWMQa0DgZFylZ+s6zEXohjON9MLcCeN+e5INxE6a4r07NsGVjE5
HDxj/YmTHiqjYBqc6VQMur/dqJH9wZm77pmFhYGiDsFApK4nMBgGvTei6gljZlyc
xeHHXmvfClHdNTUKuFHH4ODcaj2fPS7p/rwnMAlJ6bjH98DsLlXvKvFn54SSTzMC
QIcogUSBPjcnR9R/1EpMkN2uLhXKAzCdMX6bNNTE8rzpPlkPn1iQvqnBI64w9vip
YS6Er4kdCAC9r3lKL+W6jYf/U4YFgIoW89NDx133/m6tfNPZ0BPzcQdX+5Ysx9sz
5ek1zpA/4OOlqcT8ibPcWX1k7rIyvpgoXC4eP7OQ5O547MOwbteXH1Gzu/i0UL6I
bqQOTr6bNnFGMTqlZ5J+PaXqXbt5sbV152zsQTDC1/uzKZPiU1/0iXJmA1sAkS1a
goi/pfN2jhxVYSpKJWOjiaEKMDc6Pa3B5HaPMu3rS7X3epRvWf6RfJ73sp2XPPjB
cwUYGoeyGRJGPBFnK82ZZ2ZSQ6zg+UleNB8bOmxfhXvLOAJXd97B2W7LkpT0dzil
USX2f5241KZ2yDo7V9/N1AiJklQsoPxagl71NDPTx1KIAbkLBYC1UsrMwfo72nRE
voCHwOOyIVQugWHvMWDp52UIPTIdSSxHORF9J3ifmjt579PajzQCFyQ/xZXns8TX
IbsISehIRuBmwaZ6A0wFRXiAHBGZ74u47Nl4my5EDL3fGESGb47Qn3ni+t+9O9aF
Q2nmFYPmbpnSUajPHt3bzfmgayVb1iwGj8Z/XW2/vyoDBbRfqbRnEilgm5SOaIl/
yX6oSABYEPnT8XRZuUnO4zlAF8ZPZ2zq4ZDyx19x1LgW0Yij2msQFkkOyEryPwey
xCPJTbV7OVNiX9tIaI812Ftn05RY3zv3cVpSMpU70ac+KpN3Npqm4TzSAwctkDP+
BZf/mmOJswtYanvo7n8UaY2dvlBgx+8N8wFkD8siKchlmfWti/vrk2BXAwH/Vu7F
A+LJe0ZJvN6dUuU+lvtnEWLu1sxq7lQ0yXMR1Zkmd29ReJdXx2jEMJJCyYc5Y1a7
mE6fB1JVfGkb80Iuy7ANwK18k+PEHhOyisKDMnzIa5bSWwuSVq+8p4vC1RqL/Ni7
v/NhTPOOLRLTu1psFrvNEYjw/SONrUqnTY4i6RG3cdOpw5FyXC6EO9kc+uRk5Vk3
VALQBryO+6KSpwt58VkUeuZWp4dTcfrpVAyvaG5Pw67hU36fY1tJ4ksqaeg0Jq+Z
mnThkGzeFdxMobhM/HnZLnYs1rGEbBaN0xaMVSbiaCPxGFYLaPUuhAD4VFVQ2WwS
PlDHGX2Jmq01kQCiPRzdfGlbKS1517S0hqcfdJ81ZFoFZqW5j+mrRdL3/CZ+puDs
YVIgJ+xhWnbzy332q2n3VxNWoqZrMQjX/hcFvDuIAgrmLwvtVI08dadQ5ad4OTy5
0VyjJzJTG21WQcnDfaJZQqM968iAcaib5SP279azyrAE8xIJ4n3M6fA8RGXGkQ0q
bA7N3p7DSTbuMFm1aYwWz7eYGneVeI5sf1C76a3624O8IbragGb7SKOUsMiQEdCh
eKUkxV11IewMmYP3m/8YzYiYw+65rhABrAF5BoAIBc3lb1uvoRcItwhtDJtGftnU
QP6EUlOoQquMe2eW0UAIuRZf0MP6AVuVygXeBG0QTRD9CLzownHehE7rWF9qJhqR
xZIf0K8cYUlcXaRXPQ1KW4Zp1jATAVz1YB/QvtOZaAM7/9ma7E6KZvwwWDa2t/Db
7SeaIL9ur4OGtTSM3Of6lcg8+BJEYoHfYMnS3aunWK396qTqtSMWAUx/uukYz7Nh
OPHxt+CGnDPWg+rC0OwyOkOSOZ4cSpoPjdKQC99AzYhTJFh/MQ5gaWrynMMT+tiX
NVoZducQtoH3DhVeIaF18xh+WjWK7UH1ZXMk9tnrqzRN+r6brq+qYkL+6LLWWOBl
NVomIvGC7r4Yz/F9xR0+RoaXE3BU/IpTrjv1uOO5Hw94JYdqErCVQ89z3QkiJ/jK
6onDPVQxxjLnUYeQijSDEbzzW8dyq0IzOD0tfRKUy9o7ZO9HWfsXte60x8kgu1xU
wEMXvxvQJ5e98F/cRs6WHtFeJxnUN1mZ5t/wleTpO7BUTx7ecgbnuh8xWRgfOGd1
pSilOHk4iecQ/ChZ/lKXvPfNEn56n2P5+AHteD10E4rcwB/Sz9CE4azH5OhtNahp
YNkzaMcsUSe3Gg2tkwOOXezwKtdlpfmOPClIXWChSkkCG1x/uUAY/T7HGnlmjciL
/BO7dKzlMD3MDRRD8BjcAoREXcVO230XTPuVrZoGVyaj35MT5qAE1pIAXcmz2J9q
tzKcyNzZ1/hO8dXejrHuFzap82Twp7x2ijs/fFu9nfvMxtaYPdwS4/HXw5a+tm9W
DCn6luHnFDqVWjegcupFgLodzXDw6I8N9eQas7+5s3qLpzpU9QE3hKlfdxLhv8vn
B4088GVUJk7lzb++fX+jlBEp+pjflzMFEMT7gIritKGIGwm3B3wQ3VLDf7cJnctU
ur3/4rf3kQUjkL75wXTWra/pmEP/qwKvNVOlSYObt7Vi2Wc6g87tEB2BhlZIqfhi
WLlQLhbosWWtJgLKOooLQQIc8dxuTQDDjsANbwqf7ffCIRcQ78GfjDY0ZWLOYHov
Fe+ihxu7AP40978cUt+JbEHUN5TMJeoQ4NN7KsBCTyyViLETwAz/sHILlEJj+IBY
2aAlIFm7qrLR6h4fF71HwvvkV2lfwmLXrY5T95QoWhyzdc8vEP1q3NHwP0Lt3GBL
VJakhEYOeqFS8kOlE/qyNO+RijsMzRvCZQ5GBuDVUvdrMkJTQUjaRdnJ6HNn/m++
IvifA1GV5p/P8LhIZ8qz2nPjtIkMJ8NY2PYU0p5kHwz77wu7rbMdqaYtPtNoam+M
WWIudXUbS7eHnX1Q8i2gVgTDy9oG1jB03uRq95mzqixM3UbXM6t0okIXyo5Us39H
zmiNhyKnBSfLjPCsFMbSbVaCwSZ+tJqZ1DAtOT5b8HQWh7WNegGUj8clsc84uo/8
YbplxFKkrCP/E48CFBIjw95PRfvz3aTQomVoLc7CFnmBG4Vk9jW3Iuo7dtYTTtaG
U23UDbPkDB9qg61QnGT+ORJRSxHOYY3e5/dMREEBct+thJcxqfYibUXG3dJnKKeh
C2R5b3BHkUDydNIXoYpZZ+vrKr3l+LYSibosXJwaOl0MGI5yJA1HLp/hdrz1I5r0
Ow6l7wkhTBJADNZZPazVxe6Ht7OcBGnVqV+Ypt3GuOLdsDmG0o4+ommR52DilH8g
PInJ9WhxTkC/WHtoWkress8p8qGlV5krn92uxer4mAl+eYaf8wg7Csf29mFZA6Rj
R72rlS6fhte/hjXTBUd9HHu+MJIbrAw5JQ8EJ36d1xIIFsXGoF629TWg+l0hrgdm
2pXLy5CZebrNHoGKfjQvN69yWgX0iPbXBidkt/QRzIM/OslUNQVdXVBfQx8a3VZI
AUsv7yyCCydauwKv1a097QwiHtyiic9WnUcgbFyAatFtilPL6LeuXY1Oc/sB6M2n
54hOXBIYPfhVKoeCrZvFYVigPwa/grC+dTkvmFInJ+hJxfg5+hUzG4eKAViNNqo5
QZ06fgsHAmhi0zqNBsQn+gnek7QHM4kqF4wx7YEV/S/i1d644M4emTHeG7bfB02V
NHfzZ2McGuh7T+IfymER+eId12QONFslvT748NRJV44JS6hhiy7siwZH280WSd3G
xGhuklSvkWYAtPrf04JsVzm5/oJPIJXwVeS0uWU7QzvWWYpy2m+X8mcbNBgwElsV
gSQmjBlB8PuhfaZbrvkWLPh9+KPe/RHG7I3/waEqmnOY+9Bu4bI7ckLOPpIZ7c++
hwtsKCpyKLWi/ujb253MkWAQaf30Qr5eKUzKBhfEVxDTpCQ3eAfLs9aO52ME+hc0
9AJWr0t0wJQSiAA8RiK2X3lfLIq8S+iV99s63oFBOjC1WCQeSlCpE5RD7d/2Kfsn
SdYZgNtBUp3AKe9GKvUgAXShdljbj86lX+Kx0QgnLPZK3lA5tfwQpfKdSiQ9Iosw
DjCNFJ87GPoipBkYgtRqAcihqUOWf6U71Adc0tCed+54HJXepirJqR+qpFz7/XSb
IMbCxHkqd4YJ5v7YAu3UfgviLaMgC4o2QMC4GhBKJmbRnJ+ojmxtqj1ElrqXNx3Z
0LVO9qHD7qCdHVmDVO29NUBOMCvEUMWLSKWUM8BApq/OcQFZ6lkyOAZ7BS8rek8R
L9fG2tfj2OFqH8AK0Ubqx8Tcm8/xRHlKfzoYEWWIsLzy3fYsNyXX+slpFymargJF
bda7PpblEPpzVde03L6hCamEuuIF/019QR0C4fCXXjkpXKS6kX7YJfhGI9sas0/q
78ge2zmZvaYUACQzaG0OEtYuk6wp7tuPLxWmWwWbGmQN8BZ9Vn/r6yIbQjASVpmV
c/ISIhZD3c7AASF6tIb2bR2NW7mPMwKHBFloBEv5Y0xDnAQeCSRiwmm2PdJ/9XWP
8woowT32hkUBehprDC/k0uzzTBoZO+PRfoZZS0b36bXdOOdvusZH2KRa1jqBI7VW
BVI7JASFtsHlmjCjc2V/bNFdj0A8ozj4AjbCm6VJxN4BvMeEkVxx0yOtsNA2XIOC
LYRCPP9fM+EmEoC+52odTXn3nsH/nzi3u9d60RrjQHOCwqwa3sqnRzVxXazacmcC
8KK1t3VNGhpMCEeIeLFl9sGPAayfaO6C7bktFNewVZQaEITawV7txAyM7hFw2LEU
+nwPSeSHPBp9DDsGZHB+Fm5Wr6lrWjPR5NFcSHCKFa2vkUeeXK+BT3TWj4WWB3gt
EoZegbcVD4OJtDuvHj0nX4QGAV5mXPxxu6IRwe27UY5OkfJFjCnAZspbnvMCbxdq
EJhYJtUS/iYCCosFy4iIqqBXkXWc8i60wokJDLK8gel0wa+KtPircMnj2q8SthtL
+VlE1wBVY2CCmAHf5w2EzRkyilnwrS5xRwmTy5IXAqAxzs+p3+Bcw9jCkNTXxxmk
xDF3T2vk/V2KTfxcdcquAlGembgMpQKuK1HKHcpmQuIaHgJoUlGqTq0DtHqKjBtI
k3UrftXMCseZhDEJteehttK6gdAkh5EVx2iLgjeK8dZ+bbPZ71KPL3FRoBMisBwP
fO3akknHE4jy4bWcCLse0k06FfNcLWA3koz6icfmBYcs9yyiEM20rj5bDGyiVomK
evHe+pXxt3kjBuPIQfZvXY/VfCZwUymRU2fhMi9CcGwzwkmN9umsqiGw6qUiTFuQ
xE6oTkUXX96WERDFOCDTRz0NfVN/zX7M3qcENRSM7lVDYPaXVfBqUzULuhI5JQst
RLdeO+LYcWlT9v8DVbn+9oSxOz1qhdsGYEDYai5pd54wjs0x0JvDxkDGXbxuduBf
XSkNsR4BbIv09dpGgyr/+A2RowqU+tzGDlIClEByeFhC5uOOO+N9TOyYE1zrPZ4B
fOTXEsG9Zp7D6pp+GmUhUwK6HnZjnWjmG4tpBXLMxJCXMlcP2XiMfmmK6v+bBnSU
JfsghpzS8EHEkFM2hesAo6BWnOyryGE+G4xjz+4ybBvGj/Sjq1JC2TPljX6tP8oO
bcc55Ja6z+S+zs5vI4oPJR3JM/xG9n266wNo1M043d+KozMd93F8qSXZq+HYo+vd
IRMI1MO3dnWhXjb+VvvxPAflI9QtWT7jxU6ZH8/ZlcqqIyqCUU9rEYa75eDUYkYv
LpJTXjljo3wsCIxmd7PHNPvo+dUKRotVQ6ab3FpLgxXkMuNJRO59fQ+spu6ZhTns
X6y53PhRlemt4CUdkMppJbtkA6wLxBgY7CbqOlmYjvn6kNvRVwA4e0bbPWY/eVNW
IoJaOP7f0QRZE0AiKhsWmgtXgenGFAenvFY9Ow9Udz/SIq78ZnKRRV/IWv4Ja6MX
dZjO8iLY7Uv7qjyGI4Zu2S1Te8Vjdr7cioOCfEro222omRzic2xJyMXvNY5U2pOI
e4DGqUat9nFRlZLLSUesP9n2CHzgwdDh4wwJ7KTjIwiji7pFfua5/wc0JSU4vi/y
YOUKjZTSQSHaSAwK5c4rQwXO6I9gCszI1UFhONqSPKeopzf19EAXOeXpJe+0FEi1
VAbMrS5wze8Zpasl1Qll/ki/Mr5oGkNVRPrY6p6ksUN+Taey5OoFY9x+P+UMqWTb
KATrvHuJGsgp6PxNIk+eXEgjrtipALr1h0NVD6ZK339iDpeYF0eRCye7U79fXYs+
90QcYlqzRm3mnOozVZVTyR/EcYkr/AAJmpQ2qg0oITadJOTB4Jn4suWnep+ym1Ic
+s7kQ73oT1IlnSG7Y354HsghtMHwxOSSA1mtJVsyqyT9y1y6ptqbXAZyKAChj9/l
swwGRzmVwB7/0dFfP96rKO1CeAZxqnwZMRuRvI2KOX/H1l9J1ir8cfZuZeNxW2t3
IIjhTui4TjlS2vImhQowo3K0ihMm0Kc7EQ0Z/Tw338OhY6+6QtOQ8EIVJLHs/4G2
4yKg3zUbC1CniYP9RkxdlBGNYeOWrIpPJ1ql/a0TfDwLggRINBVg8oB4Cha0FmxM
ktCwb8kK6jDG8LUbrWvSHsUg+uwJhZyZ+YWKc/tkZ20c7GkL6aDPBZuAuk5PQVVF
IMUFjo55SSVOchO4+0cQ0r8KpE/jxilk+m9uBX2AhP7bIWIuiIwUnX9ct6z49oRf
7rc71hkQWwn6sqspVKoUQblNMX/zLaywmItcM4d4Ttj7CfuK9rqgXwgJiACpc0UM
3LJMObHPqSgqezDFfAberd8jXjxhURlHNF2CXQbtIIRdk36Hh1vx0M0XSCv/ow1V
1ZZBG3z6s4JGA6V7jqP+EAkjv+uckU3xuOoIyOThBDBNxMpBu37UHOUvD+Ms9/mg
XqsyC4kCj5wiMQBgLvR4h3hyj8TyCZk8Yir/4+Ero0ER5LFto/vFJ30iOP/yoYOj
/k2Q3UXUw9Mk0LxoZY2zF1TVj+9Dy0X+hHs+4+DHgDkssXM2kIrbrPiP+W1mI1+E
x2/cxN2E76cu861fBHxcPaRc0x86L3GmJMTu2hlysW4M4fdgXaLEUG+9ZhtwNCIQ
wjQ/NZq9wpTflBoywT2JIRAn0+STe86b6oZ0lJGGVkEQBfGjwyCKofUPyBDso0Bf
E4JqvW/6S2hPuA/hggRXuvTTQ++1Ua9OD3fdUEP8v4lzJ//m2QZGwBB8jRzfzwLG
JjAW/bejFQ4YN65DT7KurdW+KJt1i58JLf6wf48afZ1wi2LjJ/KeNmt8gc46IeU1
B6xyPvwRZMELpClwYPsd6cmxFoOISDCajy18rK5dNRXn5kqG8GA6ppnhz1GPjTio
TF+kiGeghDsKwwCRL4v6h3lqQOiSaPsPMX7Tglp+1fzOZcBInAQGSjFDevhB/ENs
u5/8uxO3WyiGf92RDctRKKS5s8oOTATv7nasEZDjB7fKqlYlSQOVASZHvh8OKRBA
mE5gSe4GuoRpJhF7UylRbEZ8mODdE7nibvvXeuh8QaRsyeOUpOO6GiGqqcoPTDJb
uWwM3030h6COUHXEsjEGycNF/oXOn1cuN4saAWfPJIl7U0DURt8BcT0P7De09ExA
lb0/YleY2peuw64DbTxvsPH50dHl0vAy+zcQAyOUfs3y2AwgZbrp8Va7rBeFiw59
efTXV5B6m5p0s2wOvfK/DIkIhoVFZoRmFeE+lqnLmROubUgFAXkBgcoGkQAidmFG
8XEP/hGnEweWOMfTTFElDJ4Vf+fSldVC1yfDltdHRZti45Sm82jMYR2+HxW6gRgX
1q3KyemUo243KYE9JcWqPKk4KmKafEKxEYrp7hEyFDxOfupqgW786W9klveC3tPd
gDujWElgVtSCxzeEuWVG9aCnfNA/00k6gz/TBx4T0sGSxqMbMbcTUYFlLWrYD7Or
674r2OsEkEcVZT2qOdjru7lS8idN/c51hSm34kQG3y3NVR+kMzF8bBuJwbz7mCXB
oXMQjHJwHf1EGWj6qZIm5lsXvghctqV26N9to/0teqDeJt/NomglxSwl2/UeRH3M
NgNylHJ9aFCswHA2qas78ooiddyfp1KR+U8dpFcQjURvc3rm9mn0EZnKUNlA+aBD
yPSOyO31xwfXlG3TTnNrSxRee5LkIWZ+9/VQTQYEBE63fo6joHG+wjxLUfsimftl
TE8tpU5i7IpxHoW79PAZjfMIV4iRnGEgBXRscLkmsfsPw51OC4xRzplr4ln1/es3
+1uUx+9tVQIVggk6JOaYOsJsdfAmxMJaINuoyLaqtuN5LBF3AzjvNg6tIeVMpnDx
/WurhEHDWgjcyhTU+bMpEGjt2tn+N7zJHzQcOCl2a2/Tj9TOfx42T5nHYt/pDVrG
/0ln3aR88q4hy7ARbnj0RaufPBLKCA2Z4ncBkQs6ziMtTU+wOMy2OaCHDGdscwm6
/CNUQZ7AdZqlni+iZMHXDnmF+Z6RMyKElWQIe/plQwoLpkboxiQCnx85jgYG4bT+
tURv8U79e3maXWm3nMpKoScKRqYzvKuZcHilMPU89jSr3ysf1W+reUVjm9I5MXnG
7MPhTpZQw3VWjbwN2JwhHi/9JlEKNGMtjt1ksmZ+5y3gpqO8EG3AKV8OaU6kGUtr
WxIl0EYPLHnQl/GMTJZ1zMOhFYGDMhZnSUk2ZVYnZmavvvf8UkjfHJiWk2Wwv/Ck
2j873C0KuGwN7k7UxSNTV/lL4jVHPKPGrEOjElHIQi/XfZz8BhDwJHvyiEcoY9qb
vpDuSQ7h7Lth5/gTfra8DPPALhKs2uPsvDGpQlK9aEWBhsWDzHOEsj2gIZfyBB7h
Vc3m961Qf7hpRIg9Rmb2B+X7QldrzlrZrsdyyC6QN33y/aC9QpkniRsJsMRHhT6f
GL6nm/sAn/Fas/jgdmlU7IlKZZYgzXXrUw1A4cOok6GE3F7jAY/AuiI90qAMlnNK
lcKmRA7JT7QPJR5XD169X3gkDXvW8NJZ3gZBCisdIjNwlnEEEcqFjCrSFqpKyfOz
8FJzRS4s7PzajaYJYoXlIMTG31mfKULLrXgHqs8ZTJ8FOAY3sOXMR5BkIje4kRBd
7li6u/nHaOMxm7/L6OmPpshlPhY30yubrhIMPzntEZy22Wa70aS0zJb3gD6+gDfd
fa04dOF2vofozqEUuBX2/JuOcbsrrObx1W9ralZatN53cymXJJQ1mPtpSsbKt4pi
iJkG6XBywu4d8hqeP3kdn7yGUz+E/C6bMyrCHPocOccMAH7/PVpUgDwO/MItC4mm
ZGER/pmmoSMoQDojKzQFS7anqKxZc3pDjYrHu1iNHk3kerg2AVFHJGxFvp/rMv45
IEw8B4q9vi/7dOw0dX3/Ju3maXmMSoJztji3Q7KNGKUhDCCggpsquC3GIHw1/5wP
jE2wHMHm2na6Rz5bJMlHScgC87sL3QJ6rcVbZm+sg6jt+2g16tSofQRfwjGaIgsO
0mOmJebI6J6iFwb4Z2sb8j7iBuNZ+Ui7fvdsaRJkMzQN+iNxCabww/SQW0NjPFxy
xD2jlrDzNmDLoRb5KfMqebK2fdiIH1X36kK+7vcd74ilgTSrn3b46x5bXRHA0VA6
wnq/Yn62gN5N86Ds2L8hQyThtdkIC7y5Sh/nugPvraLEKgoE3gdNI7QPXtySuNaK
UT6bXUb4eWnZ6WywdIcNVZjBQCrdHpD15S5XPvftpuj6w6peWbyTC+ehitizTPFi
cl0/SwiGYKV4SwULu6ARi3d4u1RI5SvD9sfLN5tQ7LsopGczvA9ax6q4XaFH1V+M
3zBz/A7TXeomv0BxQV8dBnQ9dincMyK8nc24hjbAbp47UlC/w5Bv7VEQ25N7xQM8
mvngFnK3c3R6CzSltSVoilbW/YeON7OzqhMtS04PLDHJxfAvGDFO3a9rGcchKyE7
nzsYjptpJo2iYeCgV9J4rphFA4E8DNgDHhlglxZn93iBgEbp7K1Ovb86Au1MEsp6
sqziwBBEhTWZ6j8Qph3iQXzc1iuujXJ3E/pQlrfMACKbcXUmcSlKRTyMnSg4EHt9
TDnCiBhhnFjbqz4ZFJlyC3jL7A5+aJqZYJ7zl1XlFm8yVLs/5H2CAz5wmUNoZM+j
8l64s30+aRITWuej9CT2uGMRtRsjd5O5NTMQmGVcC2tdVShphiofpfSMgLDiW0Mh
HeSr8nLxBPeCsUBpjlQSjp2v+izjHkU56ybcp4NwVJor9qT8NheV8hPDMq5a5p2N
bN4oidt23Kin/JWfdYwO4pfUDLWSNzooRi/IciagVy3ZC7ork1CRaRwATZIfdf8t
CBpsoV5U0ABkknV9YKFFuoa1gUNzFpL8arrkgrdGiiHO2zcA/PlolWz11A7X7SnV
8lf0/dJHJO/irh1MshtMdAYvO79+RoQ4BSo/pObiR/AGx8bTqUADLt91VXE12wYo
aqVp94MGtiEdtMrIW2wPslvs9xSRZV4cvOFHTYni1gt/NCAo42MxOzCgGFmylMSV
z6AQC7dDMuszUSpvQp9NCh5dDuDzwAQA6QZIlUTGWkX+jeydT6DAl+HLUFRKnJvh
/QE5ew6xb/mO8EpzXpgU1MrA0aXcfO4PnZtzY40HiXwDpxud35hQsTRBrLIPHHKz
G6fyVnCWKRSxl6h5zyqSOWiOMhH2R5b8QlFrYSl3Z/w3TqSEVsuxfzXJ4mYv/PWB
WacNY8KDcXoq6CyXj4Vl3yINNpLba5+YRH1U1dClkpkiB+bqFz7b9y24y+Hu06dq
kRMafq+3YGFfZV66/dRmnh8g1NU32nYRGj0tsSMd4eYLB7nHsrpcXhHY+hMMjO6r
RLjHUonpE14yGxVGbTL6QUZRnlkZe5ZvJsTppuvMIMndSCFITce228tOMLq+xiHe
xLeQox4aw7xPYTNOy4yaMhu/9u5CDRGgHBxbMKup83dzH2VJJXwpm2cOY9IAnszp
7rAZWmcCB63xqVnvfKSibXCq/WC7pa6h1J2vv0NRHTsjI0anveP7RQRcaSldwXh2
n8I0wfhD+/V+1yKopFzC76ig3PKC0ZQCEPs4egfJX8pwJ0WU8EjMI9dacx9OMlB9
KO05/a8bNTE1ORK5cqYm5ciQg0OIRKkDG4eVuygmXced++VysUxvC5sJApy9LqAX
4Mys98DAAWKrqQfkuz+4nJRHkSmrneUFXdy2kDEvhCV+f4EZNJljr+1JnFjMHxEA
5trTfm+0Mc+t6aEcy8yU514V2ibD39cThFCIle8QhhI+cLdaGIKWBOx7/ahTfzOy
q31E7AbIxwjirtJVNwBRjq8KIFGEueJocnYLzaGPrFCy1qePknyMjJrS0lbnK6on
r1gL6lCf8qEKiaDRFnpXimKGDxLnJaldyHdprDXutWCpLIIzygMkq5aZnu5uTAYe
9t4hjnQxs3OSSaJgwJ0Jz3fE0+BpV3/sXuaGC38GYx82WxywHf9jv1cE0N/ogA8M
EjUesVdn0QlOY6JVcqTp1FDRYLQyviSCyRihAnTQquGc3+fE4F9iRYCuBGabtYrs
XSI5bi73uLu/dUu95zkHwd0x4MOOFjVjgZ1kpga9MUTLZFZlYoy1rXVtChiAPteB
WWyhzMPF+jjBJInmv/lQ9vFh5UjlKwWqadpNnHNV6ghsxoUwEdLZ9NTiXe07QMOx
azsJv5wx/HoLpismvDppPQ+tZx1J9LkkWf/Jx25QCPTMUutgc55vOSdyv+L2lmIm
0yxtaLBot+y//jq6En2tHuaACfkhOuD/w6sGjahaSwM2Kfq+5bSn/lhbFGpfA8aN
WMOHheGJC+hWIlpdERhrKlTGciGEY4fbQRXMWiXCStuLSFHiajkhu8C5V0cVv5tH
JPxE9ypoPaxnfKIaT07/kCUeMYow2AArNf6xQIknJfflw1vjoBtIom3qEMi/UQA1
Yn7JstAF7xuPKQNHra3OCp8R2m8qb5Knsk5gTDudhyRqfXu8IgQ79QljzyHHYfd9
hZV0xtLc7TDS/I7kCAb2GP3+9q2JOou/TR5LQl6iwZbpv/UoLjuijLrTCyEm/qJs
pT3BiVdgDr03Yhcg81VTofrdriU7Npgvw3tdYbobeQ/8xni1e6+C+6GNr6C1z8M5
2S8oTZk/2Ka8IIqt95Hr/MXXggABF4cboRB7umUmfKxfH53BC8tcbck9ODcE/dmP
TS29QK9P/43aoUHp68KZrN6XVaAtkFyEwE/mhpWxslOLLojAgQOJfT7zVZ+5Nmn9
yBxDA56MnDjW5fIGCmIThYcI3NPa4fFzF67GVOGC/k8XjzEsG2NsfRdaMBJwNaPb
J1u2pB5mG2BwPf9PggDqtujEejser0Sofffq8Yl9oFM/xeZerw4vLmmvSDp/d8i2
10ld87ZwauJ1WohDDnCvkkucj7iciiCddWp/uV0Q8ytghFvtRjjSPMsPRhAYRGTv
8dz81WHquaYh5gmlarQt+U2tgL4srddC5DJmvh7P9ZBeygBjU2RfQutSUtu6a1IN
mYgoXSB/n0dUiLRUPLrpsuSLij9zjjttcIi1CeQfuYH4eCgcUbuJ+kpYebmqBzqT
Yh1IBIP7EFAEQ7Ei+8zXO9nQXyzfVbnsBE0qknvdwbUxqP/n8a0lieLmLKIZyb9E
cbilvHfIulLxDhdgx8Zb841zemxbt6YGYAg8gArQYmd/WdIYdsJ5cHLw4TdJyPPB
MJNYBYA8XRJlPxkyBdqi7D32EahxspSwQf8Zenp1X+vTKfPDhT3KR7/AjSzN9Efc
PXAMZXbLesbNRWq5PMrnNqXvlODgmDXLm5bWK4YzECCB2iLgySWI13CkYQcGFTGI
1vcYjFTGm5xLMp9qf5qvCMPEoOfVB7itGXHPvuxD4GXFcN/lOKeatOJpOMk4wuOk
/eSo42yqPRI54VJJ7EdGCt2Jl3FTEtCIblkebEebuq97AX8n6fRkTC6n1YEKDCw5
WePf96593EgFFCnoswoSVhJoPOS5miw7TmY/LVKJho7ig+v2i0aekMfdqFrZlCMk
CKr2C+7t6NpqsQ9j25tb8J3cnm6um0xWv91hIdITRxVbnkyHeOUG/ctPc+vU/mxe
Pb7do5iBdBCZljVeYF/dM+c1JFTGjK1ncR7gRPMEYY3uFaC3E1vEYRBwGwul8KDy
3PhSSPDeIyMXNwRCjyMYqtejo0U53AVx6w+a2bQv+J/yhUJRT7onT89Kes8qrgBh
ZAVv6EixR2jZ2bXfvAEMxoPcjGfi/2SyObI77ttuDDe3FwPnBN7F2Rp8Z6DyUul0
Sw0i4yD53IYUw44+IvDspJyP+k0M9gCbyxZ0OyhyRIRLvvOSS5+PiJIlFYdKG1ba
ELNJKbLzM8212T2k/KVodFwxsgTtw6vaJDIwGDtJFhXZU54iFizt3phHCRHjQuHq
GT2GtK+ZRbjqtZIh0szzwtpkejFzBvrdbSp2t9p0x1AYn6AB03DFF4Pgs/JMTINi
wffaa4rlvDx6Eg6W6YVJg1iDEffy4Y1NsC0dxgxCRjoJei/Y4ySw7Vlb2/QhymID
u61iejV2FkcB4Kx47Rqu9C0R6+L0SHZjxqZ42eAfiRooedDUS7oNbz5I0QjTJKdh
AMwK666EUAUxTCaB8imVi/i62Uca+uZU1+eYetVMhCn4eklGOhV/NbDmxntoV8X4
+f8Dp+Rh++Z3tpOFRLNO9dNro8tiHWrW/EqPHjTY3JmtyRnPLlQNbkdYy5Bxr7PA
QJvDlZ0R7G3GR2LwnQp7tK0PexxaU0C4uLopgupyPIfQc9ftS/x6KtXsMzyJ1qT6
Bp2/ceu5MGt7JgKR3SwHBGclQ8IGqk4OyyIpSnqTVk8AZC16AfZCEejzRis3FCP5
HxwhiUfsXmtr7wlrhMCL0u1l9qQgOtzU/hD3RbRbTVN+kv2boWrHuRfSJiyYc4dz
VdvgLwPoGrr3EbZ/angIk0vaP4BhUKtYE5E6TJjt7E+cC7fSSs0DhdZnWE6F6RhO
ZH8DJJjgI27DgD2IWer0n49GXOdKRpCRMQu6MEDLarnf//zzMzA8I+57bg7e99Qz
yZLQ8XX3/a86acylsptD4nvHTf17yInvwjDoUTM4eHOfQfbDNopPs3nDzox3UJKW
Tq+vqrH7p0Kq4N2YFFvQdeXmQShK6TrPAZX2JV0YcXjcupGnIEjVnZPG0F1NgU2w
MN0+1fY41waWHWnJCQnOdCO+AERvrvE99DZtyhUISnZJE9LzvxOhaBKo5BhIWbYm
aqSlxk68ZAL6zzOfUNVq5r+7qogH44E54ujqodVGCW2mDAILfzoYSJ3VZDIXTk0b
I+6WSP7yuHnh1hTlV/mp0vi+EoYKJ5adcDQVt9dVSbdcO0qm6ya8w0mJkdhj+Bxn
FlvrVYppvwq1qTlGaSKtTVTW/XAMTma85A8iXIOWilS3EXwDvXyjBPg0hJniRkKu
B7Wg660sblA4ax0k0Zqa5ITeS0yRqzQLSuyeJC3I68Eb3gEnu1JHnDs11AfiRcgc
HiXYL21Us//ND/OH+BibyEMqxVwdPjboG+uqWcWP7Vq5rOS6zr3he6bZyCbBaxJq
SrLrgI2DxYqrerP25xclUvLs5ofNBhs/FvQHKX0FgfljzH+O4LwQ13jbf5t47sHP
jiJlNjcUGHQlgXJ4bJ8gezgNR3/lyKZhFlEPswwe1ktV7k8WmB63YG7Wg/OAN9ea
HPsEDqmYLO4xSrTmQaNiqv25uuKSJcXKLYjePAY9h2uT2NL2nP9P86JwVUYgLIso
7HjbaI4KUNcoz78u/XfsI0vozai3kMns49BYR7thSeq7NcY8A1rycpLXY80udStg
cyBF1yYR4VABC94UCKwvJOfryYUf/rszkRs7L505UHZccaFeKRH/udChzA0nHC4C
pz5Y9GUCCnRcQBNVeCDigkRnw0HljpkdmQDeZPtc8qATcI2Tm5wNmxSok9JoDw9J
UEX2AHDcZYg4I7Tsube9Vq5jtTPHZuiH/CxcM2eMwuqL42KQF4go0NLdS9YlFM/f
3JRDDc272nRIkpcOHOvBzl+mc1TJ9G2x/lA5C+eL9GA+hf6gf4RkVLyJXmQ+mSAA
3WAxbbtFHEjkYcO3itoj3lYr2P4IthBd91Ix4vfyQzG6j9A7irmftZIlFzxCXpHY
HFgFtQMUv2A/m3veL0AKS9/gRCBBRSSadxr+W1sSdKaj1UqHFlSVM9jGwPPSlyy9
JC1NogmoGN6WZT+H8/+QOezydKsHHX5pRfqYVJcQtxnIr6nrcnGtOq6Gi4jbzqOv
8yeUA+o89e7fhZFq/JSGh8iIsGxXA5sniriTQ2VPov0gO0pIDbJrSXpO6q4YTaDO
M0Gl0iHmRYoC+bBo6JF9ymcCAigFESeWPzCMFPILH3AwFZklZNir0HExhFXPquqi
wIAjyg+Q2F6rr3ZDw5xzZ2PvEer9JyCTK3jNnsCweXLC6XjAChOSWZt8FydE3zF3
q/vz3r+f5kcIWyGOCMaMv7kMQ0xUfDYwROD4IFIZvkH+LUFHpQcPmE4InqFoI1O0
2x97iySjlc4s9VqzjZ9mVBi10QA4KO/+NxTr/R0S/OwBNUn+IRwx9GB8bsUpn62t
pcjdOcLiLic2/FGwRjx6111ionWQEHP0x5LNmYTrx2h4LNvqteoreNG+Y13X3QK5
QCoS32+K2NtZHTbrUZ2K8pkQZldMeUGRoapGgrwymNb9YXXjLoNnVjFZFIgo6hiJ
gYVJU8IiF5ZILUXhwK8e13zpiI/eYbHuiZnVIXwfEDy1dj8RbblJRMat9LmlQCW9
oO8Id/Q0q0ADbqN0GncowTiIwFyCm7YXFhU/evkIVr9/90nfEwTQKJKcxWVdwUS0
Q4g7FKI9pzxm62b4y5J2laAeXgU7TOF9PU2O1gawgp/HSUrll/3ciJMKHMclSX5Z
X1BlrVa5LBFWviSLgfAVmhIkuw5P9GlXqTo1sQIhQ4fIWS0RVmhEzD2ZA774of9i
DBcwOHt0ka7F9heUhZmmquyqnRGIH4cKHjT858byXtqbPeQZNdJ8TEFZmEQhYoXF
1laB/F03YW3lQycaV9K/EJUpW8W2n3r6go+N4eh+txOJiNgd2BITl1zu8tIODO+o
pJndM+6LvpYsuyi/4H5XJtYkH7oA2SxXumcHN6Cb0Rzffgk3WfAZA1fkKBromWun
2I2CcXhDQI4SFvzKgZgqormFY1OZSKCBQeUrvWWpZ7nJBSjsd6clO3kN4SKMLmAq
tVtAo3FnWLvduj5ijLuxQDePB3r8jx9KbTBZ2SPGIdUIvR9tpN+HtbBxzdh2lnmd
KVQHfNUirCqaCPJfkVndujIAGNHgnbv2JTJuTQ62y1eTr88RtQf17wWZ72Y4D++r
HDsnpwBIgUXQn3VjtimxHPI2D3JGAKd+ui1qwi5DUQu4XVBr0o0S7ARodo3eLnEF
t/uuCUnbC+FXcpsrA6iWnpRP+zkjiGehcq93iYfbi5Ax4JUvbgDyIIp8rIXmTse8
oJWYEoIkJ8Z995wjBavunl6S4X6MhNjSH5ydHu8HeCM7w5CCUKfPbOMDti9CP/Yn
e3NcVajWZApZyfEo2N/L7C3j/OgiHvCgQQjR+FR5zVhE7bjrRqbML7NjbH3KQpa9
QGEDIpaI91QTxGBeCvaoqsAQjuaAYMhATzqfqOm4BcRBREPzLy1aKBU3oKRH/j12
IJh2SvpIPhJcVNDza11afD5lZp7/d92buLA3U3otYENk7mCBRDwESgTQJIO+J5JD
dhyAnoHGKTJjpWa1LKAlz711/y/GN4WbzgF4roszKmUjBoo4uFWUMwjumNkGKyrF
wX81e+gLCkXlO643OS2Jp/9KANVh+E4XfDDzZwwkHJvaKBqVkLFlfTKtrYsJvRwi
yamxJsHc68NATeL2OkGhmcfb+AhWQqAZ34By6B46xRN9doMgpGxHsePwDKkubBx8
h1nhKqCqYHSzyssFtUQ3CgfuqXSW5Op32ccTzro23wS1oUIjjjm0Sn5rRrrF0TP9
TUmC5UQFpLcx58wPwVdNtcHnuoAUP0zvckOQy/rj5xE5yQHZL9L4ClvskcgyLpUg
S19h2y86tVWdbX+x3EbUTxA2Re7ipvYfCxRgMXBfYU5Axb3wrSgc+3620LYddNf9
DLa0UlgklOtArCoSJkntYSvh3e9GdN8nCdOPg7aaYD9IwdSVmkc6r2cLyDvJPJ0A
kg3kwgqDln5624aHF7Hs8O3tuIr8oyzZqbR8l/afG+D1Rd+Bf2UgDIjEkxP4di/D
30eHYdcOPswPZzJu+50vb/CLK74TpFYVULL6e0zoJ+DUwilWZFDQAh/SCZgskx2L
0eZFxsK9tqOkV2pAUG5YaQ8VAp48vNcIHe8h1MBY3p6GZQ8Y636enXuI7vHKre69
VCpya2AcxiArLzYeCnmHU93OaLdE7wUmZoC9Zfwiea3FmWL25xdqR3UzJU2hZBo/
psqPq+vteedTPXHeOlQifJjj0lEVv7ol/aA6ht4b34EIek8nYZxtKi3/0HbKaAvg
3V6jzi8qMtwReaaiJon7O9j4bQRUYyB6a9nqrMDUT+PGrSbb7nfwaDqMFi+OwPso
wAvdsGcIfFGL7xne6wCP4Eu2sh6Hb8ESwsdtFB5ce7MCeEMwTJMsowy6oGbLyq7x
Kaby/VDqABpJIPujIEjec232BMP4qdsbRzf8Dq60b0M+fLEbcNYaX5i2xAslA7ze
ORMnMwBG7Pd59HVP1EjzliqB4HeQIyZ5hOfUBCpegu3OgyCnlk9JiQbHJbK22ngw
Y+/sYzAROgvJn/XOPMOGeUq4b39eB2gem5k7BKHsRWKw+Me2lVWnkyexd3OKW7C4
ShLKdisAWwBndrR1o3EaHgsxZ4TANeRqPJBSVZRyrizG2XanvJDhWH+LXR0aEJOH
Xu+FIKefQxSGyTo/ZP6Il50wsQ8WHpqE+NeVodH+6HwKgf2nxsPsM46fPX4avpdY
25AMHA9SVjU+vDAGtdOz8+PSA4AjeEnDMigqhLIO9nv5PVUkgd86wqEDWLVDqYh3
eg+nlx3iIMCBdfR/sr0LYi3qqMaeDyrKt0w7vTMcgFIUy9opQH90vFGKRjnUVcHB
EoRTyx0Lewc/vAa9ZIEC8P2hb2iQQ6AtrWqjSBuvGbQ+0i46h4u6VP9uhZMdIqxU
9eHEQOMD9fDwlo1as00MjMkUR2llIjI84T4XV4BK4A0GaeGMT/YVkqRXR3Ymrxhu
a2QMbKZXI3Jy9RocvL8zGy0fNWtfhVSWw5z7Q0Lpz7+TcxFLsNlNItv/aCmGwo7t
jpp7KKcm9AsXWrgVGeaNUeC2aFYPFoavSfZhVRcy2n4w7vja8acV1PsHCQ1KRxM4
Xb11ZFnOdY2trxQgeeAsqSniilx8jY5U3rSjzcCxGSLjYVPsb4oe0fo9hnhK9PDF
gktLsIyaQYkqCEj6Qy1TV8RejeQBJ2LmgnokKptQjJ76XbEqwEfpwT3j7aJyOX3h
iDg5BjsIez//xXFJ1KdMJ+uFWCd/Ma9YkYhdpkimQcL6CQfNB/ewXXaNVdOxz3Um
DI7yRpjONa/jhoOFx/pCyZelSnOKHtbHNfM/mQjnXzKBeA6VmJYCzm5lwFNq35cQ
PfUu1Hli2pwxkzTSJ+v59z9bM6UCw4YuTMgS++pd3rxIyz0Nx4H8KQKCepcCIiD2
rWcoigNOIvxwwyq4lUq6EkZt1KgP+MNVONXAQyzJCN9CxscdX+wiK+dEnxkl3J1V
BRz+f4GXmXEj8GKj2fp9qh7C3t0CpTJ9cRmFG1MO4/gIyjVzZiRbOGZo9MIqbMvt
QSSH0CIXWrwiIGkLaZ4LnDdtqvwbzmuzg5hSqmPKE/drUspaaZEAn90lk1MQezDI
wFf1qoSK2Tw3oAr1EDg/B22lOIlkdxsTCXqlBtEL8K9Yz141BfxaKbwJTSEocKUA
pXsnkilQNV3Rx6wJZItGYyFMTEz3rxg6EoP89S2eLaqAMFULBuhShmIZXly4jGdh
WVl//YIgBYBY86BeclhvybtH+C0b+2YRxYipL4+MyepG/NcEZlLM3IGY3tGlHXDq
eZsjARD289zfHesYjsUSCrAurJ7grMxJKetr0D7bdG+C1K6a3SQxJkkalw0CtYT2
/KvoOt5T6TvB60fDZqFjDjcgxBKM/p1gd4QoLeUfu4WSMRpcBVInL0+9o45JF54q
0rrE9Eq59KSG2ZMWhPNI5uRBiH/fZe0qu5nCpNviuHOf8PXJclS+Fak21iC6ohsv
Wsu6wMNOYKBHddHzkMwHCXM0CvsxswGNtbLEivnIZcyMOP5WCyxQhBJBBYp4GrOP
K/GtIfxYmklPoiBhaRmiC2KV9NTFF/TxEQaisZyyLzTnXMvD/Je1rqhMs6tZLqXX
CWB7X9cXk05pFG3pIxiJ+T2hXQ/aa8b5Qj03fHqbJJ4XI4TGvDdDBGILPyihZFlq
K2KnV2EaHtZPfg2ChwOGQa0dlvHrKXF4NrM8eJIgwfuq4v6q96JIt9Zi+it0wkQL
G4bzsq91NqRjCYeyCnbveiDPI31/jKwfUcdOjNjYK3wIjDQ4sxff4ibUynKJVsoa
CBDGu66RhsNFHeZT7a9sO21SeeYek2IfFc7nT4ye36Z1iV1MObQsxW1MyQ5hcBqC
TNg07jovVeDJHDySilSAF9vWoIA2WLpH+xSMX+nop3ZGhz0zO6c9yBe0rUY+T9gg
C25mEEw3KdS54eqW1SNL2gmI21Q/+3KNH/HnT5JpCoP++lVOBujhtZQdn3wF1Zqi
jyHQjTCx9kb6Mh54PRuRGoL+QZ1krIitUmBiMSUt+WdIdtMOLPKLyK3byxcI0kXT
MUC2G4TDTOLYk4NhStZ3THbjfZfbPGmqgDpFQRgo07H3biNHl+KCgckBpaeV0Hha
EXQ7F81b8RysG5yFPhOmAmENusoU5uMwQtNTeCaNMuaMJwaJ9IbgAfbJ/Jef3KPf
Up33EWC1YOIUJLDncKkp+mX68z5YqeyqcDsUQma5B1bgt/Iv2LZ7uLKFic26f++6
c615VZ5Cy7RObuia4P5v5b+0CDZKaO0i+WcRndSiUFxM87exxJlP3QQMlQxRlpS7
irhO5K5nme6P8P/gHZdA6a8TY9XLLpW3yycA02YKDZLDRRm9C7NGbRQfmH7UOyTD
hCzqMlN1pHIW0M8n0vDq32zCTwQq/h8qDvFdrJG6LcjLVrGWmO4el2XIFJxxupbp
lsngSu/HSD0abXj63nAElvui6AuS//vCo4iD//pg2jDK+S+/kWDvkCMMKnsvNuhr
7Bz50Zfwg2QpOH0mPY6iBrXNOaWwSs+yujN7OT4PlDnDizwI0OdE5s9ZvuylsjLL
vOQqrplP0S3VFvHOvlwmqdfoeAUawc+kbtEshl9tUYxwDJHlPJ2aOiEpItHF22Ha
Q22fmkJNeIVs/G0UTWhL36nXJ171tJthxJdhvDmppxU9v8ntmQwXSuScNUG8b9fs
KPr14p9IpupXcqrzIJuN0K7uQs1kjl3oTi3wpNtEq6W9KaBzOAX1JwRz97HOooh0
MMZuD1eF5JYKAflAjoiuP9CP1OZKPhLVgwGYCuUF5quHlMQMIbCz6LuZSB5q8/vx
oixTjRXEzoETsxIcHfHGyfOyDCbbKgO5WpMk+LTKUclcmem6wQefjcZMnxuKRxTN
R/zQGyMKILLNHsPMvXcjx1hpurmc/NxKakPfxbkwjbfK022eaQGckaNdb42e8448
6Dvk5ShjlhprdXbwpYDDABGMacrM6MFjyrbxJnySwhmlPf10mGpsO23BOllr6/jM
l0ZWRx/2Kqd8J+tXrlTLQ5wphnzbl+kL4QgUNwV/hmYPeOht2TSmm9NjgCVqdZys
R9zibMMciJ698FDP9SW0JpGcRe/USaPAhh6ly0+JIFKhfHAQ3wC86JKUgxvAkbD3
uEjx47wDSBAVLOXg8dbFhNHMQp0qVMBhZCxj96yT8bsDAbT3yHd2CYkVGcBAI0pA
RHttLwsioKglQwXFu3Bh5jWOm4cVPKU6SMyqkdDhkHBtyM9MafL6HmdoO7eWtMwC
EzH4aj74akbhue1PhOSOMRH2zo6Tgnp9pFoch0d6eujj/FMtIBZxt9Q+D28D4Pz/
06ztjOIj4GxV3KLur1IwiFpEfQP8fuEb/0I5pt2yFIZD/CSL9E+c61SygQWdwjna
dUpwS7L47puQSJpLwoirv5phIsa5U3Le0MO/AS/YIcZT8bDCy4YWLqAQBUBRATJT
1fujU+I+QcIrLU3CjIxfV5BBISceRDypRF/TKIaYqncxK0Z7VPQAw98ue/6t0R5T
4jlj2w+NQks2WByIDv78xV0UTQqjKedbUDF5s23joACzZHtkQ+tZ6W8jeGGTvU80
KiMYG8kUxw3ltR1IMhJPg2l2lkC/GHPpEHy9tdSvfw41mibSRJIc/7CtVjR+aLlE
wO6kE1li2gJjAInmbzVaDS9Wp5psIj3lFbluF9FjloFogQsdqPuqbT41IGX1J6lw
SX1+28DUzR6ghUEcMwMkwnusCcXz9V7/Hs0DmG895MP/ieSfoVAly4kpDUV22Yb0
XqlMjieFq8lzrgSNgcmK9pjhZm0rbqaINQQWhhLkr6Q2gv/mheRAvcmzaNzxu5ZQ
7syKYhEIiUPhq2Ejvrq9Z+UWpY6X/oAlUCW6KG1V09z1/diNNe5br3N19EMHp1N3
xHSE94Aj1G0q/8egty40yxh3+pKHiH5Ow5k8S613kmLbkcm5l7Kg82N9n7ry/bGw
iJqMydUStPUtyBLkYis5rpSFr8P7xTrVy1YYzyI/27wmbYWdg1jmCTgYuZtIN91X
D25sUpqFCE8dQcDvUy8qMCJ6QGTfJqjI0mbCz87Gcy5E4OUMUFkakld8PijUSSgx
rpNetF4hiHr9NI2Vs+e2gGskF2fYuNZjTKvVdhPUTkGUDzXm/qotZodY1uWBTvtH
9ATHKDUcfuZlzlke6jhlWsBIl7hQToHGCowDiQDXdObT+iXb7BuH0Yg+pPVQ4xA4
S+8QVTm8tuFd7TSbZeJPgnnWihwjMGPqoJHFPRVxqqgfLlWQC3SRV+MEOAnxtMj0
uBfTUEoaXUDmdpp6CprRvMGdjQGpkL9jKpI2jrsrV9V9Jqm3nsvkyiXwFn8Ub3rd
68Sjo7GPLKmWRwhPqnxCaA6YdLZ+YJoZMKylKlfBWrBVM+Uuxe4WSJzQ5zGIxzwU
R56zjuJR1mIQF7Wz/SdTfVz0ceqYTKN1ACaEOqLLAZGn59GLpavn499GSZ7s1Cfy
mLcBq8pcqAlwWXCNwswjRYM+hbMsfwRzapXPcgy0YcgEUR28SiNXfA+Qyup2h14X
TPvFcTUqJhE4mFSyvxZklyil5E+RqJbmt+LXiSUOeGMuODOt99UAZlzNIK9Je39Z
ShT/P2ynae81P6SxVTmlexsTW5vSC3UvzihA6CTkEuoHVEI0jMyzGWIDClLt2TEb
3RDCcEx/PruOxhAVvDGPb6wpzR5lEhGq451lENs+VkKF/nZxI7KzfM8Yt/TFDUxs
S1YZ8R9AzU7laJfWU+aOkdiBiDB0TroUYDDYVYe65hAQOrSX7XM87+fM0VzvlDqD
bxtg7F6vJnn6CLQJ3WTVsxM81nVhoarMux622bjENwUELIfTjAjb2ltWA148Q7IO
HFAOipNUB6qwDumAZR7A/zSZYswDNLKDtgXVKArp3Ns+r4alHVno1BuuYKADhWhJ
0pJ3SEVtHXmzBzVnFbGF2oT89/fl/+Euv8kT6JiecCem94r+QEqWCifrR2E5wHIr
USsHhffuNFtAyH7W/BF+77/tuTEYp+RBe1CHIuy9T2KsrWwzKyos83augbFzLeLJ
bWk3nGI0tQBxf2YrImwMrrXllNFy5U42njcXDzav6GJ2u80Bs0mcv4T7Bd1fNXyG
GKBO1cuGTK0t53+zVV8y7Jj2LUrYo2ZKDj5b5I3JFmbvloX8SMy4P4uKgShbC2c1
0gvn27TrE2r/gZ55iEiE0gh2RRYGtx2t4+Av7+00O/epVARDIm036gaSWysdxtjx
rtLLlImxWRSYu/5TgFB/TlRZu6sXz7o3H8i6Cutwd4/TBBQAGuIH8KS3AHSSN11S
OdrUwCaqg/VMx4RnDt3NZZE5HsIiLRQXbe8ECb4PmP26SQyArO4Cy/EMYzIttit6
8yARdi90laaXFO3ryiiL5/pIZzt9S+7aF2rVoqYFhIp8TaiXfklY3KpbcjTtQX+n
5j235GugDmx8brB7s3NNDbZl+WkvrcDMOX4zSZMaLb99EqPj+NAsL0JxlqFHUJoF
+XsjeE8sQm/5tM415IzlP7NUEtIqHnlz9Sccu0OrzyoLoyXdRSEJKuZqrY1PmIXN
EJzT6d4eFabOOzdEdcT/SaSSfb08uXRIjbHrgvZ7fKSS5ZirtCueS0vvWS9+SF8V
IkUlG/JmpXwzq3eTjNQasFGZJjcyTRmdYp89h81n2PYLtcxLFOoy7OGSOuTnDX6h
K9Tgm+erM1jNIbg1ZSpnL70Es0To9NOocpx8lnt2crMkOvBluNbqkUMGsa6o9/4Z
q8nZAGxjcDSrQ3LlpCmFrR7Gux23N8tACB+j49ZMN16mgFYhnUuBfqIUCduwYcjz
qozduF93xkHIZP2H1k7jwuVlEMojxhYRmsAlLsfkQBh2GOFmoY0wk3bbX3HUrw16
ZeB8PE6IvfXPTYRh+y3iz43E6B/NHY0vEZOjm4w8QkdcvZr0wo9tEh58GpUWMu4D
fqYHNtH3NgFLMKNgQ0DkSpxGoI66lWImiYEUmvHi1rjgzFmvGJck43jj5bVtdmZ5
g0us+9lqqwAh9Eo8LYc/VaONH0UyM8M0H3rYwrLwVxn6Egr01nrTosq54PVqqdxz
3qbKauKfBGeinCq6dFBBJRcVlDlWfPD0QNsfzkOcpH9Ae1PWJgZmIP1XbHywzIJi
BD6cI/1DDXofLhURRjRVbkiaW8vtfEyknYmFqZIjMnRF1JI+r9UpCzlC1QkWb04T
CckW7U0HjNBW/Q486nMlQFZNK171z6uGEhStcpIJaB/DJ4M2Vj795hf929PsD8Z2
pz2HSmFqEIFqN7V9/aAC5K4yeHWdURg8FWUc9Jf/0uky+YDVz5FfIiKw+ruiyu0l
ahidl+GdMpuZZuE8jifakbnbn4EAvju8L8RbPJhHjQvk7FLaDXRimOjwDkI/fQEP
GVm+Wa53B17GfaYIWdDG8yIoHUkP7PyJWbmmA07XRykxSzIMcsDA7FeDcrIZbQRA
C/09nYPQcRN79Oy/zT1ytBARtZmjTMeFwWnhATQ6cSpCqrueA0fqvc3IxS+5ogr3
AqwpqE222qE0BN5gbc3h/xqY5ezC1XIymicFmy/TeqShw+B6EPN2QdGiSJhDCp4p
9YBPex1KcVZnXtiD6FxxWs3pv2zXOz3QHMESNlz9VDPDrM4nw8lbDzOdaFfBr28q
yFVBjSYdrAT7sqc1GqWVMA9V1h1Un/PG0EZtPXaIwCYsCiTWKOaJG1zlC+TaGVpe
OsCpXD+oRBJbIlBtXXiHOo0dfwqf/jHtugX3ojGUtiE1e0a93F6ZcukNr9ZHuYHJ
yNDhTN0m8rD9q8a/o0mLCXLz76jLr6phLI7LiGBa4WZK+02mROadaed/rg/10JuW
BKwMguH1U3+g7aD7Ry7i3TOv3fbwJpF5AOwwH+6z76FI5kS38MxN4PRUl3slmW1U
YtXIe8eC6F9427yI3yYF1C5tKgccgojoJzUMPguv8VBS+2rTSAfaUaDNttaESslq
yfMapRdDOn/ZBJ+3arwgqlMFeNCsmENDhtesY+C+3rtL6ITVM2y+fWdAaeKuWrju
YMCwSlg8LB08rR0Adwjt/sT9QC1irg8Z2/hAmH2CydOln7p0hWQe88Opd9//XtQn
ZlzMyP4xAXzFa+KvtSjFvAQC9b0qTJlJdv69HlHprSayrDUj6+R8LadNWFD/FO8u
l7ZXoXP0feiJJBlxfU2+YoncFQ3QMJz5jJoLgmeDlKXH5i4KxKh6Lk6PaACA0Z2a
O1jdLivxQjsDz4XIBehNsW8Dw2DUgKQrZ7rn2QVZWvVlULbGyKJ0qa0mHfn5os+8
Ks0roOvPCi2sU1w+Gz7Z2zgA0FzGGz5JFvwO/bzlhsNYi7aO09f8ejVf4adwZ+8d
WBJalUnsQTb1SLQuQseYr2RI051lKpLgLrvAO0UQDEtG1q4gWI9Jw8zRRqqgV5RX
+d2ianHfkNS5trOVVYmIIzZzDY0SvkL/eTMO7GuQySsAigQH8HzN5q3tRpoj0WSk
nRouQP7hd3LRB4TYZ8L5Ti1+Qkxrgf4HWnFdHfhHSeNmsf73dD7LKINgxXvwYhrk
eUPbVUN9iKlIDi5b8YFOf1i7jKQNXmQqpDCIyvJKDS5roMNBg9TuqV98P7kS0oBz
Acw9QPIkbCowGLVivkganrV2KUqsEYdWv0JkXe06ReyKaryH3A/HXD1+/jBhaZv7
4nGOcRE82garMLnHcI6ZUx1m8Fq+ifgAzlPFfeWi6Ro824DevvtoQBpuFf1aARPv
sasaDYrDMsnOMwJj06FVSf5ep5n3OPVQSpDDNM7LGxOuqnJMalX9Ho3xt5EBE3rK
Fxubka4ei9Wj50sx87druPEwAYxxNoNZIac3XNXoqaXa/F4zwCZgoiyp93B9Qr7Y
vf/Q9bVzVC/b/LUN3KRxCYn/XlDpmlBlXx3gt/pFSdo0OywfBnO3b8HWMV8t3Te0
UxYPIwahRicOzbNG1CGa25hKiUwSFTH+eQ7dFRMw0t895mAMVSdm2OmOXt6JBFaD
C6EsjLpXTk+LiH0hnEVFzIbGFsai3BpqCLT/QpoToVjktVRhWIssFTdFGoJVURjT
AvJPvug7v0JubAXeHBI8m2104MlYdg5/bjBcEAe+87o1Wu6MMTjuoQpLq66+Fj1z
7/ralcCcqLSBRDNp1QKWwZKr6kUQu8pvTIlnTScobfRiXV8zUC2v+VtfZ9SWVUph
Xgmq6W3ONragbK9Etg5thmK//BDz2kSRNXneBcgFGAo5PicqIik04bIcxsQbjE9A
F53opTB4p81nYH0w30TlGomiRTreloBYENcJ8gZG07uHlLvstpGvl/1d3V60X2M+
qd+KUrtViZFavfIJPWjB3Br0Fa+rEQ9ALTdnY8vwGmn+RBHMOtTM54SR+CfFiA19
XRMQ7FlkyyG62eddJOofxmAqHVBl0dFSMd50RpYGMPyaa5zOLDrS44ApRLn7f+E0
DC6YE7lwT5wkJ4901A7v6pTWMNPAmpiUm5Qhi+7aT8UCvZBbTqL/AXnOtGPbyyJD
1qCVv+T4I8gokUoAuqX9DAg3n8q/NGVPM/FtIpBjQMu2t++3P2vqiGxqpQLKlSdz
AvYa5Cre3WBvSAnUwJjm0Mmjxe9SAOErzGiMBtwmzQTxao2J9igA8IQnT7QOPqVm
06j4NgblIGl3sNr0E1tTjkAeoprAEmVp/7sTYOAAY8GobNztlg4rnCT0TVySfYJi
Zt+yWihQeATewDAtsCa98Tny6TjUlG/6809zPr9Tz8LwCFNdYV/lbhYFdz3RdvCA
9NwwXHCNkyap04q7a3nVbzBV5XEQvZRAFuj9n7wQVyfUOAL6Qsc74mYKH2Ahx74F
OuuZUuCCQTJ+GeGI1qhwsvPAtP2nBXsZOvzKSiEX8BVDbTW/tWdEUS13XkEoBE8z
kDgYpzSmd4TxZoWQgWt0w1coscRCnwtDMd37tpvVFymO0vLetcXmnKTaNQPowtzl
Wpfb31AJApO9tXdJkR3Xigpng4u4LbCyx1pEpnTJHFhklDWjyGAOkcxvANvOxiUM
vVBUkzaveGbab4l2aa+8d8PGsD/s+QYaC/9vNS7UWnxTB0sgck8I73BkYa/rdyNj
5wsvDVVeTQqBKOS1yFTOjsC1mjhaPM6y83JAAV+hmdR47OM5YJ8/SnH56mnDiEGm
2qCzSuZASzzKox5TyybvmL6pK4R8hY+W5UwP/cQl2FVMR3EnQRFHkdZrAujzMCWm
V//uOYeEmNRpl853SwsRA50jw9hQnEKQzPHJbQcAy+DmZtPKotTmE9bgA2mKEXNH
g1quUMoqJHODNWFzcczDem6kajtIgcoA58WophYuMUQ6lxH6abfPUr8yMRkgZntb
esoQx3l+0CKTETCcHyvKDEwcwD1B96zAVNBL6tLD6fo9/e2NmWB7rQfZ/q0iyOVk
0T5S1doHSPlk0TsS/ByUwxGgKTwFEqVz6yMlFZC46K5YDp3J5YNYBpRY9P1urSJY
XDDg9sLBVVYjTVs7TqTn8m69UeMwni8AXm+smwNRNcQ7OZWbXSFlwpGxX9p2wxao
2pF2t+k9v8vW6S8S4ysxpwaUXLxV04GAfVo+b8bVYWw885p2TjYef83iowgS24Ks
FKBipc2dycO4qJ4hfMhrePjIAvgEHOVGHYHgbwrc5xOhbR2Otah5wQoef/OWXE7a
N/g0GBepcZ4cf28GWLsCvb6EaylGFlbl/9DtHMi8Q3TSAGYv7JRImNB+IPzsQ3lv
NSAR0ZF54D0vRL3gEtt9fp2Z1knqLNGhpQo25jTeeRAzLNMl7JUNRO8DWHLY4mrb
MeWoevHVVlyCfQgtTiSBkAsfFWRZTndm5vC80JIFH4q0ZWzWXZ7mQdPZzmWoZMut
FpFPYXSys8TsPW8lKm4ME7zHJXccFSybwGloBZx5iTtsk7TLBkblkKFRkpJrzw9I
rS/cgnosToyppD2TR21PehHyhX7v/AAeopju9GcnGEgXBFvBZwAIgLZ6Dpue4zV/
o3a5aIfXZ5HONhKCLenRkLGmf9q6o8nBBxuN0DrGxbz84o6ks9rqlwrJ6wIGCBgk
hqSmtkHeuA9Zw8MKHIe78mxBhDmZgUkoFnIsbNhKjt6as5B/ZvCCe4J/MKfM+BJi
2lQ7GTr+Sk49THCMPWk31TIJjFDgK35rvD7WQarcOIgFD70b8LFi2q7dOzAuCjCM
dfoqpEtf9uwhg07Kshw8xckRyK8dq8HGPz5ppxWgZ4YCglzr+dFlYWjq+PXWqLB+
mPawf9MTZ5hxu7FvgC60WJ452oYLtOVyOpNYpn13evjIvJ8rESvkRmgBup7IQZSB
vBmrTuX7anHaGcIV71TNcG20IBEVwVbaVfxi303b1pU3TEiyHUn5hKBnKEFYrylq
XvggsxwMeramAab0bmJ0Cu3ah5Bw3r5HgAcp1aJbE7Krz7Bcjz5Eymeo2lY1KHmj
jr7S3gonIH8KOnbJsJ+noZ0uDeQ3EYQC3d3zESqQDbsyX04f8UOD4EaW8aevldzm
lIAmGZgk8du9C9kf1TudnJyc8Ki2+eP2PadbUExLx2aF9pdIs64MkmX/rSBfUq4N
JGOBWogPDPnQQ171vB+8JMGIy7tD2S+jcUa0sI6bPNbR4DTaH2zMs9P3Xv2nUDN4
8E5011dBoaLxeYEQNAovM2POW7llaS7d1QNLI/pK1LP8L2G7VhaOlGE4gMJjl4ds
d4pUaAlcZjLmYOiZxIgh3bTinzBfcE1YLoFfnd5W5NSWhMx9FfUKbuzNmVgobmW4
alGgD0XUs0VtsFpY5VseGoNG9b9qpSOMDvlUNJLRyW61x3A8WF23r1DVBeT5y3LV
2sRmoIupnJx1BZPzy4LDAxs++WyszT3PbttBzJVjE+M8iq+5h5k+no/5Z/T9ab+J
Oag1uWRKna9vk/T0kQLBj4T5S8wB8CvomAotKmEJsFFVssT12Wj7Pa9BNM1k0U6t
j42pLmDDMBDQMWB4mI4NBtSGmaltKd+az4VUO7bnc3AHMTiT98sCvckCm/P4nVKs
jIsRq2cp3Dizw7KffXsjmRm9W3IllF2brTLjHzTMa/ddVMIRArBezgkUSGqCgV12
PR/8z3bBdFD3H9dri8hUslKEV11+JSwBwF/2HLcEylb9BhcNd9I9s0x/p8ppRtUv
h9nCtKCl6ppDC9t2wA7dViPUJIFQ1wvOlgklxSldGxKwRYfRPmO0D9ZIiQK3c2do
CgK9ADHqkAl100FKvi9Qh5sX8ceAMk4f/sTcf55kjDsq6SgeMFT0YFgQqZT1eYf+
8Ev0Brevv9xqC1YrdZS9tdVNlHuHlHeMo23ORkUSM7X88GcpYJVmeRt9+rf0zYla
ZBlYuErlRHE0AJEJtygqYlVoWPgtqKALLMQJAMBWxIVA9HjuOkWYu2brGpWK1nfX
3IhUH80T4icYRhjNUA+APT57h/JzXdx6+MAdymA9MlLMbazP+yDQ5chbW0NyxoLs
C5ZYiQ1f5cOKmsguCFHI4OyHLG0qPGF9OTjaLFY76SXYUrg58AW6lYNJtNWGdSMj
XT0r99Q3fFgE+6v02HhJPB4gsQKbKr7Xn/LalDP4ugOyp90bFrS1Y8TpYtGyg99g
yN7VMo6fT70EOQB6rQB8vKiUN/GYokLkiRq9t4ZIXJBAqW5euJEBqzZsUU3rlVnr
xEDCIt5U+pNKLG2Y0yIk+fR78TXqr+fSKqPW3psvV4AqGrRplPEMx6nRKti9CvnA
dycnMvFYa+AzFPjzYQDbJCM2WNb2lNfexcp7v1E2G7EBWexLmSAqK0RvZiL6RAEK
yySwLwPDvm7l4WkmvhclENxaIS3MRBu008AG7g6exMm+xMZQBkZAqMJdKULWVwnY
Lsg8Oib4xzIxBESzlsecF9YEqdHflg2IXxh1l51Gxn+QG69HlbQGCuqWjp5j1+tn
N7ub6GmBSZAchnkFICzRQeTLLQqwR7bSgI+i69ZTMeVMAw7LxZE+CLgxN1dYWpmQ
fF9h8QZOyZbcOPCpF4xNmp94FUXpXo8Rol3t0aR9It7Wgp51cWuULDVl2VM0IL17
kP/atqemTszCoFkJ6H7qIduDNZiDyqxJK76zj7SBcH6dEfh+beQy2Du2uJhhkMN6
ZfJAeZi6RMfBtBL2Fi9jXF3OmIdNnLJIASYULnL05qtMNE2kPVoHTT+mmiUjeEg0
Ka81h4zFIpWgTvyxMUygi6vq9pCMCSL7Jku7dcM+rXGPBuHgU0AavFB60eM9FB3y
k7gQOENgXcRYsVwBTzguKZb4m+/UsmAIyBfafGeXdFXMr96C4LXfA7WmHgAq+S0h
wgdxuz5ZXFfFNa7c7Y6+yohmS9Hue+0G6RAQaLBD+xeN+c4xee11jtCb3V2CHIOc
Dbzn/tf0zdzb/bI6gcpWJhnEVk77tx8F7xRTfPbj9L2qhr8JOUkroBJ2Ktj197tO
U3hqw70HNqIhbvyPtjAkG8Wkl48+DiAEpuPKmW78+7ruA4RYUqg73Oeb1gHRS3O9
pQsLPwbtsr5/oM2C0vCYYxJ/6vwT124e16wKhWUNxFHtzaB4YBcmQLhX29Gcq5UR
UYt5zD1PKJnXUJ8EK5j5R5hA7vQhBbliihTndS/EYnhFl4a+UQWnrbwt30LDKcyG
YnXxDysrxn9pREAZe0nv1pg34IqcStzKpWsA9c+/Ixvbc6/MgJvSmkgkPM5pep4G
8SeK7Pn6q/Zojih3fAao/9hCweJtBPUXdXqxxqcZk3SOkaECtXeTrDS/JGGUSt6U
nBTys8TdekokkX8Kh4IaYCPqHKFexO89L6Pwix+GFCIqXRiE/k9u7kNwSB+3VcSs
H4nh3gCF7DbeRbSC5tgHLznlmUT676ZLJeolCr9Mc3aToZ/Mcnz5IDFJjg0v7RzJ
upgjJOfc5aZTjpM8sPiGVzQEhTEZRThXxe8NjL4Qtvlqe6rANuR3m5kPft60gGME
J0F4WYXqVkKq6s+bN2tQbK4iQVg6xuOGGKqBn1QxkZpt7+O00djToUDGr19a2NuD
H59nhPRGSSNcBGOewFTt3hVXcPJrRDtfz3mMSBfsPQY7gEM+6y3SR9du2ojkMYCa
jvr+lJ4Lc4wfUMikluXfrZ2htQm2k+b3bjU2000ZnoO5J3ACe2hhixYaCRPmECPx
fJsq/v7BUFd3+uvud+bZrV8vo2Oi6ralWaoNcP0MZqUb24Liyln/HmhhEzO7CjY9
lbOwibERgByZcPvTExoJYMJaWnztnh+xA1gl9BfJpxAB/wCEId/mm7jXwBdBcSdL
SXzL4zajE37DRMJrk2NmKK9EH8u/Fq9ZVT7ae5rgFGnQTcuPjPD8DdbHrl/oSy3N
XA0Xh4rNHKuYKwFrx7uXHMLwfWZ6g+48UWSzGtdQ+qV8w3ULy9ja4KIi1X5pBZYF
ycQFmPGn3UnF20eX0jQWiiPlzUtR55ZludckZsxckPZMkSAIAJMOe8Yv5icD6Tud
Ja0NLVA6poHRnTXAavZP1/7gvvUyZBd0/XjrIFoI5cXBha9FfI6a2ffH+1C2TDAr
kV8eb2/AqIcVPfdx6Jb7BX1InvTH5MvGzHT3TyLVVTfPxXEwUicXgzhPyBoTEEFF
c+F1sQl485wiETDdY3vJGmtltBg8BVmQ+AIKqLP8KyyyryLSSuMqSR0NFctdzg4M
QhXQPBbN5mdg7+tgCXhD+NeRfUgzBA+iKvPpjaW8FIObt4/0PnadOnZWR0o7HZF/
osouirfvzfwZ5xFm4aKf8vNkoPCSqjl5o6nvMUrLCeWKa5RDc6sOS+qYicB51j6w
luY2P61dVMd3Tbbbe0lRhwshKgvn8PWkAxkWTZm4dvxWbR1QvMvCdJPzZIMotxVb
aqdOrcAm8t/9MyCKr8oylLspAnqhAvXBF1lwCf1D+3wiAWjzDcwTP9bogmtEVhXD
TD6qwQaus1rytGJrGx+KEEi9rRRc8dbyBv7XAx0sAc6yMoTRmF4YGASys4EQGpb0
53cDjPE6Kx9ULMmflj2IYZYKNYQkzB+V2uippUgm8Y62oKkR+k+yS9s4mCrT9T8i
XyMQW6tKjeWqOxbgNgtIjTtVe44wT/T3Pl5wYw0spZAzvQwU4OWav6MUH2KLlaEO
7eD7xnRN5IhQle+gxplrbcieadfrlLjSyrA7q0A5MQ2yBAwhRk3rrw2VKaF0YHut
juOmSUXoLs7zLpgIHacwEBtejpLUMNYmFMvpY6jxuDpIqlOvuIfgVOZr5GXCDx04
UabGfc06iLzJYTZJlIR7334LfY84vN8r7+kpwDuDTyau1D1XTAsX1ap67zl+qW8w
VywJelnkgLI9xpRdjoQIW9zPlF9D5UV8mtoUNhy6oUt+6Eqd63S2H0PwL2t65sIz
h8eQnWDAvvtAJ2VrXfCF9aE6X09rNMIKGZkUPS/M8ilaO6PC+ARHqXarkO93z6v3
pUDLAYG6qPdxKH1jImlRHZFz8E56VDvITvlpa8/ul9LiMCLzqLYh0aJAedSTKRPE
QDoxde+KB5ii5DvoHskossubHCO7CZzocCBkqpLMYdASRVdWrLmhzWxn4WEelepf
pxXWTkCl/0vT+oGhpys+HsNRBDKZqiZkitlqDSss94S9zT0SD0I6HTrFDGYQpUsA
Hd4QSPxNDd1Q64HDn1QqIQora7FCpT0pz7ORMn8Qg5aKXteDI42Vmum7CIq7eRrX
pkGi8lcSJEWGXRnzGZKS2Dw27ESmZ1xDTOnYDT/y5FUu4b2baO2MQ1mFAiAREURQ
nRinIAcOqrlaG8+UBSMEBFP0ifuTqJX/tdFeO7FiMKB5Kl6td6W/6edLg+r/pBVJ
oKCgWI5jNgfUf1Op3b/aIssQ998JZyBe/wqIU3ygN0eZj5Wl4qf6/GuwkNw9b+9c
EKTGXK70EZMsE/id6oPVUML1TLpSxgmxmnldoWujq8mgHltp8qGRt2SzP7+Q8SYz
x9sm3SkDN0QqFUzdzl0x1vzFxuHOMp3olJmYq58wikM7prHpRxYpuqgL27F06vKR
wxOhuQrEe+MrBEguvSKtyqAdIylY0mwdsmWONbPtMV7zpvMP4tU8wIDetH4kik4C
pZPQ3fK/s5/n7cLo8QhjTtNEXkqM6dlK7/dSek9B/g2/Igeauh9IMKB1ofCi4ZMQ
ppX2Ey6/uGP1/e8uj9+Hki41zlm8eMM3ls+uG/UNDFAD04lvW4zzqBwNKKwLpHsh
MoKjZfuBNraqCpu+UcHxSapQwf12fb7fsiPEJJPLZKvaYqNR91ZDFCFzYfqbTvL+
YJCKhfrETJO0Oyx5R1S/8d9tKO/es6u2iHcCl6zXjCwegvP8NluE5FdXbgoB1FIH
SBC351bLC9NT8qivUGx9qW8GYyIWcdzBFaBEPrDIVWRrZjvQR2G7zFKkl4ndoOKD
U4rdsqWrTzf+RGNL9PDIowxCokxkTdftw8afHInD84JTIMyQ+XkK1q9O5Xv7PTsU
gn02fWaxnBlpJJcgqA6eJzyTgvbPN0PvY1eBwlXX5HG0b3J3Szg2FA6Aq9639tBt
fxvSh0AN1pi0Hd7eopVkJJZbmEDNrT/CGUH44PS0EOKy+BoEWMvu1mjyZ8X3emxK
YFy5D2b1iC/u6ujdzYDuftYxvDwgIGu+l5wFCZ5yQncujphenSuVI8TbSFSoY+xJ
wacEUNPp53wfPuupaxuHXwYd7OdzJduee3R50JGYUAVv7mG7gWuRl4tZDJtaLQb1
Gk3+uZazXkwRth/Zxsf4wWW6sQr7zPqsek5VNLycf+izjjT17UDs2NahyikJ4fxa
ovGXDamjhyirJW8KBNGcz++W5sKo1uozPvnuYM+FR9A4dcKo/uPW/OhJjLKO3qT+
f/JSfdHhSHz+jnvRacBBS22ChR63LhhvcQe7LEReQVpH0ytpUjkjEJpkS7zlgeCZ
pPL0BIO+n0VosuGCHI7dAjOTqgWcumoPULDvLLZ7CYD92fOzZDjccB6pzdjDtbKz
1Uy3JfWbKZLbT7Q3HmEDP/EWgRUI5upbJNx/1mK63dqHznlcR+4fVNeqG/XWSFYU
y9/9o/v4r3DVecAdSev3GY4KVoy+/s6PHyZv4YjPqpZKYQYsj5+4b87HR7JWx5tX
BmhedYvKFIrP5XFjTLNIJkmqx4SldfDl9ddiz9iyO0dhZEXKEhYi8nHQZKdZNZ/S
Kopy9AXPWRHucMpYQ0lFJXEj0tQI63bpQdEytnJChKypFC7UYcNB1/TNmbVkkmQu
pwfyRZZBfVt7MsegcF+i4CC84/yxGaKhKGSTtxv3P1KeYqCtt7TrQkrXzb/3D85l
Yxsje3pPARkEPt+JFh+fgOzB1zvTolwOF+5NGZAotw0LnsGuIoG+MK47t4leYEVu
+lvIHcluPCpeJqW9CxLpQxg68khCTyjNafWfSK7TT1UOmK0bXxfYE7WLKsIY+QrF
dGzyk+uDO3ER0cyq61unGwDMOHNaKiqiS8gMzZ8VyOliA+VHvjZbdCb1BQfc6SJl
IM4xsnKvYy1c5AbJOELOOxRrWjcuydeAx6lkSZwKmJXi7MVwt70YtOC4wV/zgCJ1
7LkeKmOvpcvqQAqB5IL2Wp2SFdQ5ln+TMazYvmstCrohJz+kF1tn006oIrXxHkEO
BW/v5DNrsqraqYXK94n+mpXKIbZsqj4cuT7Atwm5R+fWzjsg5IuODyk4bE9TtVsX
r8vuoq1i3ol8Y7jtzhOnVm6PaWtBEpT+QkPCdQdri250uv/ihJRvg8DpZVaZjJYN
aFBihQtbg5o2eETngnQiyjoRRZBaq3bZkbIp9jP739nv09sV5g4o3Z07iL2uad0E
poEuT/N0m+N2B6tA6/5yC9u1GMJeFu/DUlPxw2a+LxqJzIjZHG7J7n1Qr20U4itX
Hw06L0VfozDdfxWhMAl14qktll0uTqRe9a4AMNwB7QGaNZxCLpmZqm0Lufv0T/Au
wVWZxkG0R6hHi9MQEPAz2CbIpmzZrfJXFrJImX+uhtSr2C8A9dYi+0d16Cym2P0w
rAXPuD2p92tvQfH9el3FdqYH1NOF+jNG2dQ7yMriOvsDkBGoOT/hItUtUGjvuL/d
RF9oHt9OU1DvZDoE78XcrOEBtzo7GnAOSH+tQ/PStxauSCAywXYoKb6JRMGOBNTz
jGqkyi6Bp6evrlH1wBijjIFYAQgICfgO/4icGL/D+zlbVTi0FX15zfaZepZWOZom
bWXycZuY35irRdLSfTFZeBuqofX5hJY/wVqRE89hRU4fIFOyRfsoZIpg5hFDAsmp
ick+yzlN62AcUdhaQGxykHYfsURjep0dbgbQADimbbtYkJUO8viYjRUZPfwpGDIW
0BUkIZg+AJ1Fpq+CIvdA/Y6RXCuq9O2/Jz/TAuYOEAi08WWaNpNpy8ObQ3E2VmkM
NL9/p5r2CD4EA7nhZ3L/4Br0Se7zvLlEfJ4HHmg0BvJT/212ka+bD6OpfwebkR1j
XScdRXhN75GhW1DPiWTEaocr23NSs828gdtbFN9LkH5C5D2JSoVHbYf6hyxzLfxk
je/Fo8WzlVSTTkTKIVGSxADAMj7meY/nHAk1cQQ1TSgtIiQuRIcrqOsxx322IrTZ
P18RqIVI97u0J9H8Mn3xlXY6KKb2UK1ey5Qg4HIvIrf06d0T3Bt4Zx+11/u6XH5k
VJafkv+4WhXyRpH4Y2+idUuUqb6eAO6SzS4pwxL0mQUDlTLxZGoTR7iUjS6nxedQ
bulgqdXFJ4lL4bnTmS2MU7CyzzABOT4bp/1FXgxmRW0B/zZMQc/bEMRMDMuF0rXr
nZaURhmcjrEnhsEL7T9ZU1t/GupJzmn5o4ybsxFiyLhHai/OdBhcASQ4R5oDfqMn
hiTlbeN2H6QjZivj9crlwqZ2cE+i1EPCtRk5SQRzUKmuQMOnL+vALK6PS69FAJ5d
s7ssJyorkiLOBAjPsTHKhSAiL101ypnTMU/XlQ2hUO+YuX8TP+aZ0kCa+xUL4Fpq
wnXoe9vd1H5WyHQaVfP4YVsAdXkRZxF4d82LhF2RpHgIoDzVrydBMHIb5RyAHVvc
yjcylm+oQmSgvwoHzVhs/nMHDp+hsOPHQ2jEwuK6UTskw7GqpgisatAKuJqjM2tM
is0LE5IrzCtKXVxDAv5lGrI92/cXTlcYYtewuKrg9LLd03khZcuiRFcFcoyg7u1T
u3TQ9lCez58ZO3dpDuhvzwASJW1Cr7k0CH2CeaFiL/rFguRkJe+dVvR70XXrfOAU
POHxOP6c+xkOYiJ9P3HAEibQr8UxeY9+UTwar4l/HJbKxD7ngP22abi8qUfG652n
nxW6UmhQVPYlfeEBbHQEMTCMKkUsdsOSA4XnuwMQjxfXm9CqzcAo8VDQ9EN0CXxg
E6O4T7yxL48SFYSEp9x9gX4y4sLx4IrfVcMSnJjyYvfuxLJxnOK6mykDCXU575nb
7+wE3mvxmiBCm94GjTuJxA8oVXOqdQ160cvD+srkk9oV3M9GIeR03wZdtjTIOkIS
KxKkqxjCxQFpUtZFF3EqkCxKdr10loqvl7OcC1KXZ+iWfhRWaVBiMJEimnbzof/K
pJb7j21yJclAbpPxbiDAWJpYZxfftoAwnb7MpSFH9EBsiOra8/5HU3DFw27AS6V/
7Eov9IiIEFKDjJ6KKEjZW71eUBg6OJ38aIrtktzqjjnqTnpXQW2ghYgXOZ2VaAH5
G9JlKKuCjSDlT6Ao9QucU5zxBLk2N4NqJ+yA7SKxlfmAsa6w+ITlhcHX4/80eQAo
I3Li3J8snsB6MAKQMGkO0/dvn/6S0kPHy3pY0zUVMgsYaQsOqTeXXS9q2RnWCyq7
PjnbS8E7OZiAihVidPKvHDt2mMEzedba9oF/AUs7AVjpAUDse9wdPvI76gbowFO4
JiBMr8J/xP6H1Ob3xBp2MWQ/l2KMohbqF9uDS4E2dprLn2hcm6ZnZvgVtff1b+ut
hsACPGLgRQd1ia51InO/0bBCKAiXkw6kaSeRvqScpCGT/znI4W5G+DSSEwxJd+qU
pdrB994oJ5GiKBfoQCD3BhOShz08n8TYlBHbN8OPV868ol1q8Rr2UtxA4e+DRM2R
wPhugSoF0IDCzAzmbdPsEGyl047XpoOYDgZjI0XUCYr/5XDPueJET0VsoIcIA9AB
H2qztc+ztrqvHQ9DgecZgyEtmGX6TbVZ9uveL40M2hzEClBoLB4VPo2euAXKJWNY
zcuTCLOQ06+Bqt8iq8an+tIvn8vKwfcaxPciHjQc6fyhwLenGgUI671wTXABGNC2
WVFxiZ2mlU7H9K79jAunjPCPK8EPNOPNr2UUfGfo7+YrdpZ/62cCfHCqpaG4BmbU
zrOpwdhpxGX4musirIARkVYQIV5Sogs+aIv9/oiof1C2Dmh73k/isERMqJnBIFP6
7r/R3/DC1CaRYrBhHL4iIjo/8FMrWLxhHT69YlmWjeKbO5CL9IrWudiTvN8KOigQ
PXRf2e6V1xgNtowO+qTux1mzGuLwrDL9p9pV5x286PAXu93r+MH/vFnGk5obCp9h
vsBRdkfORYiSr+JpISlhnq3X62GcH6d/8okQBkS84qiBiG2qVSt+JUqzUmPtK/Bo
pBhjbRMoTKqt3FZO1nvbuy+rbQSsy55pZZAFieTePOd7ves6rOznRnJgyeB5qISo
5iyLN9FGo8F/rOtU+KdZtyb9VZTyerBVez2Y8ReBCE8NOA3A/As6p/3xaPIbWJYA
4/0ll1Rpb0VvsvFOYfDuRTMUeFtrW0/3SRxXyf2AQ3c2Y6aGvak2Rkzi6yb71K6d
mhgcxMyy1tyQqpba9+fwWkdi4VfhzHiFRBGnIU3c7qPXGBR5bz53h6VD4WHgr9M7
p1Iu7WRzLh7yX/Tat+zKaYQR84vBJf7Uh+w5U2NtZTj1NysaAnfKS83mScTk2ZrJ
VaD3IuDIPtMm2b6sUxBwoa5XjKbMJCs53vWdxiumIL/2CNochFU93qB74YpfletA
UC51lY0/PLOz+t1U/ZU3gs1wnvLvs7OZHGmRqR8JTg30qtWqff5xho2H1fJ+Jwqi
f/9OYJeZtLtziOBPT9DmHZz2oxO1WebieGX6gjyXoKrRv88ApEWuu6y8CTbtoJmH
f8vdXdISxMm6Q7f9MWL8N/iaeFe02dGlnShOUin05xLU9IIMr26ZfJOGGg9DHCUI
5xBqRxA+gPRPhVSWM9+VCyYrnmnPLuxN2Ss/TBn44efZJvht9d8BnZK2Y2F6frn+
WCX/FRQq9c/zNkyMtFJ5MgvEtI0+30OnRMsqeLgJoXxz03oA0opN3aOSaogQzBLU
DZ1WJhr/rL1V29YCk0EOixonM4URjjS3Lc123edaMZRk0wiYXd4dwpRk1uZOtDah
BTqVpAMpAhWypAhLerhwR+9lf0PSMAvq5LLYmdkcqdY+4B6Ts+1Kf/cWlRfLZ1Hr
NsYqnL4VclozEB6eRwMYeXBSVavaIuHFXiR+wYY0f4jR0el/GW8vYnf86N5scPBE
otrKJ6Fq7bEToz9pjMbUQu6Uavn/mwGB0dgEFX78Pxmzp0JBzhbIelRV8BbDhNzY
KrxeKbDbRxib/QWCedc4O5JXIod+tyNZg/OFoph98PHIPlChaRJPIY+KqJGszj9y
MaURiQdDrmE1mTYHRykV7seopxIA8vxPNYhX/EW6VGStcVBJKw8jUytupxDyohnD
zDLuqRdaEHESPl/TpAOuv4uWV9m895Nfj3/r/rc6l9q6WVe+qM0qrtG/UUpBdgDg
qqLzi9sR/gWMliztFjE/RLKEMf6hTr310gqQHJCnHMWYk3QqihPjzlWfNVSe7Xpa
CRzfbZSmEnPRKSSO//hAH9KXYKbN/NVnW4jh/gdBTASyo+RNVZrCZRotr2SfpHMO
aqP4WiDS6mDjxSnV2A9RDTlNJAb+fmKn5o3MsLdVADlVVTQWeLc1tmo3g3F1zYyf
psR8oacn1f5Cqwn+oicuJ/R7BQkRerZLgylqX6/uWhDuzmrkp0FKnQx5qU+B1vVz
hX91G/GKly8cymxvBiU7R/zWEJWzrFb0bpiV+AN5Rm7aqFnQLw8GRZ9ajN4e9l+p
U2p0mlFfS7jeSie0Akq6NcfVI8UKILTdRxmh3NAbUNmcgD+bMKJa7zKIXdDmJRjM
jUJvzlcR4nlidOJZUk39kOSfI0S4r5LGFjsi6q9Qt5yOx3axK7GFoh04rYq/LXrP
v0haMhqWOLx9D7hs/07PZwnmPv8Ha/PIi0niwGWOFa8lSogqxqZKwR/TnUM1YTSu
N+zaDwGjyK/vL22ZUno/GXaj1D2jZ7r1lfSloigz8xjE2Y6j5pgDTwdlFSmO3bKj
LncvcGKndXAVWF/Za7vC5HFhp90BxH+cp7ts5UnrqpTkB5eSFwIASzeb2MX55yC7
8kHhJJVE8QGXPy8cNpq5mS1t6ujY8E0lR5RfAZFnxCXHmptXkY4H6XoEb7QleK7A
fHHh5/9csUMNIK+CfC7zpBUoE9rLuDW6euM23FaPPpGnzZlnl9gtTZid3V7GGxPF
EIExv+qsKHmT5fBesNQGiYKSksUV24+WKwJYrrB1E62J0GcQMQb+9FLakjpGraU2
lXQFvJimmEiYDNGgBRDr1dnkETjyvIT9iDTnLgjj/Khmq7G+W6XznkA9yOFC/pd5
5UvqiqWDU3Kazzsrk7qX7k3l0+GiUS4uwEizKDxwTVVeEMb5aRIzKf+r7K6A2IGc
HJv9LFuoompENu16iyFkZZcSdlht2e80YQxVNa2X3kT8D1I3zrfk/6EAIcvqPT7+
oPsjXWfiS86s3LOuQZbvbwUzOgfsu4Ypl/YooSpLBsNVuhbVZzNkSoHuUfL1qkSN
IZWDbHOcSeeTyjG7bzzFnYtX11Q5eaDTcA7nd7A095GLAl8HctKDufs1nR01hXJr
UlLEgX8pS2hHhQWfyxibAXqRXKkSxcBg6CbhHwddItB68LNz0ehMPC9lIWEHiiL9
B1VJwsPfGscuIH83TPPTaZ6gS3ivWdMexevtO6GeSW062u3EeptKVXo1b/zkDcrY
jN5ZWBvejbGqKS+xmUnC9POnsTiXfxDpauoZbp9Twt8+sz3a+6CTrFsubtAOSXLi
S+1I4/9LqeNwJUIddamkD8NuZYpatcytgpvezSxF00Q2szJkNT+aJehusPmVSPaS
NY6BmF1mg5pcTPqpY4OVfvessz4BmU5y/7F4k+plmDaJeb7+GRIqvpywjvoaHEpi
wr8wi1qQcIds1FsvweHcSGRWy0MRiD65/tUd6XG2SPIY/EqYWE4yxAklG0W4YOfh
Lp7m0Fxpk8BXgeL0Q3PcbNMbIlkFEnD35zoSLMjEkc2m7QpkR4iXcckQRaCtyo7e
Ywa0YjjsbTmgZuqYtQcoxRBpm1AsDx7IVg//w0MVeE/SrD4+VCWj31m7ply6A7RW
3r6bQjoG7BApX4MpPRGMT/SuoHLIhIl4RY3WTIbhjNPy0vjBh6GWKX7aLuxUJ//r
6xx2kFuATuVZ8Xj3Aeq9aEb1kemk3QyTd5bgkKo3KYiFUAxgotZame1E77BvQCM4
gWcCpWpSeMjLPOZ6/PwMjxpl25rq1toYO+UaHWIzUCaZ/+/yXJho+XwD+OGnOtMJ
PnjjcmVjW7XIx/8U8lpedywKmPqd6g1rNUI1Z2CN/DqJt96v2ulSbSulaE9Rk0sd
uOQI/BUBq9yuy9KPrDTSsocwoxE3H2qrWIuq17rGl5QhOqR6WRjX1hTl4umlUoCo
S3Q+18A9nsRmz+6FQk09UmdSF8f6iS2DA6zLk82ImY/55e984/Lj94zDmMG/gDw4
nqqUxxSD4UYr2pVa1VPE3Yn43jSlcYO+VITCirwvFrcf5zIygKQRaPCyxQy4DhbS
VzivqEGrYIvXOg+Uykg5cNRiukK3YQW0EyG1HIUYIXxq5iAFDgFr+pk+iNfiq7bo
NHQEGBI+pyTSTNsKBAJCTFzpE9ZeAYFyvSjIy5MH5gppqbfJo9wmTSfHvpvHDFU/
fiOYMohZh9A4TZGPzhLUxOP1ZKKdlz2HT3vDfAr+BIH18t1fX5arXHiDYAWNHs61
NfDXpR3jqoQkQ8+lKxVgMwKRd1OX77b90v5DRlGK9ZI7NIPVL4fGEL1t6Zl5R0bf
bS1hIGDzWWTJSAhzVVe7vk0z6Ck/20utHu5PbfV2960G46vdStiA/OH7YUKXOeUp
bMBsUMEpKPPsQABa5U69x//G1gn1/EkwX09rugcI9EcGQYyDlxreTKp46lPmHejp
sRV23YBfB7lkral0+ilcUNOSAdZ5RvhvacBIWwUfNLOlQ7gENAaWDabNBL10za8z
rNCdc+ZzcckC3OFq1yE6sZTg8ALuDqJ5+6S2Jv/d1ORoxBZeU2nccKLM0FzuP58w
Dz1F/5u79DNvl6KI0SrL2H9U94JVwz7wdmXb7Sj3/9rzlwnnombYRKi6eN1taU1Y
ZiU2joBSkHoWdVepMZs1HxRe50TL2fov/C8yFDPQIrvsqqhlzurgJRgEJv4kMwes
VeYkFsiipk9H0DcSMUEPiwD9qYraKwOocg5zjHYl/3w9ZFICb28hxdnYCEQtvf1D
a0/3w2zq9KB9hBfwwcRBQvth/TgeYbsRYMZfNfW5dbHx7ZXb9h6DDZ8Y70hGaeUF
kdtZyWlizawS1FlHMGAJc0VJ9MNnH3K42QKyztZ3gqD2GaMtEYnLQoILEjK5QA/m
dtX5Z2QdaLkuXjLcFFtP82A2ln2rxg7C7susPEk540Lluj7Y1C1P4nV9kq5hPoES
49ca30QzsYBcIGYeca3efJJzIEonYAyuMwsTIMh0UcWCLjISiCIKmCkJZY34aBIg
MU1A9vmkpptuMXCX9nSyzb6MF9rhZ5Xxezaai/MIUxCwdSJLmUsX9iAk5mKmNWyI
qKM0KtJmXDtKyqKlfR/FP0YL/7LEirrdIsTMIhg4yCkkeyD3caNDuAV78VuEfxSg
UQkwaRGcKep1B4rBk6Lwjj+pwwRdHavjqMARQdR2pZCB6YC0HEz3qGj/7UR1f/6z
K5bzQePZkfQ/9XthUPV/FOVlt4EtCfrPf3wRo8P73WBmvhbU2ZEpza6DzD+2okSv
Luz+jGiAGyUyKODzbllB0X2lSaE7WAl7Ax/i3KBxWlGltxF2tMRUYSL0hO2a34mJ
zJ/79YfoyL7ru7PYYuk7VKjZkElQvSzys8H3snQfcLghxl3gJHdYBS5GuCJtCYmu
Wn5fdVBZOs3WUuEbrLYZyszIGmGq/eTf1Z6aV2pnqmWvvf9cAtuItYrr/9+FVUPl
6s8hZ1xrfbNZ3hUNB0LY/PazuQoAtLqrkj9RD/q2vrKxztdhgEg2kGLm+ErqpWa1
VLxRKb4nAZN9E4tOtWkg/SJF4J9S/5Ds8fk7iE2PK73LsXTcOeRMl3i5IDJre0mQ
Nw6PB1g6xMS3w7fAzS319g2bNW7NkGMN7cLn4PpLTAaaDEDI7d5TQuRM23FCvZps
51ebjCXWyDgGAD8u3AKPSMiIztSkb2k3DpXPrhA/zaXpNFnBfWidBJN/WctGk3ft
8RfVVcl8E029nEhGpp8GvrHms3+Vo8boZYuf3z0D1W1cSS8JcTX/85L0GOvyAsFN
N9KVGPRIFy6qZePePLyth3tLVAs946wM25DxuyAGqrAvRtewxuOmjxNxzABflVvJ
poNRZ6xeX/FhtA1gK+5qfDQFXy6aqrIwCyogOdcDWekqfNXdDU0AwpXjsoRnP0nC
4QRPAwpmxGvqvJuYiQ7I9J8Vlk9zWiwOD+bOPJsnnZMpN5s3LBvA5WP6qtsXF+2K
AfUfUc50JuNV+UlRcZQd1Lyjxrv/se9vCeoFLZ7znSWimt+/JsK0QbD67pnpS4OC
ekY07OGv+0LDkRSSJrSw1niVGkJwwwgWYrRdonPJCar3iXL6HVcjHKUqtPdYKzSO
2QW0RMiNF7q8m/XE+DT3wVRVwZ3bJD5dusMT1QxXE1paid5P5g9DCifs2IfVgfzR
XSVkhjXG9uBV3VLWtpM9zCVjHW+BvN5UgUl/K2MEmgIFQjE216G8X+0D9sYV07oU
yOf+rq2ozNoqcgRb9nkipCHds4Hnr4bh6sZ8wvMgGyfcSL1hd7v17Rb18LKQflTd
01ft4afEQXcBss2dTZ7soKGR7lQo+NwqlM6ystUPgRl6gOiT+OfluYbm2lrtqAhX
9r4xV2hPY67x6c6sgoOqRmaEWgsXz9G9Fr00gynXwSo8l16CeFzozymXVgZMvyhR
6jMWWvMXGfoNrCH0rwgSuv0nxHoBjgemg1HWbOgPSSWOtXgEididSThQ2MV6pwM6
fDBDSji6KC8Nf2IxPdXIDwaspI/n9zvfSckhSVX5EDrlAalAikaxGH2xtSfg+P+G
iAIjZmCPh5TQOz5A3pTa95Ove0zkFtQ8tWuDtuqDwk6WmOC6TaeFR2IBUHpCs+qY
mAAt4+JYVcJcQVoFqW4w9GwKHORJySQBT9jkRuQLzvwSl6gRmuv3g6qBncszbQgR
V7HR2TA6NPn0Ye6DZmbhxBXK4vjcKeLXrh9H3J0Sgm/aEdF6FACBx7oiGSbCaRsW
HfI8CbL5m9J1QFr15QywDaWNfI8kmmJsvguAffAfz5xqr+C5wjBCrnUWgmZr9Lbm
ZWSsmtBoYpD6H4FcxMRk+V9+ZJCgaHYiTkAQbUVPYSwKEfQiy9ijaBHkW6VCovZB
vszdIwUxKmEB/DBcgtIllnbnFQok1Qhyyt3ftl/IzYDbwTX2uw5MYtDWGNH4PiDJ
lHdtOF38pzJw+eF7aHj7EeNu6Ob/VFnYGkuia5/84eeaxmF1oRnU3hgiLL8dJ0Q6
g6Ug+KIgUkX2b/Kz/QhPUCXAF7QHD9TCLU71Enpw6fOCpnFHrP/OzXvnFVUB9Aup
NG/GW6oEgYveDjUQVLMSr/keND2mIUmL/f9IeUUz1AZytlRJLVWXB87aXgQ2pVq1
ItKW2+kwEYutiMakl67ELeJ8XJ8HYez1yr4F2n/0zrQbqFF01H6oSITFVkZZCdw+
tJxxJh65W1SvTNiNnrFq4Wy0BScb/UXNi7WegZzVLy9LmbC3dXzHZY8vKxCO6O0S
t9wOupCcUG5mAgKRulszoizGrmk4sbkIru2BeWOt53EM+s0eutnq25UEqaottdFZ
1aGtLUIy/ezWcs3NKaLAi6So4l1jWgTkmpL21lYLwA5XkHA3/j+Zmrl1ar7liepr
t2V6WpQ/7dmWCQog5HthLTwt2ktFXzxHefAJxVkzI1GttD60wTkQStsxdquYLoIF
piGgVaXm+gOacdP468YhLtoWI3/uCvBqKfZ+8Qt9dhE+OBB9y8x3rI83YYntUcKf
bFDst9sSH3nbwPxqvaIXG8uLD5kGWvzguvTxzYZD92WhyJBjFHEdxZ620A85z6qK
1uFvue4IuxxvYdO4C4b9I7RtNLnEY842phH929s41MmTHE1URxuRb73rovnxBwpx
1mE3hxSJVHBScJ7Oc9kjUQyIy6JOHvKeU3Lsl4wdSn0OT2dQ7A+1Y/AZQK3m7nH5
yVIdlQZ9/+MFRFXxXMwG/bcLml/yiPlurRRSqy+jlAj1wMLfj9b3iMkVai0wm3Ie
oZoPJukrpEf4vQPk4rtCKexcUkemxhGMLSKFaTSLWEGWgR9MFw6+NJ6iyykYm5OZ
X4q0MGkq85Tlmk4wF8RtSzS8HQ/VCKC4m+mXInXmkJ5XBt2OIGed1g38cBt3xtpi
L5Rf3geO6uxRB6faiivBBtW+CD405/na/bIZR3jHHj39wHRnds+2Jti45sqBLt9z
ZzLTlJd+MQVTaBnJQfGO1fNXO6nbIu7TPZJfOoEsb88kApmV346CPMviqneEI7I0
9g7gS5fgsJJhbXw2k13a60p5c+qQaXrHF7rQ5McJqY5qsboK5NN9hKrkN5qU1rTe
tMNfg5PRXqTwG+7/qptEMPQQFfchdyeGs5iXhZyMyxrvW65ag6FQcQ4tk+8RNo85
ig4KYprH3i6cu4MZyDQTkJUxFfOX2tJSB3cag9bkP1GACIh2mA/PCJcrRu2p+NW0
HJHoSAVvGPfZya5whaxo6jc9YzgXLMjJwaazww+WfBQ9wdJhbEITiwN0/f9bqOrG
cU6no88J9bUQCQaCFtVpOdWBpULzUsAcF24J4tIRlfwNCUGN9bMSoTh1ysKm6NTc
BO2xYmcDS0t/swBou+gnDVFRe+tk15K0fd9yApE9ex6cOt96+7wLcfl1ceW5mbQ9
NaubR8vr7Wpa3ecYyicYgNPyE7RmqCE/XiETnNmlY8GMm8CxYZuASg6LFxT3d0V5
+t3HCXAx1w02CIVdAvRDcwtdNP+LuHL6v9NszsYJVlD6IuKWpsVPw+XNzV4YalUE
n9MIbMgA8thTFqkGP5uiMpjOkbYeA5bTtEj4ATlj07r0UvtRt2rsrLL0PMo7gPDN
Pi+bUyWJlN44sqDiDWpLybksa4792oNxBArZXcEF8+viabF560OxBZT5KLQIrTlp
yq/OUVe7cszCmbhlHJmPbn5aEZ3sLjgef6FAPXjIJyxkDgMzHtR1qeBPr16Qepdx
XROFZfljL95/9eBsuCNKCAtadE2IMFae3EtgiMQdWqXXqfO7piaVsm9uG/QtBatb
5R8aHLCfi9YjeSKn4qk99pPWCX22MVElMRgHEwnxN9ugpfkjrgLibrDjBMtawdKE
ZyKxgN3swBO/sAtj/145rkoD3e23nRkADoQWlaVjTXeV+zuzGGg8N4ooQGS/ACxa
xlBOK9Fe/KAieNj+Amsj1TXFhUfIBtUcVnMY3a17KMnY5LEXAaghKtXj5fCfS5DO
Ln234LZxWc8MvDbsJNDz7ToGtuTmuyAPLxZYEKDrfeD+DIWTGd1UEcx+mEcQgJM6
4wVoxhum6HaiOK/jK2gfA2+3RZ+JS95BhgojMINgJo3qhrruXrJ2uKetUrf3s9PF
8KqYjB57Gu/iTCZMd0kaYi8WcXA2Ul1+iXSEh3sY2EBzOn3v0oX2k5py9Uk8qFMh
ztjSOlc312mNU/8APRduOJIpjPD890hOVIcNsjQlLPTnqM0k9/H+LbxG0wbQW3V4
Y9g4XUKKq4FbnQyBB6sb/0UogMahvmvJB0ULe469QL7Ov5el6OQVLLbFamERczo3
FOSqeaydi167MVXK6/mpsO+SCaatGPY6mrfs7LE1hi6eK36idt96BAYzUnBUIXpI
50svI3YSHZpdGi7Y6YCWOxc4C+sg7Ai9Wu2GIQoZIRIFNPKbceUMwn/OW0BEBzmK
I+wZrR3+bdmR/oE8VWPyb10M1t5TV/G0+Isupv/RqJlDDgl6eI3g2jO2mCgaj7ka
Siq+EX/J3yDcF+P/7IPax/6GBTpdZ5qgcXcFK1IT2PNocHzXAlYyUBoopkRo6L0a
+Uc0NM14iRxClp84g2m2u5+9COJIql4g4TBjnNDpAZ9yZd400yCBoGfLW/yYRZI7
p35Z5inbKnyysOOw1ZuOnF91SiYBDDeezc0mubys0kgOTKrUvBBsZPcbQyk8G0dZ
XaFAbF5F1xF2ACPZopEwvOB4y2jM1Dzv/6UPg+1Dmhq6vZVKSYiocMuTQb40O8s5
5uH6WVKiGg8Q9qId6gXioFFHeOSFfqVDOWmG7G2W4ds/jSQdHUP+Dahp+nrBA4iC
on/7mqhjqzNpa2TmyEj5weyIJPkOk5efWxNJlfHyAmGCr3tHGE54047lL0kTmgDe
eyyMCg4cBmHiHDTrlavpIVFZbTEBF7eIq7xSnH24+UkQu4MmuRclrYhGRu5tSPv0
VNkk/cOrP8kDNE21XJdKaGptOh0vot7tIyWvekHzos6v/7fMcJH9Cv4otJkTTiya
E8UgULBY9Ow+pITsWEbL6s0Qvqa3gT+f54JDVCfh2JrgakJ28nHNmPMYyxc7aAWt
xaEXLNFJyA8ktSqPVaarUDNKaIsg0tiFGbU8zdNUWok/3gsHGVKF2QAHYMySR+fK
LTPqkMoMeMl7Xox3k3siiTW1omG6KxWLTPSZHDBaXD+NhMpqu0tYd0Ept5kbtAmx
elPyiJj/zFDB+/svU2dWxc3DkZCeZ9GDHXaSecmoYMXh2MUkGVZExYQZVdZO1qj/
tmhGGU1/ZQwGkpsL6tTsyzSg5amZWRE6qmf2Xm8UQV4L1+SixNYz+eZ8QvVvNjTO
imVPYJl6ZjDKclfpJfmvTQSIkbcU0WJCmN1f4W4TNbiMsolgzrqovee3iYB4DLiN
XBZdwg1D0Tv1BCdOvBKgileIGQbjWZ6kmgYdbEMjjPbqU/nDOQaBDHOZE/o/hbqp
Sg10yfdyUiuMPhzDAbyclWxNBQRFfuCSTl+SV6itVQL6K5+pq+9FjUqQszv4KlY5
Qbsp7mBOTMeSYPIsOesgfH6xnQZ+7FiME3ZIyVQq9dvgZxF+Q/cuvsu74ZLyh41C
p40/Tnb29Ge1MEwbBP+5jtGycolBGtzykgAOSJDXIzDXOnGja/uBuIXSwYfWnhiE
3+HK+D1MENow9iuWG6nMrtxc6FE7K6qUaNJLGhEeGMCfFHALcLkvOOsmlzZka4mG
GcjqpKS7spxdMMmAwpbWo0QCi6SmJ3nByQdSLt7PDxsnPJaAROlK4oRoSTnPTiI0
lok/zkV6Dd2qidxuMCoOymT/z0x3KOOnICyw+h+9Qbt6+/uX06FLbK3fuqGhc+6W
7zKtklnRFHJ5PqpVxpuyiuGdqo3SYURsgaoH62jlAuSM2vigPGy8MsroPt30NKz4
ND0J/EPpqSpihXXuT/8pXJU7V29jpEARC4vVPi5OHGy1KcT6YUSMUOSwbIRseCPt
Lkfaq2kf4Ihl2eY4gPVS80Iy0X5fWpvemJqm7p41FP0PuQxTbn9z75Q04D2pnqKg
KJvlARWnMfHo6kDm/iVUcnpdJC1CHnjSMtX75nqpEDN5/8mdhnJGa2KAg8G0qOpj
z4F+oKVQX38OiKqhRYF9ci4O5MO5I2ekyippFuBjZLZQU5xy/h2zSHNcJ3GDH4PT
vTiT12Z9Jk7TFMADoI1gbdZdC0ATCLaDs83KSfppmdht6pEYnVATFufkA0AmOaf9
YVDKTVK27J3Xya1dZHyalTBX2sI67MrhA7efekeXXEz6sal7LVmwPSZDCAMlmuX6
bh3zkjh0Ssyo2S8wU7u9e46EwjbVl4MdFx4+bf50nKXkpP1qRT3jX9inrfQpUDaj
dPCeNKmM0sNAnRm6P4j0TThCRexs2W1nUGz4U0COPROF+XJEsD3gFUFezr27BKSG
gAERWgQISbRZyjdDb+LvvuIU/uJooBQGfYrvRT6L0GM/NJEBdd3Ke2/S1IOiqWkD
i58KBu5yyo/UfqPiz8ArTrH9VTASUsUIzEgemCPe557LM7HxnqBvmsNVx+uNdjSS
LOitDNaerWqqfJ9tZiVn9CWEy6e+hu/8UHS0nektgtKnmjNC9v2T4sYuJQodTp3b
/DPa35DYJbv+ShxmrOorUY8QpqfBVeSB1AqVda88wCU7f+cM7MofkC+JNSH6/j8o
tUZzFg0o7nygWaiaHjl4iPVablWg595D63Cg+S+MMqQEGEZMXQUAuozXZvPZFRgz
NjhSbCB4OEHWCG4PKRpHQwL+doJ7klKWQuUnKl+/wwxbDhCjwQ9PQXkEHfTJzJj5
VCJQIGqyrxRWSldPQ1DosOZp3VmDMcvhHo+7WhFFrUrcudfIOcUeO/kevs/ZJdYz
pwkaGdL+v7EyEV9z2d63OPWQW0KaxoX35fLgm4JW0akxxOUZnJhzpDVpXEh3Douu
G57K1ipSjeufnzBYolOXvlRh5pv9Lb81T67sKQUTEC7ZLrYVMgeMcH/kcX4lwWnv
uuCRu3oX2ziScbsRll1/rSatuo4OhUnRsWJIhD3rDntPYJsBXhRNqsV2+/DxVw6b
BzEvxcHsSHyTbBzyhW36o3CJU2Aqn9jprr7NYIPEOpEwR7XnnzF7s6H82Ky1HaoR
wf9mgoI6vXnlzyitJQTotYmP/Af4WrFzCUTek1fmcuF3pPIQIC0ZEaMbxdT0atSl
k7hka6/iOeikwEmLaGHkwqnGUMAd4tamhn62LiSyBYU0eKHbizsw634TJAC+YyvS
bs+E9BwWoV2In+8s9shPUvqATxh3YS9yckIsQq6OZgbVZv6uGeq0zDl9glcKCApN
1h4tsAEpizgEQuuPiDujN4oD/GrWAA9CgQn5Z7wd+d3nbfQ93GR0wCDI0f52X8rb
YwXMqnM+LaMT388w6C97Pi1jVmOQwdHK8CMTt30vFS48A1TKxRCRzVwnAqdPN/sO
XsoK567CAy6nLas5QvA7tEbSMoSfs5u5FdopffeMih58eayjWhI/z9dcV7D1GEXf
tu2Zl6Qr3HkILrwmYMJWXuh+TWe4H4UgG1FqhrHCTncRdM3mumgikK4mFiLX2RQc
j5dwRkgi8Z7Q4eb9tod0+jfHdDWXG+7/pvlnWsJuE+tW96mElpvpY7kelJk2gGD/
isfHOTK/sk7cED/bJfsLEVG69qQ7TZRDIwynCGytMk67lKukvRSkdn3+i2gNxFl8
oNdbYIg4vco5NKgyAZM4CHMEJED9/kMrZSYxFajJqYGj0JRzh7z5Guw7jcpJCmAJ
1cuEZcsK8aEJM4551zTs4N7o36gl4gJ2mk2T0UinIxCojzz/ys6RBAgfmauirrpm
zYg1aWNtWMUElScBZhsqk7hLSKOrLZOTjm0olyT4Kccl8n0Sba3hqivRkIJzv8ZV
2CW2nPoPGrm4ABWl+BsiCn4dNqAV2YOZUAr9sWT978Kkls3SEyNfkjswLW+Li1dI
1oQnEN4swJp5sr4cYacdLk48MFzBxrQdRyxLZRqnS/vlp46if771V1wa9E748lfI
fpMXnnZXUk626yVia1fZ7KE7ixT7r6Ffk31s/T5XviitaY65v3EFCGG3tZ+S9Uvd
krAD1ZCXlyg9SFIpfTO6AgUJ9CbaA/xkfj+dPdcjxpZg/vP0UMJZim3a+TEFGh7+
12EYB+TLulQ15u4j2/pyAdbDG7im7mIwXpzlkAUCgqH/uMJHSvNBRtUqVbKkePwB
Os+2nD0yhi+c2Bjhgvz8jiZ6iPh053v0J1Z1tsJOB5VPYggiBrTHZ5MnSq3oRhA9
GTwb8xl9Q3W0h/PAZm+ulwy50CuYobAcnogHLE4ehHOMgKTfklY47pCU0Lg/2/zi
JRSDNa89HzasBLrBED65zYvmgAHM/fbGGWOle0rIKyL4rAdgHc1edzflfK470oxS
tcOKGp/Dc64WMLIZWRQACoC3RqGzM1GUuccjC3AhzdmkVVnldp3tVKVg9h3n9Gml
Qq1B6ZkGsS6FlGYx9fdNK6OqIbrShzs43Ll0tqa2QwrPSmcocbYpkl/hgRDAKLO/
o1K4vl95S03TY3wPrYvhVV4Utxc26sF+M9oQ9BGRn/wbU5aG0Ohhcnv1r4He0sH7
Xzg3BPANfL7oZFZe1MdoqAqJsvVPnmc7cXhAbD7+UZfYbZXFjJBmpJSrDg46BH9I
c+6ZTgaLIs8PvZstVo5UShjQy7uOgkpkIVs3ZY6Hl3oyLB/kb5wmAt7tf+Cd0H0W
vjRCbHaK/tZrAutWvzqTXxMBD42D/s+0bq4xxWciQreF5KgadbZ4kr6C1H7/lxT5
CIbiYCTk65uhhBzEL3yYwC2kJ0v4ZA27CNnixqiewhQ5K2A8dtHp8yaI/sj+rj5B
xB1EX3mjIrc86IVF8CxNwMliodNC4o1AyiDs2WoPiKwfOUOoEWKr8YQu2ghjVKls
aLNWQ/xhwi8mEiKWUPW4J0MtLzSjzt86HKZLyi5zeXfG5LyG/zDtnc3AQFLJS8hd
jZ9iFOnoYolTT0KiUwzPepSjnQ06oTS/I5SNDrv50JSqzn9uxyZLPoBpPdAn2m1z
x7fK29kPkuH7F7rL8HeAlOydmxLlIHnMX3W1kVBZMcOg+fO/RRR04hUFIoOMWVPt
jiD10IkJ1bqJ5jCk9SLPMdpwfw6dyogLG2Cdk7CpPxDaNtwC9o9RDwQj6HqoqZSY
7XABHe0sV2ifRwJxKseEHj2t5qDF0PpSibWoInCDJmD8uJ2NhjgVgQmUHgMRSMX3
zIgUM7j6/Echf/mdOWRv484u4KhGPsAJkE51kkC+ZJCk1ZjDEYhUT4Y0h6bUMcNK
GZS+NMIFUYFOhCVy7wnFXBSrIg+3S4YlisC8Y1bBjU9VReCD0hIiTQhdViqQA188
gLrZATA86vF29B9p7MF6XCPB0mhMaOx9qASuQ6EAxMC2bOhWoJepxm84kxHSIwKg
gWcWpNeg7cD7txTFdNkPK4nGIsDw88y+e+OoPzs+HJcrBTQNYIYE11JTWvcrlVaM
z87PImkurV/At5b4V0vE+BFcK0olJygVv+VcWyiGG5Y0SeLMLwlGZHeQJE4B3G//
umSzWwx1YewpfVxYVfVpA/wvi6GMxCj9ZN97BLRbuxKur7fSg4PeX5FhGbPy+pCS
DBuELN8EIef0/EeF6ArDzxYsM8onUdja2fZk6cRFr/HvRdUwZe4KadaHhaBECfEU
iwD6bHLdbk9x9Zs1GbiXX0rOW3egDPBhUsj7vbR4pYW8LgNpo4HWSrRoQcX415fZ
RmMHX7oDdx/z3C+atfB5VQH1hmnobH/INWnUR3yqKnZbM4AsCz6EzzD942iZNNyg
BE/+7P/IqzBKiyhgMipnVtUK9GcH7rug/AuZ5l5Dp5AVIe7or3IdoI1tVbEI9I4N
e15nvEu8aCTH+PgQqO5GInHGhAV4dmt8xZ/RTpA0c6wrSJaX9j7WPnvAk9q6Mo4h
QPLzAUsRimMh1iufeFHgtM6JZl/eN98Oy9CyaQIgV7BdLmfwwcj9VVMRiK/IIn7F
FBjLc1QReuiLPDteGTbduZqmu0Fh2j2ocab3Jb56oPRCtsk/F7+fAZ4a6SLdgcll
8TJow19REiLlQyr8SRfoDiahSabgsVKER3VCN6HmCDNWMZTiRG+8VIEbfGXRNtbx
lsTurDHjPWJFWHiAP9dSDrDVzaScA7VfIpVdvf/HGxRo08W4vTtpAAblg2JibFvf
PKMIxTDf4dYKfs6WpSTJrejHQRziDZ3Blq6tpYzrwXEExUdyNEftn8OBBBro7b1x
mDow9jVp8tL7Au70faBb0GEforwMh1HCf+fxlTCcUaSEhrR184gLpTK84qDVfj1b
7d2cLYZ0PgmHB9SUTzsj4PLgF06Zts4HasrTwGqCchXbatuiAOs5Yh7ThqZVYgFN
xRfHuu5zoyE046iASEOV7+DwEGQQjBb0UeNFXT9KSrig7RG0Q/Z0PtAnCMza+Unw
j9q3CfdedB8fROO2+klXeeCNDYMVqmYvpPCPbZLgSAWDZxB2JloT9AjHJ3or7e/U
DIOBBsxkHYzPv0mj5czAWYfAmYflQiv9juU+DDC/mJ6Ewz9wObxgIPiy6ICbbG/W
yE9zv+s61RNA7lVz+bL+hJSsr9iHMVqQLD747nw5WXXpBzsadczIALmey1iquhSL
j/A9YoTMhGwMwh7X33IzaFCfPvPzZhQ1kiKLABGhiD7W2/iLueplSzD00zB5k1JO
4kNvRGzxMJZIZOq7Vf1OXcYJOPyAR6S9rak7ib8f0Xp52yiOR9K67rowtLkHXUII
qsJXKbUy0bIF+HLceHljUyZgGnBepNxWopx1KptxyDKyEOqTlmMcP5urAOc/eRcN
PiGf6T7WkpvtXb5suBNb+f+fT47GtyWWzyUsCeie0VrBpwq9X1Nov1WYa6Yswqgj
bnBe+JciAYEFfgpiwAXre6Mtm2A3aW6B1cXhk8qF+2ldQXRYohb3V6Db/IvWc0Wq
2Rvmh6JdDEUoOdrIyaCMCB5c1i0C2YNVX3ubRaBUjTQ2VxwClHQuyJu5yvfnyiu3
UHrNGpINEOSHpW0lUoImmkYyYrt5BScg4L9FpJqQm8ZGft0yNK1tpeanL1iBUmvh
y10QDYNgvbVHIz4JEqN0jkgGRY+wWGAphzG7Hj5njp+GrqfgNf8tPqKTgr02SwIw
g41NgTu0K/Yc1NQFnnmN7b4vFc8a97FPCsUz9gqXplpRElVL3oQFVrrbds3kzNaY
NLzyqJWvETr0jyFSKPYuygkezKnPIA0GfW7pA6ZUk/T3NUVRkVHuiS6XOqUkxRov
PFG89K0gsOZOV00bcyPPKTgEH+43p7vmZNrNRXMqwfXqWGdb31exl/LnUBl99Mk1
KTwyXEzO0t39a2rkVvLHVcAC36xaswdTNgHB/FbipUPaz7BRKjR2EztP3rX7DTIM
KwzsaQaVcpE9hqj4qgIScXCYU9z9GYAIRy65HeCpmar9BdG47LlA9Kndb8lypQwO
cIBSRrbNg0Mic7SBN9+tsyCkJn4P7kD3Z5RJob1y3C08WZT5x2Q83CHqJ1f5jIGl
lX09emiJua838WIi56gGzSouMzRAKFx+ulbwe7Ru9WPpcHr3j7gdUulHz3fCOlGK
c/teov9Q4j/c4lJm73l//RimqbZw1sch/1VKKgY+sCFLD30dPC+/st6BtdwTYRWV
jA0MzJHgULJwtbumK/xW7KmyYd1unJkP3lozhJcThi9zHro4N3pg+j2cVPdOPan6
hDY2iH7UaSTVsAjzhBYg8/+161ZgtEi28rosXn7I7gEMgxBAY6UGtyTSlDUGmFBW
9sWwJ+WY1Q+RMG8OKWZ2GZ25jCPXSREU2KWV5xu3DKALmsVRpUhzJeQQHrwsI4Ef
/NpBKQbdpOG6b01G3ueoaE8zNj8LEZVePvSdsgJqjsmM229qnsOCvJkEX4Ki4FbT
hIYSeJa64YKrFFisNYnMHMSHspinaP/HptPzUDLxq+nVgtW/0MmZHMkIEhYsDtaq
va2/UQlXsgcGA7KfkARaxHzowVgHtx7uAOIU0BHnREjENX585glB0Lfm7Ck1vHZ1
K1j+3X9mGTgOVZqMk8H9dm0CHqbP3ea9LlV6PkroLBuzjnKhfwrdjzqe26FbCQk7
m+j4m+xjKMTl79lWGdVP+reWWCSgAuQixCLd1izOeMcv4BUj1wB4i4MlEIWxtuyY
JU67aGGt6gK5ZLoYaF1mQvIy7Th8Xvlw69lqJ5TKpeBLa2ChQdifciGZfA7y2E55
ampqlLoyvKS37cnATNm4XXeAD5HayjP5I7nAh0zHumT5cz+HIRIspkhm+4fhIh3x
e6LeBPwt45uPOcLpA3gCnd97HR9Fdd6fIzIs/+OWgVh98XZS+b1/5GVYn6DZ8Un4
/Coyr4EWXIhr8Iotz/JHLPOkRkV64mz9kM7E7yhqM4pLW2spt667DC/ERRcB3gAS
i1eQdyXbSk5RXxiRap3mgpmrDgOA/a+ksndYpqute9vLnd7W/w2kAioPRRB55XsG
cjAtM6G1XT3A9vIxFPAOQnPpBaJu/NsWxLqG9I2RUGryi2cWHbZC3X/d3xd99cxR
tYusRJayQD5KrfI6BgVsEXCL4J5fM0qChAUKMssXCZR7yC/gQSiBH4/mQhnlYMkg
AMt0t187pSrvHqTN1nxvOnECsM8s4vkvk8c7ynyEHfLwMeN7o1CFFx7eGp2ybRSX
knAVM5/3Rtl6nN1Sjol0ipPhBOVsjEJgNmGWJpfrHfaz9mGVv8Adga+OZD/LGsfb
acz37eCISLnDosdwxcBLAupRWQ5997S0ZBRVISLRyl8Ye9fRYCxb0glLsUUUL8Up
wLdceIYEXAqmpKVZ4drrjAd/1KFn20PFPlGBFxb1pnx+ILnmr9HL3sc7/yZS1Bpo
ju+/HYg3vEtkVjUmbCcANGC5uaSeIwFGESHuJiqgtcKzNb4k0Cci2BPMSt0xQNR/
ctokhgRlrrpV1fWYngxj6bt6D1TYCgvsdhKyfXtqBmXftnTqhQfqTZRB2PBXmpQb
gnCPUMN7K3jNug2jJbv81kFQzo8hJd1zSFSfLt4FWobNu3k3prbV9UA6Et5rlefe
KxTF/aQ1TViutpbtIRnUkJsS9/ep/2PW79qp+KFkYOQ5PVsau47U0IToZZjcs/G5
tpaJ+vvvykwrkSJbBesrZoJFZJcIoSX+Tt3RFi2WKa37JJS7vcfWq6nt7qH1/0WN
1NSs+r8HaZ1PEyeBPpnM9TPyR42j+SyWcF9S6TnZvx92GNZE7w2bw63nIuFP0Xb4
U4Ob2WcAaKbZBxIRGRiPM5xflvHSeVWVOSTpv8O++8TmjfI26czVzdZPTM1ydz0t
hKcufDXyVhhwY87255U7TXvSrqg6Yr0llBbjGJvd9WjebcPhQUiQOyUlwwjnQUeL
oTyk70EAUFXh1bdsK3jcVJyQ8hIcBbKF5OvWtFqik/sNMFDB01gu2n1Mnxn49oxV
SDPcBB3+7u+O9vxq2IkrFJE7N1cx1LFEigGMxbCbF/9EzkS9+lvYJhIbpY59USqE
fL8voSYOV/Ohzg+VqJhPEbdItChik1hbdZGymYWMDqHhqDjpkNfKN1dZzmcnOhjQ
TP3Wdyf+1ca9aM7lLDIZPYd6xD3vCrH8De9BntZ/7KZmSDMNzRRsMgGpJE59IqhD
aYkcBEXIFRMsxL6JyS5EHyCRYHRZRFz3juCddx2e1PIv7kwfObZbFwlLhJcEISK2
kQiBNGgFuf0RS1a7Y7H15ChpdwR/gwjCKCZKs9miNZpdWLz6L9vuGP4TSRauzAkj
yplARrbPvOQXwJ0xdWdR2ZJwDcpyV/Mw0HwAcZ6QzA1hxH7anBeQ865MNZ0xlJh9
xvP3xbfqVv35HLzj8B21bLMiFj/XxkXS7KtEpadHDtGaHmKu7t5lnbM8qKCXXh7W
PgKdr8ssiOReJTg4QYmN2tdoVK01/E8PDK340Rj1RagcDfPVTmm+XAXZxbfixXw/
VJF7cvIHk1vSPZRcQM4ey4K5NGoiLDsW0LO2F/3OtIswo6dbAq83f8TRNvtro71x
HDTMBQ9X0ZGilgKGKLhlej9mU9+CcC9Oh4Opom6l78/f4ubwSLgP7X2P0E4/D+Ox
aWfuU8wS10zndq2dHOJ02MDxQwwR9KzAvdq3qYGpQ3bpD/83uPB6gvJuuZt4bKHL
WFgphdv4DLKf8smD/OK0qzs4SpO/xeTkAQrF362BFUAxdB+oME6x+BFgoDeu6z5a
+9nyDqu9fTqeDfBAaYCsyp71fNPO2zETOsGynu6ssRaE3wzd8g3+FAByH0vTiruG
7YoH6AoOyS6PfOFizhlwZ/pyPx2sBYJlAWj8ROVhwHu5k81nRaQyM+GmtCv5Qqat
kz7CV8C56JkTI0yIPlpH7s5g0g7aZXdBl5ywucwlUksf3xGcJUyM2zLz3t8wyrum
WPHPfYAVXgCNbebp2yIbtQ5WRRCbljKTMwle1AI8hCI1RxcXp/rJbioXEMS6SfZt
j8P4zfkxNOAMr2mE0lglk5IllNJWgyh6iJcKOvxv9PzG6YccOgcMudCXhtAH2rII
szt5WcYSp+sap80j01yRQbo9qRBBJUq4XKrDlclGl8iiADTLASUZvjIAAH0051Uw
lPhrz5RzU4wyn+uWnrmEc3ZAtuFbfyy7y+rDJEVyeTmQSQFubZrRnnsRKaobnGOm
TJhZ8PIzsb89+78at7IOXcFfCCqCm7UOApmYkiAqjVmHtFagbKEE+ID3t/lFvWm2
YlAOg2ngtXl8GAfRTYg0iTWD0XZZMuQlEFZVBj5Ak8x06BUzKheh7M0P/A6NbiVf
ccH5pQLCwRX2RoDYBa1X79osHCoiVn4rSaaITcuexSmiTg083k/XopJ2pvXmoluA
9/zBymWOL54DIV3Gr9niU545SlofsXfaR/HLtWvZ89BXrQDPWZGcqfKDXs672BQz
ObrDr2OPJSAsCxj6nSw785632aLjs1Nb34ew9VsM43Fj+0PnYS1NyvGXdbh0AU1I
iK/AMzsqf/EWXOMhuPW28CbcJQUp2jHIY+bVsAQaibOCyYUwuaPQRLAhhU+79WQx
ksSHF27pxexfiqWskiCnRUcyhWd4jrxVmdFJZNmFIc5P+301bHVdh+Bc0sGoqe/M
TfJRxSv+MPtClhxSkLfKg4RwrD59BWBW/EqWYcxgPSc/hTV0eg2A7GL4QshXgOvM
RQRPm0/RQLIIbUs5LHJfJEr9bmOeTyM5nghyhZulHVMIDziIJtd6fjokn7C4gW6u
Icr+wf9vRNbmjOsyBfuDSxCS3hFYbNfVuDFfBQGPJJLUMTpL485jha2tQr44FeOr
xlCgLJsIBrJZClwxUFo6zTlAaJSDpmwnrlc4Bt81dlfztEqANuILgpGdILerWRpB
eQD8sQkccQytCUqG4XABEr+gpkynM34JrDQmgFYhp0WPD+cT441FqGuqtz0ncb5E
lqKmVlJfTRa9oTHQm2wrUHnOmCCHIF9da9J+jfsrlAkh3RYBtDsqHQuA2xY8DryY
UWpfoEVzvDwN2BSGSiJXVStBkhfHv0oAKVJZw+BBEVbEQ9xYu+E6PhyI494BgrHk
IslD9hP8gkBatH2OTdEalc6jg+9cmN4Mu97oLorXHwK08doDze7NLwJXm+TN1ZJU
c/DgBPoUCGFOUc7khGl7sGp7JJnF6tPkiDDKb0CDdkdbTlZYh832i/SQbiTdPWBO
BKQIJr/gBibqCKk8IHltFFPgC8isWN40KrfrZjfuHoKPnwrIOk4d5IMxqlqVLsF8
o/y5chKH+gNr++E6fa60o1cV8ayqB98u1ktHi2HCDSvg8tFwvVYFIEfW9jXZKq6b
qo1GQYNIpsaRmrW6dhdf7RNxDE5NwLjw6CTn98Y3zC+MFtqcojDR+pkpzKoWr0jh
H/kTqveHjESdzzY7RR8BRdO80bKtKqUa8FAIfhPfmvBns3QaLRmveShZB81wqrXs
hJvV8gAbe7gdoXAh9aKLCyPYDjgpir5gnJE387v+XZuBr0WxRTQ7yuLJJmHRDyds
1crNMfkjZTuh3e9t10z19UtLbZYreTmo7yYROiuO9J3UcLTA94tqetX+qo68rapc
aB/4w5yKL2li2YuepoFOX5mpB9LdtG3Zayauu3cUo9dILWzMm4RcpYXoWimdvNG2
AB0ByKFFadb5i1NJ8xN4D6Z4xfvUeBw/f7GLeeyzabuIIjcrkmXvBi94mZhzL9JI
rwuOledkOSCrNRmh82Qi7/l82PNFsetJptx/cK+v03p2v7i4/CoXVRPRynM3yZf/
iNm3qKqwbG64hXeRkMcMUa+JZe7jcWRKj4rhx4dqbHWebFI2bD539fHYmaBkYcE0
VmPPoYV2Qg8tdllZnjIKEROx6LdaWvHpVjX23dLDuLOCxMdwshhIQolTkUnU6Bo4
aSEE5EkaqwwGY48F6X55Ha4mlCMARlvZxtAy1GS1okYmCAIFQ45z2qtKK+r7F7dU
dbPqAYzex4YtFWu5cjXZSBfv01csoOwuCBzttOmfDexPLMyCYsZUk/iOf8lyFzkY
V14uR82hMAYff5tei4sFLf9e4HACmI0zhFsTqxAYEC/FX3ADZMsQVU1gOO2Pl7b7
d5MQWRkxslMQVn3n9H1b1oQ87pqYpfYaS74b/jXABSNMgcDylTvbWJ5Q6Q5AsYMD
WKKJWWOJF/7SpMa8qC91YYXOLYBAJJQ2+S/qUVj0hOIF4VYHzk/Jm94ZX7QyIKZy
HaCQP3602YMWdB87DVlTaER4kXtLrHVbbkbMORC6ehme0HXSpEZxHhoW1yxRv/Je
Xvz5OvCO0nt8dHjJKJ7vI9G+dzae5l6BAl00V3C/j4RiFs0iTE+lTaOwp1h03cS9
GcjyH4E4mhiWhxXG4PCuswSP4HDVrs40p2EvhdVolQ2nWAucvePKsfg8tYuChosx
df5JFTJ6t+BQKy2bixNGwSGEax3dmJG1K5JjuaMmb6gh45ryp8UICJhjPXbFcC2V
CpWu6FQlyWgX7fk9IYFZ6d46UkRTFXgFAEVfphqG32yni/w4F/EGrycDpS3Ys2gb
sapcVH9KzcXhqZMbpMg+/xRSxEbLbVEG4rTtUo17L5r3JvBGkrBx3yA3T1AYmGsX
KsKEo3eK1mwd/O9sa9eKC4SP/jwZ2mDD54eUp5sqVJELu01ep1G/PFbgJUh0BxjV
ZvDPitHkc/bu5Nl0UbgaZa23N4TBx4Ql9GTW2utN+6VXc60n/DKXxWE0o3Os+nJc
o7dEUs3fSBNfKfm5vCpzwtIvePjBEF/UsupU1Pmp5g0K2kInf16hRlkgqJs1Xd/O
jaZ/sYk08KVJIyCNh06/p598UG62zSsuOXOlSwu7WWIzdaqqG7+8C4cfEU7R1GuB
5u+RO64N8RHm6s4y+dVa7E3FU12jtPoPcO4gs34TM4Yk2+/8VhO66p1bpJTA7SGw
Dsf0smasmB08Fv1SzwruipcLQ1pNkVdbYAwlL3d+LUYgGH5BZ4kgE3fmVoOTX6XE
DAbf9tAYph0tiUa5mAv19/876oTZVhnnOW+XCjxNWajmlj35EneLWSNFxhrawKzK
ZJyROz0DON8VtLgRBmoTEOKWRbe00X5n9rwFkI69JJzgs8rvt0E2j3zPKVZF4OdW
JJoF43k7KlmxTKeDnHqKM4X8FiRBYX8eZ54QcbMcRtPzmLTfPSy38BXT421SAt6m
EZHGT3RTpDUrTBjpM2vYPa+ncnQdOMYLT6EgvytwcuYrWVq8zgjNQJumxdqb7Yyn
GVIUSEeOCQCvm0tFrGR/miGcpEAO4loaOE94RpnTwcNca1fTW4MC8pDE1scNJkv7
3rmsdPYVvzUtroYriAHbssXpLKHodAvmnGT67WN3S/gYjWheG/4hQZx2e4DqfRLM
VIhupo3fgT6cv2NPlClNtHkJCdhRStwPZzj3p8oZHlSDcvSsXVP7vqoTnDVgkvhj
pOhmOO9KvdYKu1lYGAuE2SGnbwRdGVzWIVpa5SPbrc2Vs3RNRVScGj00hLxtbKAW
HPQBH4tOa7VDcsoofgnJRWHGicEVJxuB8Oj7L8UynJryMERKuLFctGdsbGZktoqi
/h1J+eOZP+8TYzevKJq5QuaqtA2UEaobc9CqkGBy+8oaE8c2pj+tg0z5GCYGOIWP
VsEySQ6OfhAYhzQkdBhfIJyyfjF0W9j1+ueH6PvyKysShOnKSqiBxoAi7c6sFfOX
IuPuam1U9vNCR58nCDRQaaSUEw/PyLGUEevyoTHyRYlUEISZEarT9akNVBt/hz5+
jExZ2Yn/6QT+OFgpiNwCDaKiWyGuT9+Erhs3aGt1KLdYEz6eAqsf+cJdYo6qwSjm
9y6c/6zXCOFYTSKZLD/eqqEiW/JIkt4GqrHaF2tM2uNLYwVc8EpPX7jrXmfulPkF
hZAzvzHyitO80LCUxw6zS3ev+BSR2VeM5l2Ks34VFKIyzqXcFeNBBrTq709TkyZx
fwLVc+jTgGoOWRQIMhS0ph4SiTu6JXngKTCPEzgjW55RbIb9X5gnCZTFsnNxkRbp
ZdEz78FN1+fu8K5H7tIyjouyhpo6ZxgE3tOMFG1Yr+A1abEBv2BV2Et3uURc5nbO
/FQ616MkiuJHl+vTIQmYXSR/yhmOpG/OBXzSOMRG7n1xnYV5pUuNiXKKRRBSZiHa
qHulYqN9vvzMign8iYPGQIDjOvUKsip6YtUaLxk3Kkq+QIC2wYN9W9U33Q5eAcuj
E30Y+eCYU8SPNTTBHzi8zNRHKu4a6Pk5OSsyugNQBSenKkAUdG5Rn9GRrO5Ua24f
/gB6h+5ECnsVfEttukkMW0mB/SdwVvRXweUqTeDa2/ZpTnPLV0+5k2Vc32lmHPSe
SSCAj2RyI8j1rnQMrIVqqGLuzghKTi44m4TLHvEh6gaQd1YwNbVdslLw8fAnQmU4
vYnzL1wPTwItQZK/JiF+N80YjNeSu/dmMwuhQyj+onNeiyx9YzLdNnM5HbvSfZSw
0kkAE7lFRAoZUYeCO5GY76eod2WwqbeDWk54Ddjehgh7626bzxuZc3hGg/eo9AB/
4HExU7XwMMgD/9/yvHbu7JBV0uQM6qDiNK70lYNAUL1HLUjuUyUJwLxv5hK36jh7
I+yYPxJzvJRwkXluQgl4W3VyrSGaeLwMJbnsoG2sqEu7EbLvHk1IDCzaeu7O+pxQ
xr6hV5+4u57Vy8ZeNnwE+DXKNhSch9JOhEkoLU8vQRHl+FSDmBBsyEoS6V7StVxw
bfx1eamK3ZQFpgnPuV6Wq+AnfEj916xrOp9F8aDPRq6Eqb70QWgufWLU9wLDAkSA
bvoD/kNFkPLaFgEmFK+GSbYV5L0Q7l2l6ilTHMZReBA5whnuX+tBTI8UttRSySFp
BgP4RLfZXB1XSGE+7RybvambrNhsL0bTEdT2sv3sUF0+5XjPUVQFHcS/pE+Rz7bP
cjHHFvEWEk67q/pOjl+e/4NmkoKGPpY9lDZ3/z9m9/g7u5dgSE2Ymhdq1zICCTcG
c3HUUxXqp+ZY/91MActFm+yBNzAOvdiBCRgmUz3F2oVsBeQcASJ+ALpRtgZU3a/P
xlfQk1lVYs43sZ4GYLcjJ7AYGUVkVa2hVuWCHyeuvxvBcXW08PHd6sA48C+TErro
wDW8cYhc4u4ves3OHiV+ueqjwzmTZpy20cvqSnVwUbshgw2SunUat1gzY/Ynwgyg
8q+LCGn1G+XFeAIiTw6ykZoIZ5eTqYhattvTLdLe/b+Khq24fY+BTFyi1gzhERpK
tUnuhMsf0xchm0SYGyiaRjWDRxr9x9W1Khazyfs4TfGS0+B0S7QPpmrR8qve0z79
Ag6VJdfJn7tI8R9mq0YQ1B9VJLIUQgSNGT+TS32oEvPeVRI+E1X1oyxl8x+UEg4G
gXPKFLoF01yPZm4EDPLeKpPV5ikpAMZcxCNYXsIVt7U4NTfF+IYoh1zQnWpSbuSD
02H75atRCqs28gww7uY3U5T159p5qvPOZdGnXAIImGIBw9kJU1s+2UyLlKCS0aX+
YkRzAmgB0d4J6Vh+z7tK2w+XMWNghOxTLW84N2mQ81Gugcl7iGUYDCmjqIHtzmps
ZnwzA0PpfsDEiD8SIeKsro7/o8WFw6samQsErGESticK6sHMTvBL1Vc4X/anOGYo
W7adwUthQa+hgJvhsnV9zLLTk7z7RRmoZLYAQm9E91b0h4uIHS92gn/y1AIhkN8b
ZBQ++zVlTrdpqs/bpOAvAbXfYjZWwYoPAgT7Eq+aQIze+7Bt11LBgx1ddQ6UQYUZ
/LzQp/YhvlpH2GBOtXtFJ6I1pD1XEpM3bVT2OBQaomqTzM7xK3GnbuZekYi7E8JG
JMYiCxmZ1F/dK/j/lPVJV5rvDpbZ3wC2r6jNV5htvvhkG3BcmDXb1DCHfoOefPOg
/wG8p4jsO3EjexMDZTadGAeaalP1uC7OqndcS7lZBlREKlfj5VnN0ROxUfJo4USH
q14q+FpvXlx2eN+XYI9ldSyMt5ssY7874OfAsEWKj0Etaa0v7to87T3YQghYtS1p
mDWSz6SuSnWzY0GfAoMb/mNyARybhFoTfJKLfwb1OKfDfZX9u2mFEy9t47Sr9P9P
rM+bbIZn/w8A+3h2q5C7A5aK3ftBO9ltTOAMyQaggRLuTh2zj9d8xhuDWeQjXRbH
jq/ptG1cMGqitR6M8eEy5v2ZUVyiDobX/zKmjVWawO34gsSLKqCWNLp3NXTrjj13
67AUb79d4fGd+MoHA5KoB+9WHIpbnqByLpRStKGDWpD+dsm2MeqvG2RjSDx3F2Vz
87gOAn45copf783m8QvSSQX0PVAXFUr2YnRzhsnJDe3A/yVyS2V9ccS/qJChdn0f
XFGjRNrJlGMdZUVhLKAKzui52MLJpREuz1dULFCDudbCQHqbdbDUoHpt7eq9RkqT
Cw9k92JY+JxhbJmu29aybxnbQxdBu+WOLNqm39CkYpdgom/UMv9ZUENSucq2AkeE
+gLcQvkCFzw90vMjnQ75PDRIA86WZ5Ykv3y1H9UpP4Qs6Kuv24F8nd6FVhyYs0/X
QzSiGCojvuBSZFSFtb0lFX753FCTb392oFCGuFCE8TDlW4k+EOetrP0tEoI/smeR
dpiddZti0q6bKZ/IMqaGVoV7fAl4Cbe1KzOPciT0Ry0q8airdhRZL2hbc5ZmUFmR
x3d6NHFpU/QAt1vCpE7yulCxuZrZuQCOOIqs5jvfOk7tbGvkelga49+GsN67cbxh
NOfMYpIJVrDaRnxSey76sp8yfg0SdOGn3j1OMjZj+pgvwobulPE8Bsupqk1OEjGQ
mBDBd/AyI0AB0261RfVFg+1FfIBjvVHP6U/QZb4opiH3nhbNnFkEx5BmDQY6+/LS
m8GrARGX+9VrhjP1K3CQ7U9St+Ko1YDfHC/ukpVfdXFImBQas3Ac15VExwOyzIxf
0y29VHhwz2STzME5Ws7bi85IPfohgO5L41pw03cB5sVZEgpIXQ6ZQdJOHR65uQy7
rXC0GfFHTu2CnreVCE/RXlY90kSi6P6jutJcQrmnhpa/vYhsAaqP7SFvSlozn3uS
SHYkSYRFa7FC6YbB9V7lwGV/M83jTW+6QW1hA4eJv/Yf5yU6tirwRX19eU1nK0aU
vHXLXgOtQEvvaAa6eLWAd3GYk4uCBURKWhNfdtR7sazOtw0GrjXxk8thj0xE/sho
QfExJ5tVvkH9Yczz0z5ca4i4E64/QT7Vr1q+p0NiSj71SEhoYc6QgCoxFdym+xPD
voXCNdTI10VMceUKR5Gw6epvU/t6Gxd3SsKhJMvdY8YzMOMl1mHqhh2u8AueX4U6
X6bhIY0LDzKzK4s6bgYZsybMkD51ugPB1lV9rMiD8t3yUfkN9DdvUATf7yuH5Pok
3P51j7LfM+qsEg/h8NbY//qHDIb32sXi/f4jqlNRSoHeZU8b8RWiCNGMSLquxA0J
gtg1/BLDZTfm2z7pDvaRCbgI45dmxfh/T1a8A/ZxhPHE1J9VC5iVS4Hlw7gQADLs
MQwXcs6i/iW5vIkZfbPuULMYAFkejWJ3bt6pKnvbFA5qxJb8ZMOzlm/RdQf+dtFy
dDwQjdO+770gJlMAttnajr6tp27sSYSXsSybi7Q26bG7zlEga3wUkOgfbNry3rPD
koroNcVDvC9LMPVb5yMcoBwSm96vlpRF2d1Zcn8GxXpZmdxjNhaIBEkqlTsdF4g4
ebyYxHav5gvB+/cGjdzo9tsXw6vh0X38Ukpn23XN8cldY6Z3ex46W6Q35YYpaLIt
2PdsEuD3mLslkEvUfOQKJyOrC0VZbegq+LHS2XcTh7MfGukVX5A6B2paFW3WFno0
J+vsMOrW0WgZJuX76L7MVXmGs0j19Hlx5MzSzhyW7W+g2eIHmLwDJ80yq7QFY1Sc
/tkcHLAVO+h4oIHHxrWRSL4fIvlovVyg361x9QYqdEc4beoiH2mTQxfb+13sNU36
gdoiIJrgUiMRTuirP9Vdb3b/tQVytQCTwzx902Jfe9TEqXaqaDlTOahv+da9Aa/q
el8e4zf3jGsZNFv5Ch//HrG4yHf7PnTJTvWxKkh8RMvS/JLKLzL4okpLWNHijFHp
Tdl6kERlP1Lj0twu8OkbKYWLhY1WZBJPjiT9d5ouNyoRipemrSWRpeAQRwqxHYeE
KvoELl6UDRetgah/b9oA7kfAFTm2/TYJvcnN4UWEi0eH09VQcEnYO2iPSwUWaK38
IktKuRtt2bzeAkyel34koWV2fxHvtsNy120uqY8jO/hLE18n9JDk3ocp9CKLEmoT
FyuJBkH1yEbAttJH7XtgIluI944nzySioV8ByQ23v4lrq8cZJ4VCOLu80ZGBXBpM
PHbwW5bCkUFTB3mUfDH17Cmw9N+PD/epnWnNpGunmlZOJ9rG1YLRBM7FF5jaM2c0
gvkXkrat+YEAbLNJ34Kutlm04k0qcklGrqb341+BhNsss3naXmQXy1ZQZY0tyYBv
8UNueitFalwjJEuO9vo/AB+yMLRyN7whAnAEpVI4Xqjg/vSEP7TpI8k9FbNMKspt
wjwqaEywZssjBKkOJznrBNVrZw6XDYqIFWtq3KIOVccj0OFJzJOV7jgfdpm4fJ6Z
vGqoFkInKgCnSLDTF5fihFxLT5esi5OJ6zUZOrfku2Z3ZlyxXq4vp9d8fj1WM2DK
1IaBcplDaFqRpAzWdXQIe6L8rdA1+01RWF/ozn+PXcM9JhnUXJvcjvIAtwQU7hOf
b41wEfnS+JV7Mdg0TfaGBc93efy98AjMdGtW3gM83q8x5ZCgq7v0sXJ93+RWB7NK
6LtTPLF65jeT1f89w3gdqUd/LphQtxonZide4wcFM474A2vqukQUFuZyDE8rd9fN
wyeQHl7e4Io27ZvFoS1fnMslkqftPaqsUG2SJpNvbUAopK5NUwHqfGpp0ySyRvev
+ZT7AJxKmJH00EvwGbxH0xaBL36PsbvQbWIyWvpxpwz1Apz4W4oeP4ZDc8mdZL53
TF7DS4N5W2oHdENeFwts3WvIg8d/gO+aXt8tTliRdoWAZPus2PfVa0FbZkt3NIEK
vvTWI6TYZn89RbkJmcAD2CvZPM2j4R+HddIAHG9SEEM0ZO9ChfRfx1G89pv4SfOX
oBVX8obtJV5ZC26eNa2aiJV15urEBCgj0DYgycdZr74RvTTARiQmsgn70urEn6SH
AkddUJFr+WSfi/TSgeL07jxbew8g7vCmpAEHXV2tj4M9iWrTbF/dep4erh29M7yS
sDuqq8bGkgrhhVWLTDWkgKvZlnQn6sNeSNajriJ85SQJDoUmaXeG85OMeTjGgUft
jMBeF6WO+oe0tBPSHVUmt+qDYzntJQWIXRmZgftje3WwhHpcysT3ouFGf5K7IRUM
PfsoAyHO/m3ZH066kZa/IbKvSOveZxkhK1w+pVSLA0m8e+gnaA+FL0ITnebB1jwU
tTUoQcgxjtpUOWpKh+yRo83dsqxoiJikgT0C8L5Wy/d301b1MdsYiNtHmOX8wVIP
sOxAhBDIYgZSCJ8zwI4wxrmKF6NuTnJ1dCkx7Scaeq1XgZekn9Cn8NAeMMZ6Scry
bDqXk/p+SdCdz48pl2KXJlORoWj6BcOB22l7cWFanTpIt61xTHYxmTjFZ1Bg86AQ
Q2/2wuUtQQyopDzOrza9IQ==
`pragma protect end_protected
