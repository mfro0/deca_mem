// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Ev7Su9pjtQX1BmHVr2ZNki5PH0v/ylvKySKjPCzR0ZucUE4UBQ96kv8g08JOdjHm
FqqF0EVks8fY5vQvU/vKo3hyyRKQEk4Vxzig+IxV0N0slm7PdMkWjgnb7ResFXak
WjpQr4LRKIgj/keQsTm9haAz68g3Wu1Rup7zWFmNZKulgYspUC0oWg==
//pragma protect end_key_block
//pragma protect digest_block
5OHuD1Dx7bd3saMIjuxoTgSxeDg=
//pragma protect end_digest_block
//pragma protect data_block
DEZEYOn0AQQbBMS2Y6HM+oRpkA6XwZlvK9RXcA9b77W0Dfyhj5T5BLa1y5A//i6N
07BNquLk0yarmw5c2Ph1MOaxrMTrHeFmkvAnkafwkcnxPnteyVEc+xSYMJX+66hX
YSOAMeqxWDc+LZmPevoVGkjbabE6XXD1MC38XS/MTOkUclZUYScMqgrYbv3+GC7t
eKbsBl4a65Cu/7BwAvHYT/FJhZVMTK3nURZj7s7Aecrcpy8OFdK9s41ARJPxGA32
OuUZ0oT2VX22hUU7Pkxqanyn8nSF20frH3MJQMPZ5YkLNMGLk9jqdHd2r/g2Umrz
axsvSNOjE4RJWErUI8oUbooREKZkyNv9aJMhiWIbydEl2ueRZBCxYrEHmIwMacb1
b6PpwHCt2kEX7L2IE2ZkBk+/8nqubcA8Ny4nHrLABCk2h7kje8nRrQk3mnZsTnDm
UuSog1F7h1AsceqoNpWsgOTVTSakjWoepYOmPswMbv7LoLZ0G5oEji0w793mgBhJ
yW7rixS8NZ/d/IwVlzIM98dgPpMNEa2pnD1893twCE6jxeTeKGwjXCocE2IVq0wu
AtEhe3jeXFd3i2v4QrBphSK/cipR2Fjtg1sKtx16pO4ILHNnPjs+OFjRx16Ab+H2
Vx9Xt9iDNk18MM7GDsOPfW34ZP8BVoPY82FQCHWdFmxhgI1sLjFXk5uBfun3AtzB
yZW5lXpJEXMwlRadiPrK8yaQkXZLr6pjABB92beAqNRx0oYj35SHwx6kSB0eoYdo
CpTGqgx8V61WCPHPJcqHIRWZyI+B7qvSQgzxjyxn3WNWKlw6SdWWRrTOCfeR/QqY
UrXltl2BcTZSa6wcmTmWjKbP7iM6E0dXVXQiJysdSagL+zKFHTpQJDQJlVMXcYaG
pmnfOpiZlxXrT5CmA9mbJRMQsmkJGtkLJBRCwnGzeLLwUbYD4a19JABOTbvy28zu
Mv8kxfD/5Jt/v1f5BTOlvLXbOTlXW2ggjxnBgjgPADPzMWsWIv/FOyB5fqicvCTH
tWM4nS0682y1yQcOj9SVrm2MmeebgBrneouENBvS7Jism1s2p2YAAPX5hbGBXFeQ
BPZK/qnbYUVfxUVAwURsa8HBj08i23Dvau/kuL8z3+mQ2O13q5WA4toJGhd5LMAd
+DZ/DxT+teLMyhF7Zta4Xo1PFfjKWXbuHbbDhWXeiK5X7k+9DZwbccSLSonYg5s+
F8rbn7ShRaRcE7j8+PAqrjtL7GcEdVyD5pOnxNeZz/AYZPUJgSx4vgCCmmiiBeGu
cTys/FioC9PadlKV/hvFb6G9e5L2alabHRXrqDjeDphCOdaQd5pcrZXDKpYk4GFL
exRThYJA4sqRrxX8kcgb3kycU8R8nBMZcgEFdVCOigaFwT/seUYgcllJLAYijbr9
ohgJZHONmPdRmSMBpjsQmBN1cowgFRCuYiPoTzAPTqTd3FyKQTyBo7Mfu4lGaBxE
pcgoqYOYLNbf+jdNUhU67RITPtqynjNqNhxEwkMWRgvvb9q4cKD+pDBatifl9rAA
tVH5/tS76VbbizBGqwjy9z6WFVOuodi7AAp/T/yJAY23xle82xeYkOi6kItOAvIF
MwR2sUJrmoQMkuAXgdMlsyZBgMyZtC5jIOf9Eyhsu6Das49VblGklMisH+ZbqZU6
3ZjVhPPuq0cEAwIuLStKrx4tsOewUfEieTTmrf5NUnrYG9dWloINjvRgXLJ2jCo6
r5qOKUPNI5W6gQzEkhcJMZNgCxtlzmZmrS52TyFfscApfS8/bKdmn/mjw05pXvN4
o14YeqGSTzc1jPnxqkOP24zkdHiK+bORu7Cfp3TqgQwIRAn/AsmoZUgsN15A/16M
zcDLNgV8zSZMbXIvW74Y7uGIrlKubtjKRddykVfdE6R12GwcczdOj++pga9aGqaX
90fdAfy4URQ2iU5XqdF6QAIFxX4JjFyaxhqES5V+Lb5Pl2qMeOkKiri5gUOXOQaG
WXIaUS9G6MNErPb+0/GWhIdDmQuTea4FmpEZGZIpK1cVfrGYGoTMPemciwJVJc8H
dAMaBXxS7vIojZVJ/A8wwLIL1Si0A3ipomxMKr6sLwF5hLgH7a8+6zfRmHtIN9d9
5BjxpxJ5QXgclirZcjao0W6fyLkPZhDcytDGfhONHRCiuh/c+Na5AFgBjc8OSDWJ
YScDLaiOhxDygLoi5zsInIDKueUlLcGnIBKW/MhEcXMuMEdXkvU7HRfggsZ7dzr6
Oo5b2RvNLCywQXcJEGsibioaPBl6Mb+yaL92cEPn5ry6U7SEujbO7YRZLt7Xd/VI
rlS62HpS5s7BettQb1oQQj8I6h3k5YH8kgSdBdxc4W1WwQ6fSclya5d2U9+pJYT/
BDJJgadT/A30wcKuqFbdDmjQ61RGXJqEEuUcvq5b0/Ued6YpaBBHLNwsUlGeFnuC
F4+d7F/LmXAYUfy9YpmggmYIPGEKQ2ffMyvjlywBEdyT2tDIgaVwfUiQyFGlx3iH
WA6PphS+Ztiw1Mv+fCErD/b1h0keEdtkoEE10kXdHGA8U6RF8m5W3vET8Ggwlp2g
wHivv3ZkCe5z36U2JoKYI2UwooU82nX5Ml5WPNXJEcqAWek+HVHIU82oWACYDGzS
Ajt/6QWIOd5zrAwyZfgArTaRk84Geap/K+dzU4viOTmQNC65gGC5WbWK+6wBX8se
I7x8u8ZY3c045kJAIDpOcDxPHh9ZBOuZ46iWKViiAlTTbxoAa6I6xJ174uEMh8lj
t8YsTB/gEmS2zLG9M2q4W6Nw7LykdFwSLieOG9tW98iI9WkagIuWC80lYSikU/Gm
UnS2QxJOmsDZM7qYKkeZtQOq00kyp2XThP0Am9brSTdat9cDR2TQnWxjr4Gh+dvp
Nqv6VyqUm1LeGiXNJPW3Dg37c6YmUkGtxdiNASMpr6Ef8eHmMibOFPwgmw5RFpS7
uMHXbbejtcvfbTqLF1R9BS7Y2irFBJyq18ozNsV43lm+7ZCNV0xZOX8CNKPrqz3y
ChynTrEDdysEt2QnttOd36M92RwPaY6lz8x7Q7+33Ig3ILI6nvHj37VvTkM276tB
d1Ex+nIV/5EPTBvPEUFZ6sScGNn4f07rQ81HrJ/RJJbmnRl3P4y1x/toVjNLq7FC
lBAaIDfXvZMpVZ0wiMDb3HxYlVHEVCa5JIZbW38NxRV1KLNA7B7k8oVK6rAf4i/p
w2s9eEjcDRZiDvXP05d+ksbiph4Vo08TRXrnA4XAsoEAyJEUyYat7dFWKJ45Xqz3
NOl+Jonz1qcnsX1mypmMNq62ERR8GafoBoeVufXTryozwe2adVKOB5TDn7oKICuJ
FK9+FPMaPldOJmAggFNPSP3bFnTpgEw6WxczIj05zBYjjfh/AM5PO5GBeve6/G+k
zJsJxqTrcW7fB4fVEPRSbSdacomhgRVINqTo8G8rIDiaUUAJaqg7pr7x8M2IoIZk
84Bkgh7JSpETW/b+eS3p3VQGtXKXaKoPRnsuepqfb1/6281MpLNovZyIiaTrq2SE
0xdUN0SqbU3Nhs6zskwjgcrij/Kpcb9Ss11dd2QBb07MVBmeWA6XSF+lA4YyL6/0
4MTrM6Lm+27i7oEN4hxctegOQvUNmgVNqtx8spJxnLPVG+B3hojyzlcylrqYCx7n
JK5nxR1BjTRcCwNVlWs47cgTiUzszXJ0EQnYjIAe2h3KjVzba+nf5FqH9MKy9Gd4
GK8UkmS/QYbWXfCh/r+55SesJE9k/gOXKz3IkDXXCwNXYkWrcL1ty0JU3/PWcIcl
iD3/wmWewXzPj6QNLhMVtB3EOjf/OUTQgebTr3icPwhy3KNFRWFrNy5qOZx2ISS1
qgbQHmEgaVb0xf3Gg7S4BGdxv8clL9i5S8UZm04YtJgK9hphy/I+ieKqj1cJ5Ref
PRcBEzdhc1KUMif1hZ63PKd2+Ymc9OEGpqSH6PSfWlknbuo0CSvqQ7kqCms4fjcC
maxCUr0hjOf4kanViYqfzYZf2kiUy1N2J2+ssafttT/XII6jaEMKNBXVv1DFzF6V
CUitpNqEcn85s701uo+eXUMeuaH0OGAYr+8pkUOUDo1hMejgIt6Z+DfRvJenJ3By
laEnFfPKON/B+rYaVxGhTsIt3ZaJds2fFqoN1F9uR7OqxHwvweZMCUKzfM1bz5iD
N0JH2/UMzCkcDSoJH2irVcvVnYVsPvy9/a7v0BDI1LMrD2KZQibyviY3f3SFEFbM
7XMYjHA4jLa8Oorna+nNoXfC6KSs2JL+QyhcK0NTvackp7BrDZmPVOh7Mn5+YTFN
vCztjSu0ybn4Z+JH41BKmfov+wpgl4oehF/GLc3YzO/Qtl8dAY+y+OMH1fMK7Ipt
NpjgMtGPswK5wq0Yl2ay97KmQ33lIgEkpjN4xglyhjVzb38LeSi3RFtkkjTcOTVf
eaQK6qljlhxKbLSrLn8gswXPA6KOmV8rdbZWYCMd5vWJi2X4qNkfSuhAVhJo1OTe
T5ULk9cRdZwt6GiZ0JvwJtzGst1DH+2qZVEVfvaWdDHR8apyJM1+n7g3D1giq7nZ
j3mzhvaCWWO2ukz88UKcwcJ8Bl2G43nl7sddrNVTweDtP1PPiE2bOwyq8ysO3BA5
NMiDw41G1DpbqnOPNSVHJmKWruvL9vlH2kdq93TqC7b2pD2jQv2sJErrXI8p3KQC
g+ZWe1qrkZAzT5msObyfgvT3hPKmb4DRuejzTCae3EWOzcv+CyIkNjZvxozJty7e
ftosFX3NzMsQPFZcxF62CrHO7oRm6jGqoboF/3ItC4Ong5LSF5Bj0FxygHsf/+TJ
bfGqsC3hjCTBL+64OBmGNBcpi6ZwQQMEA6mqJN1HJ5Nm2s9c9A4fbc+59szQEkRT
SzBn0htOZKfG6LPJ6Hwde4vxiq9dh2/0/MaZB4+6wgEyVNR0KwEusx6sXlz2SJY1
RDiY5kcK0dyRnPOfog25v875+gj365uq0WHaCPsLChUI//0gqqWcSEyDjpOWAyfy
2QnqUIw9snFLFRWFQ+IR3+piA2bO91kymUuJQi276tD90nymrLjizKwb2CJKg3aB
UNiC2LCCL7kbHN1eJSsia8X6yx/Or3pd27OupXUgrQ9MlDx+HacLvgmpb+bc/HZZ
8r86SQVGWdeQsqG8AeuEhsPmwX/9RmF2cpWyq819LqI5jMFNkx4CjLJIqWK/jLt0
+js4ntVjl/AxBqZObhV4PAyQqeoDFWsUbRGEgewX5g+oIRtJj6cXkXq77qoanQXy
in3ZkEH/QmxBxaNMpL4lP8h4VSt0xrYU4x4NZdQ90sf4s4uswblW9Rwb5lb4xrSp
2afFmogGNqQNIB3rvPznsqhVWBdqwumirTp9Ro3YfXZAyfwauYY8bys8G941WEew
nvyaJM/kuN3M3F/WtzvJlUVKWugN4lhUG6wGmr08aySqe5hr3aEfwGm0+bh5CCcC
h9tUpvGfhC5//xWwlsqPEQNPUix0zCiJy4qZ969Y+FmToWVVMJObrKp1A6mYWsZe
GcgK37YEx+wdW5AVoX4jHsEejzVHp14eKePBRp0wcfkB6Ej4uBkqToEaXRFE6984
Are/YQLFQq0V2Di6p+8az5ML96W6w/bOuAhNnifNMoW4Z3HoO2m7+W/YkrJPJIMC
uXKsuLfLEXImPsD+0Vkl+wJpA1DUdfRWE1WqgxzsgkbpMFUt/oiGhz/IChly0tRX
DGdnzROyDoKVdYU2URP4mELpacYGtGGvlwwahKVl7sJ1HGQ5KviZ7h840R+3y6F9
qF6HC96qvxvwmHOOZuFMeEcqPCIKXbWthDd1oteq3yrlsJ2Trvv7GCLyUzVAat5M
FEO5G3JJnpCuhPRuf43YvtcbByP0koRRR1QMszXHcWUN/gtBCfW8myC6+XC7LQIJ
SipYBd28z4tpzKfxj23nesj6cD0A/fWAhuiGczqvQcPToCAFHINpLKPzoQhm8OVA
V8k/+S1NWYN5xiikoQmkbzRpz4ZIrWadPk54ei907jytQASRll0fgGU26ZdFuZzx
rMjGbRgOnL0AkfPdBV38pNuXAWZzxY8LMHG12sK2xqFRY9fSc35u9LL5p61tFrwK
M73/IxH+GNQatcw9VnhVl8EMbZ6NszTOwfvYEnX5kO7dnj48VobKzSlHAJe/heD2
pwxZ9kmAUVY/qUYJC9PoGbDwFqzi2Z9USMGTUOFU6TX2ADaNq8VoCljjg39rq0oA
pLRJwsb1/euZm8w/ugc9fCk0vN7J3Lm0ChkrBYjTjL8TQ38h+mccFrSqXK6/kgJY
7LJ3JTkrlQKByYzNDwkENGYyIW4JDT+VfRZ3cxKWc3oMaCjNkdZlQhZ/5yt31QOY
uLmlmXcrtw7SlMXmD4TuJ35dFj8x0ptD6YObMsEfwMGinX5jKppjYXdHdLgONIjN
ckIksUivuAjDSmwkBwDJojeRtArQ0dVBh1ZA6n25foa7S2OsVPqQQ8DG4eR++oPv
+GciNP9h5CTXKPtBL6EuFfyxLjH2JmpKi9OyWBUddLxKEYfnaHROns5mjhatleqx
LUoyRi3NC/+hB5EqBRHmmAFhQuoUiK/L84oIZ08cNvHhXcTdaCMPBvkJyCvAt012
Fa7664L0bhktMES/oLZRyUr6iSPCdmdMjoIsEap81wRnd+ohpow+uiX8ZE5sC8TR
dFH0dwbueDBcY5+YToUI67WB8ZewkApnXQhcw2VJLDTJremi9s1hr1KA8iF2lKSn
Qpvx1sTxrrAxV+R/uVflr31Sww0glYEUVNDaflY6SLkBjJV+gxauzAAA/LJjdSET
GQGJccwLh2FLi7rOaE/OJ8Ykhl/9MNlwb7B5EHfKr3uWqSEL58o/IJ99MZndBWJM
SuyZhqn06jo1hwh3L3q4gaJcgcd0TUleEIbD98HPsZUH2ebEiiAMcT5NgDQtDszW
Yyts1Im0+7l93XNJ875aaQAGbPX/Qw/vRachUUePKbinBbOxjkSk668DjB6UYBqp
KjuIYarij+yvkNZe0zY3oIdU4EjMmD5og+6Di2r9WAL6bI4UjlC93dhXz2f23I1d
rf9YzBWnd4ZVACp41lmLUlggNtBf25tkTg3iAtmX5bw4aKLhrw7ep1fNmDctS0MJ
p0wSgMVektyb3okpTP/oh57hz4N1UEFTqyAOFfGodNoQOUhoL1yJM2y6HXI/WQ6L
XrWI6iDb9YezUE/SR47HRhWJW5q55+XdolcYemRI1pI6T+p5Bsisz+h2z5UiSYPf
vAzF86jJUvV1uCN0NToBgZ0sKDz1UbDEFcvKdfMzoKO3urBHWtVEkcl/oz+EOgpX
W61ZNXEClvBEpLZJb/zJZtyLYxOyz7JfF737YPv6yeQOAZaRtKrmndM0YmHjuqUM
Z8Zkmtf0TN0ugsH3VXwSLDQ1JW1ugRu52OvIQkUgCRKSXwarK0BXNn2C/Mi2YbDq
91NfSRKhU2N2E37DOMxNTW5dFCh6eJjERp577QD7cOY5VJFQxDBGrbAY8aNPvEbA
ULqP9VDfdX575qLQvcIxc6A5YKui/J6tabgNi4t362M+cps6vjqXgNSTfSIV4TA7
EFXIxfXTbcTIuaAdv3CP9tmq1VwrUeIid6eJ+BvppZ19UJZX6i6/YDIUwUeJvJy5
xgi6tXSHtKZGx/1F/fWR/UqK8ySYVHsBgyr62EJ2qOoQlQd5qAfdTskLNyZHdOt5
V6tnHbwb6sboDydInkinykjXILHIB5ltdzmmlnFImOcNv4weRW1hdHM+WP8KrzWw
bOTwBCNqFjRy/7FxC5fJrIqfSxIQ1QiW0l+w8IXKAXcPRMO5qjZZ/gfrDqzRILi9
wDefKWfRs7ZyiaV+E3Ll5bpIvb7I0g4mkKnIfeEA/bKMcatt5qkPAFL5h1cjZVXk
Vj0lI/BCSijq2nqGH6tAKKdBNvzlYoq8XZ3S+9DirSjO4BTTFtqPaBqb/5ZWixA2
RNz7/OoYmiZGJaRN25SHxeCnoCJR5Tp3D/eUF9nO7ZSorLLxpzc9OI4ZpSKDFoRy
74KpzxHzsYOpl0xk4ZnFlgPrh35evsClmXznPCoz0ezHIySJk6DRzuHM5h6IFogQ
ETZCm1SjD3Fv/OVnaRplElvIGT9ulKBRdn2iwnOYr9K7dnHheTbDX3dDGgwPZSG6
9sdgottN3XkqFqLjQ5/ZsA8cBH5Dmb63GEmVTLRCzSCiNiq9WkhKuXySXlkIuSqi
xh+yUGb8Uvuc1uttJe5hc9cvkGJu/BPUtRBmXPgLZZyfwCH23CqxOOBhknPqbQwe
APSdE/IePKDntzqgiAr9A7kEuHduJOgaCc4PA9iTqwbimyVZonsM6fzMMvCUan2d
Lx+PPMZ0rWSf1PZyuKHF9uNZMwTAizMeM4H4ShwgSBj2/4Gw+ucwOCdCyqCSt3Ub
OXdHcUbFl6lnlAshvZJyWwUvznYr3n2to3i+Cd8EwEpT2sRzKmAUtkOt7NCUjq3h
oz71ZS/T+39pfnp5ViU0M+/U3T9mOY91ZuztcrEKMOU1TTI2b+idgzk9N1QA5nbn
R1HoSsXG7eIe+FGtoKCazi725r90FcYvUVdEEfUgaVaawRRd83/ETHfZg1PaDwyL
j/qEZD/6RtoQ6cKMVX+j9FKXSQWJifQN4ByCt0zGuHDH97+VkFMbKp90ltX+Nhdc
GLCJBhJWbUWEy646Z1ndLHBJ/NNPAr+DPAWGwSJuZxdg1LpVnXSbyCpAu9vxoieG
ueEkfbAtO3ykui49zzJjsDuWPr5481dmGtxei4jJ+Tg0KNrBOmnMakwe70ra0VZw
25/jQbyGfitnqiFT2UINLUjYU5t+mvkzYhgbKf8iD/IlhN0NPNsKh9kXRkZF8o6K
6xAM0GQYgA5iVwVPvN7M/TO6YpqAU3p4qqIK5WkuHQiee855hfO3bFnKjJLrXi2A
aiFHtI/NSExn4eiRgqrMS1M5+TNBdrxHZ9BONUkx2hVIYYuqC/468Z6heZaipPoo
uajxLhnewp18Xxfq+qNelDzg6tMfN5a2RquezCOAWaTUEnsryYpKZZE2BWMrThYO
KfImAuPuEXU2u2uV0j6pX0ZJmWIEyoveTd/PLDBTGQnt2+r944uyiidCjqvC4vNa
0AKgOH4ehEcAY2mrRkzCSc81B8tXMelz7yCwcnobDfMXQxaxbVobzYMBwuvkzYbk
kCwgWi7R/7M4qYvXJfsIhhuT5YX3Up116aIjwgZ038nlY+NbEPWuwAgeVxTY/x3P
6eIZ2/Wii0rVlMS4+yQa5su9AUfJ6GWq0wL6ab2okV6M5n8/8yl1HLXWVSxi/uM1
pHv79aC5QDHX88FsV5CURDUqdDruZmWh8P6YPkCD7iurV3TH5rDnWOdxuSA5VFJq
7ARYAgktNgPD7ptZQAyyJiYaNGL4yHAVgaoPnmuLKP5mlq0RsdBWVHzgsu2s+ULj
xw88wUHes09+zQxhTgfmXfb0OL3ONQ0LXoNxAqSJ1onHt5syXQSqE3tyWbYjnUB9
/QKNhxTL+jmnV6nRcsbTgc5IymwnSBvofRGB7DBXti0md4aUmbzFBisPXAcT6ExD
E6qTfDQifNstqO5KoKcnl8qKFrrUnAfzhbmARJ6NtoJmfJ2DHGQbt563aX9H5kvX
knweoq43fb8RHRQGrVBx402z76IVVe2wRxBzG/eGQywWs0f7NKkESdXYD32CGf3m
1YThT2td9PiCzXXUA8KBRgLEHPkgbIIeH1K5IT2euSVESss/tvjo6ED4EcywILXH
1E2s0c7pUgbjCQiPQlhOTFiNYAEnuZY2nAJceN+lMqGkQ3Dz3ErThJN8MFqgUBTO
XLc2TYiN/loK7by/35X4E/VLhoPM6r4LixAgczrda8O9GMrOqkKOsgX1UH/KLtt7
ZDSFdQ/y8Bktk6lFcVo6ylwGfioX90Btb9w4mXnWuOviZd0MX0rO7d0h8Zl06BNM
aPjTngE8biFzL9jpSMRPwnELMVSDWNOkEHUpKzFOrbmlwuplRHdiJb0+cJV6oxYw
AQSF5PNIq9E83nai9HUZi0+tSTs+hbthptw/BG0EAL+8Uvc2dSEOtMDkd4T1+FJe
EYb6OEGNlcmpE/57IMMpLvGFXo7Jv3J0BgR8tSIZmMO+8053Ek4vo0GCinMga1ja
R9R6MEXQ6yTqqWsfJbM4HI6rTlYPzOqs37+KFXtq4edmjysQVULdJPmSm+/iaM/f
wKsdINZ6g96NPsvftmC9R+syK+4hIj8tNN6c0FaCdV/ktUuDtn0920hpt2DX8cBU
umAdzC0QclZCA26Q41ZvAxKSDlqJr8dVH0VQFxpvma40z9ZbAicKAWjHiFz5JiCa
GaD7mxdL0FOhcVq1YxztJbsh+/fEIz2As/EGnlJ4yJyvJQlIrP3NUS4FE1R0wo7t
AidDa3G+WA8OQQnMj29VmPDHbdjJ/rKef/nTCAV39uJSdUMdWvvH37wwLNQOj8Dr
uHwhbr+wWebTAzWPWvR+IdxuNQFraB8aS6tvIC4pU07e/HQ9QhYx3mrh77meSJWc
NbT0N0lLvVaMgR2JLOh5NlqH9TPmJxRrEOZHYgEOaXRoGF4tZ9uR1iTdbIBaL4SB
Wv1GeHqeH+5GfY8w593+XmXP98ldTbHExhmeNnXhZn10pNpm4+gVilo7pUM+IrOp
UR8iqUeORIDMk+FCb8RoAMhzJibD1nTKaNELkyUqoiJXQpp9Xv4Otn2BdXBPflLB
kQzDVvb0UXy0hq8f+ELrvy8cMkjjbB6B1MCBdgBNCZQIXYZ7SXTvFsa5gAVtQDsS
ObpbK8Qo0PQCBvOjNYDqO8ValtodVHuw6xYtEde7yh1HbSZnpanLBLhtkXcnLKiJ
QhDJX1KJKfYNEurbtE+gPDHr4g/mZJgptA/nEdZfgZ4vWxaFWAPf39Gie8Sf65/X
Abj0Uz7d8E6oY9o07NoyiSCJxKwYaDLheiLDfXIMqdj9irJDebWJspiMZRGOT3S9
LWa/eHp8yaiGBA43QPQv7V7sUxQv3wrBBCDfMWZ4+uH+EQMVfvSqs19ZQHLtGI6r
M0iA1Lop1kxZzPH+gOgMCEKsWaLDojJIUcN+LvG7DsMJK2b22cQv4wt297iDuIal
BmoiJUxpzHJPU/xHH8QFeScvxd6Il1daBXqCD2UfIsvmNGFDoQAI8tDH8f5PorEI
7GXeAijuhbuAVAL020PqYqsVhxB5CKGzF6j9fV0miUnlY7wn6x4yq29V5E0QH+tN
BhefVEUjHZGuQjPCXgAHq9k8eGvr2xTNm/Fctj7Ng9JeudbxxFBi2VGmXOgvaF9Z
33VRb2NcuGzKOEnswOKzVyleSeGW/x9uG+h5GN3aNC+8tdng/LLYsXOagnmfYl2U
3MonizpmvOUNvi4JORkx7/aZiXXQxVyW1V81Krhafw3y+Z9mvTl7HLUsfRh2BuNU
qm8vfOJ1GOc9wVhgJdRQxrY0y0SoHD1zT6gkGdTeF2nNenuYTU2F79NBpHecKogF
SDsx+QwXmUApJZznW7sJGm0YDI6LAWztr6eorUovgmac2VlhFZ0Cfqxeak1PyYgn
oguFR7FFHcIcY+ZivD3ujBsc43Bcg1dpsqEsUQ/U0iAf7W1E6EnvXnfaxVK9QVTr
L5SA7TvvwQ6LgrbOMc8Yr7d1Pi4ZttiqBfVsywHQ8gLp/fGwWkR9qsnPkWDvfdpJ
4up2+MUKtdiw4XppRdPRA+rF1l6fcrsU8sCWglgfsXMIqi712cBnvX4s87EVkaVF
AJ+4+n49XKaNM+FadVEmGlAqQAXZsLDyCzMpzPvb4uO1/peronwGq+lr6EocCYxV
f4tuRwZcHQaP9YU7UMzVsH/LVEyyoUVTcUKYc4i+aWJweE3djsY2Y652zVnr9Sau
G6CXL4LeDoFgFXMXcs9+zD5dfwVaAk0pYAd//ps6tIt+rZQhMU1bj5jGXkLeB15q
Jh3bC8jPPU73IZNq1s+NPRvH7nFNJXgMN/HyAAHdlUY1AeB14+QDJOHeW0Q9lI9o
RvWgKNaqLkj62g7P+fM8fXK83Zid61GQK0yJAjKvlcM0fnKgBVINz5d2mPimOHX/
CUdhlMJdbLy6VApxPTJUTGP8wtGYWtQBdr63JpDPFJalF9eyOc7OGgkgCqAx0XIz
ZSsxbdbRc2lqYeeQB383U/euEnh384jWkXsPGfLr4rMmyj8B8q29HxcZMMbRMd/H
bcNobrCz1bOkgdhCIQCXg9hxDY7FlLnpzzYGf6aqSAfOxcg2HxVWVHcF4aZfUYNA
9rY+gS8wLyfoDGe0AoUDACxdqs9fNh8XkpskzCbUnxi1L5ixm4MAx0lRy3YPpMfx
ZxXNBQt0AJQlBZF7N8sEbTIXEZaWhX8QY9R8f3+MOyk8pwtz20GdNiHm5thDNold
LK1T1B0k1ZDo0SBPt0zfSpQdP4nmwhrTA23/ZFErAnu6qNrh+sVSROaa3S6vZcY5
CKW8GHLtJ8SYnUcBuEmjR738Oz9hXn7MYClsdWAavrxPDj7LgAaQvidFNJ02GPKz
r39czK/5iz6UL2cfVhNhZFp13YyrMekwnsSPdsn3VQ9C17it2NhJNWEzXK8VTrLZ
1RO7X7ULpZIredIoidjFtLIveuzgwU0cC7cuJ4GKmNoKsIhNP0In2/sfJEgh3xeM
9TCgDOImjOu/GZUdpog0qcKENvu9Za8C4nO4M4DCMEtAH0S9mD2ACUUxFHWauNEz
wocU7Qt4NVkk/X/lFHGLliBU2jy+jhYbPRRmjiHTYE3NsBKnccBrh0jIP9HOG3Zw
wlAgo3qBqMDTRrHzqyhOgK8QSEViSt2hZadirPTeaXsbzm1dDsAvQG3e6DycY9WS
ltha7iW+uHfNUd6mpqOJW/aUnzCzJyPpi2J5xJDmr1bR67r5o1aC+401oEe6cDTH
icHwRG46WI4ZdnWJQYR4csG8eJ4sgbOMEoBq01YrCfKYmW1GglHa1dQ8KERMXCvC
95MbcrF7GZhMXuf9ATMMSMOoSkei/yLQAn2tSvwfuuDVMoGVtjH+QKITa+odYW25
1HDceq52GoV+its9v5tpatpXz2PT3rEc+r8BEs4cLQHELFQXSdSaAGcI1CEBviZZ
OEy533I7VyUewJ6Q2JbHCVF0dDEAeiJ8usS37dypQAhJ6inZyB2E6FT21WOWUt8M
FKBeWtAFi/GSJTjjW0y++6xxw1ae1Cv0ZEI4ScwPSrnK+vWPhTad97AgHxiBa63i
Rg9Ut+P9UUuub01hLZXV+HsYabYS+Ug6RfX+S3QLDF97VYE+W1p41LG3ijQY85IH
00HWfh2moCeb89qPCq1vhI35A1nBUaeaHhCy7wNqJAYrwNftqSHiOUFrOlfO52e1
fVMXfCmZSsMA3Tw+dv9pt6pSGrgvHZGBTpq+D4PHtbjqQmGQtwGcK/ZxVi/kf0eK
IrGm44lQlRYy1r/YNj4nfiD7bdPZFhIYquc41eVXVbsrq59oMCVpelXqSnp53poX
ROt9voN0wBhDFaFqZoqxvHtCpzsxzaHUpBRXdN6Lm4efM/BJfVdxSLZqw9jrt3Fb
fO91C+uL/4vvjvekRzumppg1PZFVH+HGWxZ4zKmUuWqlnFytZttQss14+wj7dAjN
QPFBiqwjT98I0zSGRvOXHV2V8U1XkO0e5icnBhu7iDhrujCGq/uDe9DZTRAR9sY0
pAXd+gE2+aIIpzB5tvb4ohbYDKq2qjQlmKGJKDiw3Ct+TSWE2OiCJeDK4FOJt1Gl
cacd/JvozGzmqqGpFs5q5mwwHvB8ToFbrIlsNrvERWuQPwS1GWRJAF+T38DcpN1B
H++MVcxgabmkKH1aaRQcvFDlrnEC78kBAzq41ocYt5P2lZGRZmShRue1kUgvRtTN
Wg29FRDedbnOAu+JULotowROSfUe/8fQJOZ3myAq6eqErMfDRMVG9SVIzvkIohhr
PT8tErsPETMMQIG4kZ2dLc7WA+xyhfrmdEeJRr/8zQmlxwRL+rFAODObcjoJt3rp
cqE1xyqQoRTsLA+IXDb5CfRD6RAA+fxAlWylq/Z728g0R7H503JfgsgObvFakkY9
CnVZ5Wrzu8MLiHIiPSc0J8mqQj6aK6ZGPZlHP/KSz9Zsm1sOrGo4bJK1zI4IyuQU
v6t5hL2b9Q9APWUCHi08HZWtJSQvwjXBOdWmZezATzuyttoBDSDuZj4RMoh3tk+K
OK1QtTnyq6YgeAw56csfnEg6R1m6rbSlEFtYiMsNVOkbiQzuFDpiqoisaWvIPIHj
MPcYGjs87oz4Xv4EXuhC2AIu0HuidxsewJd4oKlbpZBNyuEdkOXyU61ApIGalj6Q
Fr6MuVIOzNnfhUqGUUKrhKmJ38au/SB35yq1H+xktcKnDgXnYsAi+v6pdo9QmTns
fCyDJer2h2wNP96bpELrqyjhu4ZAUHf9obw8K9qRT3S4KAvndN8XFjTWldrM7QII
g7hAc1HKruVRLOoecbHMY74nQ3GTEKRV9q2H790KHJh5lRzzNXnmaRLLzD5i6Ry4
oxQ7IJb+2IxzFL7nTNst5qFalVmPfL6tPC+AGpeRg8u1XHIMO4m8ajfIWr3WHDIk
9r/Xt2qxHYhE7i+zlUUQjVSdIbo51Ag/TmnqKIII81yEorFcCdN/chx7eWD3nHTi
oEfwkWUJS34+qa1G9CaoZz6wGg8/mnA6jUjFQ4PHno266DXK7buOFtahUmsuyTLj
KNJe6wzu6MuUBdlM1SzMhOLeeWesZc1mMvWC6NSJrL7Lrf7zOCxI5qkMNkM9xCW1
IbcKeUhco0HeN68+4ngnIRAP3VJBzm6v4JJ/d3XHigy91jSICWl7H5kELMtLgFPQ
dPr6TVjN3aPP2o3Q+5FZTI1HJj1iW6sb6ncVbU204eJKzaZAU5nvrtkDCGRqHlou
GwX5mt1o/W0rTshjQhjzJNAiB31O1nbWZGMzE0UYi3HLc3EXxBr+6SGsTbI0oECA
KVj5pbSt6REEpZSATDcsYGySdsHkJk7IsE3yUGcQsQkkNTqZgs0YksjH9fUleWhO
4Q9pl5RHFYdPZCaL6XUK6r+QCZaN8ZAJg1CphTsm7ItccURk8MmiwxgOHeBGnPxR
wt3ugxlhfdJaIk0W+fSxGTQcaDcZQSuYSHCvsCaZZYN4OCN7Q9GU2c29jqOxTCul
q/JT6MMPl5CvMB7dUHo0jee1AzVMakbTEStM+8ASvo0BXcGJzOFCL57KUR7tmY/H
CZljiPeREpnC8Zf7/lQP1RQmMSjPCVSspsZK40OANGM3hGF/CMdApz3xDNkmC6ht
M4RSEoONcgRCacvkweKnYsKgh4QCHYaa02QDpURHiU9Zr91Piek7aoQgYQZ1yf14
EOVhf8its4H0PUW+5+WOenNsI7krPap0vGCJqKpMZekxey5OipMkghbjuLxEaFEk
jDRrxMqTmGib6KZ9ezTctd3qaGQCgZnnCcF6u+zJCr1VObj5mQaljXhiHshMTJv8
6ph3aX7JwgzvXP5+zZMNZdcmlcOLu9eTn5dodhX2GIGCCTGIZhLlxmCBOBfEjnLO
9axd32K5Fwkqsnfc38M1qubROdx2Emrfnln9iLk3luingFsZoKP9Hz6rdpCA54l8
BJsOeLBUS1ZZkeVjEmCF4mIESepn1uKu6feEwMWenm8vMUCbTrEo+LIvKDI57jMZ
fmiSEjatzjJB4uUYyAdFblRX0tplJ3L+h8TZAXJQWsyoiKkN7AbJFqMkEU/XyoD6
Z+00Dq6/Tozyhoh+D48E8zcAv2PdpD2+SWI82pTuAHWZ08F7CIBHAkYEWHC1G58X
fwHZJYaHakIqxR4cXFnHqi0avcJntcsGL0NF/5Hu9Bz0Vtkqx9uQ4tFAWxKL7Nlg
KCP2JC/j6IMs/9bMMsNzDiMow7ZsHR7HpIIvjL/xgMQ+Njf9aHVhHgrz5isiaSVd
bXww+jkjzlmRe7UC6EcmnPwYm7fU2NhY0l8/MUFIwcZf0rTsflxGVfA2tfwecRT0
O/5v0eEoTpUTvRH+ZZc6+Y67JP69nkMN3S/x1/hD7pZiXsjbJIIMwlXPPBJsllvj
SeCvTboX5tRMPCsSo8Q+MmnvJNS6rBjn5cCMV+nAh4hlNc30O3n62eUbX7WswzV4
GHSCBZhbJ4juP/bYAlxE2juxfaIqVRX1GacuXGXaE0j/H0gHZEeXm3mA70S2Nm/B
vb7s6CrC12XQlqCM+FibNvfRbPyKgjw/FJNTbtV0lvB0UDm3r0q6mXZM5AP/pu/z
O5WI/xhFWzhXWopHWD0mp+fMn6wZ6IksWQB2KA2oPHQBiLPJGx4zSeBSMEcJ8MIY
0I7k/fH8dRzOv26kZNu3/cDCfVa4V9KDXfB6IchXtWNcscDLicfU+p4SdJqg5CLp
bwZZrM2x1Z4wAeoZ/nGj/rQVr0nVmgZYDUiaBMaiFvAHxqSG02FcARL/cjS3Y/nc
eg8PBsavwhnjaX0JhfsfPc4gIM/Mm8lHZ7laF2LkJcVisCaDicetEsOJirmevwG8
8/9n5U+sEdeu3rbKo1nZpA1fhaqWAoWg0TKD463tDwIuhaMSx8TZk3Cn4H49R4Hn
UcHx/ujK6CjuwiiiJVc4FZ4r3xC6H6wOpvxo/njxDjHlZY9HTUZPR0ZO1rE373BY
ffqeGPIbRMhhv67QDw+62O9xJMFo+yPDgomX4YebVFv41ZVrEmMFPSjzWC/w1mOZ
wtDGRl94ZuuXEFg+g7Nf7pS+zk5eUWAg8EKImV0zIW89+L0ggWpJKSSQ3vE/hdx0
vuy/hQR3lHgT+r5CB5Mv4QhsouG1cIzIVvqzxtpblUsv9/PLUOqR8IUSmRJhZihJ
u1tcKSyXYuXvu+CCmfH5H4AwQ7nxXpDNyzBmDr6Au6b+c0evPoA2FWLpIt2ZNf75
53zLY5+5hsdYR52XaC1BaaU3MzX4BPCzHVXLWxCYywh9m4ND017vJCQHs8pduIBd
/X6TL1MdVUNT2tc9gi/QoW0EHVJkXeikEz+xuE5UXjcjk2qISjHxkfyO88JC+WZ/
KD6MqT8Hc0C1ZrdgGBlxuhpviMsvOQOT2hbJp+ZXQfA+SV9VFKSWwIxlg20TVN+S
kGI+pIgAD9W5PzWCj9+4nr6dSLyLsyoULLZz1MYuJqBN9und6whjlGxyACwCzNQ4
Nl6xq5NbfDXEydxCqC4yBTqFhQsCZoRjOpWmOjjrIpQDmqsVtzD+57SxFqFrACAa
9bT81lOA72eX00/11s3tK0Wna5TaaE1nETEENX3wg7T9VSmHC0Z4NMGE4NxacaWd
6kycHWru0m7R3OJRu1h4Fy3xxEZQlpfqcNQs3EUHhBm9riWB+CA3Pe67TT4AFw7d
NI+9DAtVbGocEP5ebOVcRh6aOdftFzUyo+wLf/YgcRBTnALLj0KUVMYRvIhMriLb
o63cFyFdRAD0h2eVojX87ru+se20fbrYTm+OfjntvifnULZkxXf+PnIcPjloiPMP
EFxk0a6WuckmN2wP6/DUfcoAM9O6KyCwqDR50aPXbkzLfzVRzGyvEcNRnDBDeuto
mtG21qhhuMyorOn026YS4ZiBFvzEBJ6rHRpu9aMVtdaB1faBoUA068Ur9L5curdr
sLKY0aCF47+LJW9UDMZrLAIqhUDcRBwIiQ0GGV67rCCZWgyBVI2D8vBrlFpSEpLV
+Fxm03Bnn1VLRkTgfRf9XPA03b8pJZx8TSvTkU/vI4oqw1R3VGPjOYalnmVzTEnJ
BVwR4cplFy42vzm7Ud9QNQgi0riMJxPR6E3A98+LXCawkqlP/6SVrGQwHZNvdThp
sesKSJ62Pbb908hliI1RZ8w1wt3Mx6Zm7OmyDf1Bi0PXVLpe67fGckjxk/1nm3kE
vZSmzzidh/iMwWElY+JVd06w0Fy4kEV2eUura8oavCWqMCzvxWOjpUqMF/ayRVaD
AfJgTXLIMqHj+Gg3OFlewkV48jHXN+nBbogZSw8mlHOUhpIaokrtA9DybAuDGGQ4
C8xlSD0uqCZbT/CAsRSFxZf5Zx+uiF1jM30wJFRjO2hqyltLnEviU5++IL6WcBOi
mfxM2SqoqxeOLx8zAAA4ilrL/bXR55AVRk75LDBhp9Eo+I7rMR7dNqahEQImd15O
Tk0klkqE8TQWmTUzlYCfTbpeku5bDq17jReDoEDLxsuuI5rSFVE7e1Jfs7wWemfx
IiKOUpL4M2piw8EtkZxxFD85IbROPrFbpRXKAXIjGYNnMx14fiHqFIA52826n32S
z8Eg4munpshpInq3blv5IgnYnySfPpajKdtUi+LQRjYKJtblQ6pWOKR0rsxSs7sQ
BZIucLOXwgWyRXafiUEsAd3w7LfzAfsHTTRCiFZUnBAYEGAg8bA5NnPX3yqHUJZf
0IgaoPGh6rLPuaNUpykwtgAwSu/TIL2vV/53m94Mq9Pc6syKLAUGZ0et3Fhu99dq
8EIroDDRLmy8vr//EoY+dhBfneVryrPEO3oKWIWkh2vAeB88Q7BY63lzwde+H5x8
D//xTmufcxXu0sGB2uv2UdnlzO91BNLN6tL8IqCmjwyFf7oOHBtKkxAe/BFcQOTx
2rpFAkofczomfnVvMI49MzoNKkyOgU8jTdRUq2iX2VVDabrooj7MM6xZ2LlFUyLz
I7V7t33U01xUB+ucIkX65JtA8miHr6fwUJAd35UN+2mNKk7sL6T1/dwGiqspM62j
vgG5hwl3cCJ/uKXSpkTFtDSS+fsoECBjKdDH9TKzQvIhBPmZ8mXCWEVW/jegB6mP
Li2RpbM7nrcZHusBLjKH6+sZmFlZ/28QUNLoUNdYhqyvKXh56aYpO8bBiuBZIIR7
yKY/A3zFb8tbzGvKizpA/tP0VbESq6Q8BEU5LTvC5FYAd2CajYaicvbBWrT1fCCy
kjazwOYwyzBnXLfoMwjo/8G8oqlpFOR9fKXLAcZDbesoL/Xo/v7HZuLMnPLYZiV/
SPioCbFHvJEIoJXBorKydmvfoCtzGh72OzwSsLecyLpSDcYaagEhopiil7QSblM2
XyZ6JUFvluCKSDn7cLpRIE0xp3PbQC0y6a4HlLLpZ56JZjfveiCF+DDH9+HBtyAl
CYkmUDCfo4uAIha5qzXtSDX6oH9Y88PpgKhx4DIUrjOFbo3Yd7UFyQ6Fw4gb8VuM
lSV5WqiuF93kpp89ZtqIjvLmv3HVUjrj3ckAx5bzpE10DP20JH4G9G4bZtx6Ju6U
0pHmxxcInYfpQolEzU/TgLI2Edl1P7M+ulX2UsIUXRf+ERwZL+kzeS6DGGTdQzDb
4trQAH2TytNjRS9BKy9G11Wc6xf5U7ADadApYRYepBSY0ZE9zFiqc3Aj+2iLTV6A
VLZ2iiHO2HE70zIFQQ8wWwNZU2wgP47onN8xOJc3IGiFJnTup7kLeX4V7y57nRjK
UiKN47HZcdH9IgGkvvPP3IlWnkkT3BQ7UAHMtMUmUL3oUr+7E2VVl2mxquphODFi
bknbEz5VcIXz6IbvRzV8ebo9tArExEigun1FszDWERk7bMEsXNI+wDJBxdASpavl
fmkS1gk8b+GrAgzbudwWG3RlHVqvvl9mt0egBmR2HsimfrFcPv9z69DOiy+DuvRC
GGMcNF3JpmU1d+OyzNkEXJNRC739FzbW3Kjw3UxP51CeTXZWs+kc/IAcfP6NX6hC
yHVhiLHKlCy8UlTfydp3VdBQlgzoFNaK79XN5pnkxbSxxkbNqgqOlBiPv1e+VUtr
mo9ybVGBEBThq12S/KNelkJbjWTCstmFp4xsn6B1jAb6ti7Zrw3ABlBb6ZNroi5W
VFyJmzCH/kwUnC3BeFnGnX84l95gmFqlI9FWLOmv+YiluNXeq+Z30LlxJbcWwIxM
NPXySsFGTgdMX20Au5C05WEm3WHKjv7cYMjCDch636sVBAzTRkOcX3LJcBSQn/BQ
tLU9Cid9cC+S/aIqLY9/soYxvioFmb5U/g9wyEN31LZY6Cu4P0x0Gs9PCYhG4ZA/
+nHaMm62iV1YhlCytohe9NHlhltsBklIMa4ENJHQzt/Z94goy5/8xGQLTV0Qc/Z8
9C5Q3dEg2Pc6x7zuoYMZwSvA+GzXgFfmpKurlZtY+q2EeOwfN8jK4K8Or4FW59ba
QoP8ZeZRNSZt9KsYjXyE8ZkmvUKux8MZdcVVBvzWhi8TGOkQdGFDvpI0YXuY8RAH
iTRxcYYgGqch+6rHDkv5SF2ca07GjetAVa6qhcZZa4vsZol+rZ1iqzNs2kk+nYbM
HGvfx67DQRz2cDWlRBqyckM6Vy5evYWQ9iWWMfHtkFU1ZvdiSmMz9DtL7TGs2vKB
rRpZjAF0BAi9AdwjVMYIdOQ9RkcExC3+35xf0NNSrTuKmpmw5laJQ9dwFWZX+F/j
U4/uxGoXm0wbtpwGMUOgGOD0yUnvs7gGlLtBJ4g7+fcYcuQRaYtYYpB5YXyMS+C/
chIC1aSACrrWH9JBopgNPs/aI2RyX4Ip+XWTwxkChUXmcmHxiowJHVHJkcW4+Hqg
tveqyd01IM+rV9K/YWD++RS2UAcb3nYstXagzkdBpMuuWSdE7XYfzJb7cju5gyok
p2k1IL883hZa6rrpuuL/Zg3N8HhWrmJKbCOxYNpvjssoonH5TgEmKIyugcDupmxj
6+iy0zzhTB3mrvvWlbllvwJ159pp+oWAWpKLrHy+YewfFTSTyERpDA5/X6CgU7uG
yIZrO7b85nu1DR80Bt5VxZXjlxAxmbq6BZVqVYeIEDeieprNcWV/+5o6dAXLHRet
Q48QFaxIW4INNHsdRrZQjtj0dMJq3J9tDyx+xGfzBRzQhW166iFjahTjucEtJvsE
3qA/UgOZ+5un05p4VSmLraw9CwMZ0tmAEk9kaKy8yFbCYtBsmutIyaECMQ8vDtZh
3l7rwbcu7i3pCGXdMektr17c/I0C63pTV0FRZGQcuTUAX7OqHiuzs9UH/HhdX4/K
keeR9/c9m56+5cOpczQswBIRZZKgWU3Vwgm1KRss2+kFfqP6OykFv6tNHpKwBIl9
U+9hIN/0QTCjsgylkoS8cUpRjXB6XtKaCITuJ9SPbmU6LYChfZ7GpBi7oLcD+mnW
U8ZrW0YYvc4EZHnS49UyiiX4vaIpShEBSd3cNHP+G6lupMIOXu6oBcYq7aHqfWhX
+/LryVuQZjZE6sE+6XGfXvv85pOo71g1tXmR4wNtgQLKrGMy94B0fwSYDzz6Xar7
T34F45cZK+SpxybaGgPtd/luLu10/GsYE517KbCq7ISEhoiFRG4XovTHfwsv3uOR
5/C+SrK6+XGOczBYSfRLmd46mH7a7zR0148ZBEDSlARrSUxiZojqQW0tNoWfdavC
eHYkHWC10cH16EOE4LN0lB8YZyA+uV8S6cIob967k0OlckFs8MZg3qzwcMCOwu9t
ENa1+Hy4JHiPSRvxYG9PKrPwRrGVXJuXsfkMJu3SgMLlcjG7MpoCH7YkPkGJ7qkA
VylWlD8bat9oSRmrvIlk3YeGQc9YBkONSpmoN/xAscNNU2PqExBUInJoK8vr1g2+
ldR/y4NiphD3UrCHM8JaR0mMsCwuLPmxpmPk4EDHt/dmNuIb0Y6n+r/C7ZKRQxEk
nLQkdNsg31SR29/zZbFWq5yJCA+VrhBbgNZZgtkZEiHauIHcRAmQsIvx7SrlzOjN
xce8vbzGlhtco6w7r/GKm6dBrjklDcjksYf0vv389LmhXw9CokFMNbdbTp89yXIs
g0sy7Ph2Fl9RsPB850CL59NkSrCdijn5XB8vo/rRzGogYeHVAqT88AMyUAlUg6qL
GCc8Og45NXs5EGpgzujB4ZAIPBYUIUFYyNFLUbywvE8x8VPCnrNiLlpACfG7VxBX
SqQ+pLi0Dtbxidz0n84l1YyuptmkIs9zBW2VBSQfCVHqEu8XKq1Zw8ELpg5XTltH
9dWh6aeLEFgPMynFUu9DXLMEMGDSu0DM/G9jLx7zW5guikCkO/HYDif8cTMgyl76
2Gt6vd1uTgfS1DuJRioLCqZa69Agxhd2lrVNQT95uGVFbN21hDFQCUtFIFGeKQ08
0rI59xe7teHw7GfFALnCTJb0xdVTILoNxE/SgjtDEvMl7+yyD0XnVq+Glpj6/jqM
fdvKJIKH9g2SPA75l4Ow1vN5lZykvqrA6s8Yks24c/LrfmqsctOiwS99VGPxYTG5
A2ERaVGvU2GrHeZfGVrvuFtizPdlgfK39bw4Onghzgc/h7CeH4NvlxxXczsCQ6MH
emkDi1Wrw3Fja5EyZWEDvShnOkdtbR06Yx57Slm3+sgpAj2zgY6uUEgVBICv8P/P
vZUpbMj78RemxNFL9RG8M5R+tZ7d1p65W8MnsucdhxHXI5xXVXeudB2w41SmWJ2S
rMoRewrICuOFW3ZIxxlqL8+xHT3EC3+VqCkuI88hRiVtmvbCJIbhQ737n2s7FaT6
CnptPydPfStdKmUIpep28ePegwfYEkX5aiE6z/0AV7Kw9GTcy+IuReFC+v/CsuMo
fzuM7P56qR19IMmswPsBelwvGlwrpZ9xtpw4unSIh3XfrpbQG3C1BieQsWAlCUug
AVMNr/0jJjALFSgv1nNyjHbQM3X+0PL+pjZstI68ghNn2I9VmBZYcd/nGBq1ieZ1
jAgSZ9H6NwrIJy4bEJvtPs7SFce8KaYImYAXN2iTlwc/lcYZ3kBNsH1d0XqFNpWY
SmJDwnhPC3qfbAMDr0FzmjLee9l7/mXor8S+SiB1sONqiXj7NWT+/raNizIadpOJ
HNbFjB8CYDd40anxN9wyt560YSbWolhKf+ItbVKbjmSWm4hYA4LfR7qLpgthoUCB
vKgw8Y+8ELsNpM+GLoOW8jf6RXrvCE4uYjUUP0j1mV3OpIS3DxH0U4dea7Pe8NWX
0mg1rMG+AtJAXi47nvlha5hxY8q6Uq5b/psjMQQf4Rs=
//pragma protect end_data_block
//pragma protect digest_block
zPouHssevdeof86Nbm53CzwmpUs=
//pragma protect end_digest_block
//pragma protect end_protected
