// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
RM+E+cpdxVnj1cY/heKlSjtYhI3mVpki25nOYi7vhftNcksk2mlk+1tW3dr3Qfghxsb9Chcohfzu
O5q6Y7I5d+2YXsw5XhyoI3Etrv/vVkWVpqOZm0SZIq1XF5e9Nf+zpHhtlhta6Ysq4CuYJHo4AsFF
U4U8u3wMEZe2VOMG8Mur7FH8fcPJHznUxSAG92Kk8IU6UpWAquUZQwZI27VOhq7u4D7hcTzf8TzR
bAXderp9KJFDWtWonzS/jxA2BVu++gCMwHLDW8ufdi5ATs3gFHh5DHDRCCLTKX/q3sieYokATilu
mTJ3p68An54JtRMV35+UvSm3oI4GZn7+gQxWdQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13456)
fI/xUNGH/6Xhf1XiAt1xZnpZEvVkl/JrUGxMWEBMsUng+h9TYKQhNtobfhuL2WBcnZKzRLo+iQYC
WLuQ7RFWaIcOo6ZB1dG7M0T67PCiwI6GdruQFwhE9SmxWJKLAIQlZiAzjGbzca2sN/MVKg2nYqVT
uRq4zKSq2uKOF3nYijoeKy8NhuB+ROGGwiZ+yd+F2UThdNksiDM30EdCVt/MQXWkKxSu+Yke9rJM
f5JX59/Jx7WG65EystUIp+4FQ54J0xzrdcsilahDhYFA719QaO+iuRHyyLSWWIjCndQ9RRuC4jG7
THkTAuFI7ck8re8kzaqLGGgqkW3rj1JyTOTCDdyim5HcEmJgeyyN7kXRsvIHeghlrg086t+S6g9K
kRBUFyXynf2JvMthRA5tymVevEwQ2ik+PdFDm8vGMzfKENrXXYTJUVxuxQlot4gCu5RrPTN8K7Zm
s7PserCbaLZ3kV0GL8L8Pm0EOKEQHQxgErMGENoJgK9i77lLnQDo9wtBp4/0G/c21r4tqWWa431x
1vYHPIz6jJQkCHwSFJvSuQ3gSixezwn2IMYVofOLP4zNmhqsbY9N7v64+RM97UbXYIP2FUwM21O7
Yr7Gym+2ccVBiUNa9HEuuYw4JT23fi4IszREGrDpQ4XqMIDJ+6Y+hTtcys0rUfQHLauvybs3ncLf
ZrQ3QO2rJXRbqu778iwK22M8kHT5QOOQ7qJc+O3PSbLHq+8W+Nq70plVnIvJ+Of6EE8k5fUg1f0M
T5ncDbhIrNf5VLcCnM0MNIF7cL//3sci1X78DlUONhcUUw5fd/ZxvUQd+aT58P6kO6iYQc/fIOvQ
NpXcaT7vMqoY+6By44sPeZKOsSqjVoaEpDtVKar9gm2zZPZ4xq9e4nu2x2iibeEmT2SKDTSLculM
AIoCfYy3JceYEgmD1UiSIelnZ2NdzIvAnYxmA3+DDFz/Wf8KnLoaegzGLQGgA/bCCnUyiCDEfW2S
/+knkvPsySk976e2fyt45TsjDpzZo5uZDezjf9ObOmguB5Lz6q7d6Jr3t/z3tJW5Qzrp2fy0PvXN
Jn45OTP0Uw/QeXZKiObPDFyTZQ3A0RNWW0hCOhkgetCE64FsJT0RjOgdY8bt43w0iPvjG2Xcb2cx
8qUP2zhyzqSav/DxJvUMxYrFgktOL329+5wznVGFhl1YxGCEThrlDGjY9aF+AzEYajMQAv6UcKWT
DefKdxDDLbqShY0Gs3S+IqonjW26vD5mePvfan05Bh+9uAjZt423oiHOXkjOBtSIHWyJ+VJdAOOE
q7qhCoUcRREGfIwaAyPAYO1MJF3OgHLPpIt/Pq8DyIlcyYDSJM+CQqDpySKi0qs16/P1SymSkhKl
iOJDQq5ggEMnqMIUx3NcT0dUnnGc190+oLWgcrm529Wb7mb2pISBBRImL2eqMi++7ieqXOv3yfcB
/Fait9s5J13M/wI/mrdIS93WD/FNKI79M1XMZDATozulb4/6M1ja4eeTWp/yfcF+3C0EdnzHZ5DU
B5Z1Pg+DxTKCxw4DFIXTGiZB0y1A/8gy8o7J6yxoRoDsB0AfcUuQBK7uU037kVdTv+Rf4gM37lO/
afRZa9e4MYD/P962fUU28ZsC/QXNe6GFrqux/e71u/XYqbxSNkwgc3yrzx6OgS1op2Olbrh7T/Pi
Eist+roBVg8M8LQD+OoCE3BcdebtGVN9busSqpJhB690/hhuOV0d2HuqZB8qgiUWz+2pgkHasP6A
1xuIXjuF3MAW8+PuXVzVQniv2eM+gloMii8VXtRm9NK0X9PoxQ7ZR+/daGdCZWLdb80AuvMCi8tL
wZGDoEvzWuo7pc5hNnqfwPX8+h86hVBQMzngZY8pTmmED/hs/HgS1MbF7UU/4yP+bDBhHQxkZWpt
Q+U05YOn3nxe5djxHP0UMDKcB69Rn5Wm8VZtyihd6YPgFX92EbnEt7eAfW/8EzrwpnbFPNr332rx
NKskJC5Mxg6Hm0TcxFGZKubI83bF32YqoN3qpVN2LLmg571cdTbjTDjykStbr0r80wytu62NA72H
UbSCQ0oPI5gaao/FjAKXdpPVPzCRmfVlAUcsllnBNh/yY1z5cs9jifpsqun0ehyZXSjJhULlAE20
JdnDeKEW5ECwbzAY5e1wrdTsE9MECxJ9Wt2crZa7QAufbYDI8h4IXewOH+lKNObZ3mHeAHnBGd69
9fDc5DZMfC0wT/uB+c2FMJAd190KttkT31C3t8MiJzNMAeHCemwXHe+TxL4+pLsVC3NWxGluIHah
huR1iTrW92mGDzFABzGFqfTd5oOMFFajiy5Os8vSY0xUe90U1puz8hB/ociZWgDeExmCfclEWlZJ
wyA9pzR+9ilFZULeTD2tXJoOStm0DV4QhFDcmNarKrmNOrvDPwqGaH+AkC6Adw1EK146FrISepys
Sq4woghYtUEajoE52PU6szKVXUADcqH6B25EETuZaklXwZX65KF6NphEG7RNI0e0f5NeFO5bIz99
zoNdFdBaaXDEi69ozfw0P/7W8R5Hjaz/7a6no3xSEhHvGHkE8IstOOkjQcZatdWjfVHiLzV1cJ3P
CQUNT0MvvoTTGKWBtYKGHpNWgb7xCv0ZlxNyrdImOVbWU+pkgXUzM2RXFAYQkNdG4p+BU9VFAV9D
Do5n5EpKhbEFAdE+UnaN1X8f1JfQcTweGbbSsvfzHIKc42HykBtLxLPZAAmynwctx3eVg1O6yiW0
tK3alz69ecSzRCfXM3cfOVvkiy3wjm/RGfGwugxDtDCKKvDDtH7p8e165YyZ47HWB5C1pXH4l2/0
KzouU+w9VyhSHwrMsGuZYfXuo0ZT9dWboJzv3Kimgdq7WBCWPSvjQk/58/6IQYdohNjy+GdIQE14
jrzbkKWiZEMh9duhx0sjkCSrA6PiQ8otAzEhSFOSC4fGS1AwIX6CY9oWF5naq48B/vfZmdu55De4
iTXZNf7NQwCkfNzWVC28YniHG3V0D4ynNjNY2tvuyTRPc2jNh0GQGWO3vAXA5O7norycrfq1JfDl
04BfIc/FbBKGelf2LHh5PAaBxSJNIkI2/n/hG7Rba3eGXElERiNkt1FsgHu4zUSR/0qUo0MZBiET
//ZF7RB8klqb89C2P+GuiNTv8Fe6LIH3rqsZArTMm3mnWeZ5OaGnRQkBcKg0Lic7YAkdh11xOkoL
3WLvzHMvtHZE2WouTu/oyx+OMknJ0LubU0CAlqUvF9jH3AaU/XTZgqkTcCmcTwEGo/GHThuBU6Re
LQb08VxqOQl9OQDaWoIin/S+Z3HzZt7j5bU8dK2KaE+lMRfTfTXjM5hYKiL8y03uTi/y6VuXfF2B
cNPyeuScWTe1c+iH1EOA8/VewSj1nV2Y66pt+wo3bTrssxEotpb+hj2H07w0g4sHNBSbwfarCkRI
atBv+xTIoRv5e4XWb63JTcLK7OTcMLN1vxL3+5yxVAl3Yuq7jMszTsQDgkalwueGsC37OEyVx889
AKKamRSh09CXsQn7l2RCaXoqdlXfm/+3KE/jXnwOBsyTz0NUFPD9bOT2azSv9tCTAZA0GaXKtq9P
IklQn/qysAfkAmlXXyqPSLBkq85LmdxT8L3/13nl1U24Y4yT5eeJztDorDbLsilMj7SdPwI+iUeO
5HoB+WxupWJFcqJJ594g2Lwxp/Mxrg2JeZlgTejyevvnlaS2y7All5bmUi2G8KeuXWNrX4F5R90x
68oZ0+sWx2T/AbsY/BGAEhtRu4Snt6y104jJr3yfHMjXf5A3DPuyNXEj1H1kkZFC30gv07djHcZE
vV8z6aZhWDdosdwKJ8dKAIXF8en5SMuAxhbru7e5/UdHm5k+9KTxQ9fXlIDeovBBitsP2Owc3wTd
GjgnEse1zs+33sv2FJJQCF5WDMcr8PpyCPvwTXE2OiIDy4mqcX0tykmVRQqEybx9jsQzgM1Wzlv2
L+yvWN7tT/ubireR+eIoXPK5jq9fhTHqfKCufqi5g7OPnpYqbnZtvHVSKSPDov0R7fBF4ReJIGYt
j4wl2M7L87UoKw8rvTZMRyo00nDgmlHVM1ijKHyg75ZGh+DbGFVcmr3Ka+kUB2PlPDpLk8Uz9ReC
hAVv0l3W0tX5O3UL+siYK3/ipaAI9Pqdg7KhsI5JmYFSzdeu5YP3CMkbRr3lcLeJriAFxocN5zE8
D4kn4xd5YOL1G4eus74rsH6dJhQPShOo5trTa1QmjhkXqesabGP1/1fb3GT/N2KaqEdedbU/pb49
s3m+d7n6edHrQz+RRyaR0AwvVFf+usMY7vxGo+FEgfq6o5XclMRXJGpjmmI1Nr8MG8rD6e99UL9P
gDiyOhWUIJEgbPGmydWGFzLAUUpUBwXMNj+0DRAM43Yiuf7Np75ORRga2BCL1z99Xquk+qXczCuv
Jv/JKnD/gV3IyDckcarlkOiGV3hBp58LXfYaVcqzUIYC4jeSmZDB4VAUHmlwkuQ6M1Zo0RrbWFcN
vtrB150rJA23D8hyW2G7O1kV/lYTK9ayEO70mkBZJS0ojRWeTinq5UAh9rZGUBmjrxxsDYwYGHnj
RqKPW1ePNejQpU8W0dHlnmG+06udjWBYKUmLUZyLOoodgsdgzNG0MBKJeEGG1Iktej+YfEpqBMfC
lqqhT8u1lz53uk7b0GvlwE9OSM/+0l3zfvHNXqOk5dFuFNQX2/OCT9RNO3exCe4Eig6KCfQRrlnl
n2HAr24m0hQwnq6WSVIpen9xcRBi8xykk8S2GIcVMeHVNv2gRR6GtO6oJ/saEvrpwxn8ASwvZ5Sw
CoJi0UjPNQ15lBYMcXrJgpSzK5EbAvAnWrKIWG2tRUCTMk48aa0c3dc76mU3P9g643PbOqWebKmg
/v+cy4C3eM2cwo5iOwqCrT2AUZfrB2SXwI6BQiWVjLiRqE1oHTopx6aSw2Vxg4smXIVwHsToNnZV
cO7+DRYQ6vrswbXVipp/paLR99OkEeCc6gxaQaqU6ClJdcyxEyk/N3/rGNatIsuGdCqdIXIhGXqA
rpLsQUx31WXXlLex387yf8rqhsHt3ruxf47A2JyPOIhfUBqwosaU0t7IEFAXy5JG0anGLZE6cvmP
v6Ci1ER4TRmeFk5JiWpisI8B+z1qgLvNQJDGSPFVhPTildgPvnflAxt8AL5MR6XZLb5UgwW4U/wx
x/Q3PTCHj3iQhdcNdylUvelrxvVIIScMUGBfFxhMP9PQfkfdf/BE9y2ZnDGUyKuzV7ajU4HRBnEK
RMfZkxV4rA4YxhUlOgQRKCCSh6v6wwsIsyIYbRBLMbCS4MZpL6IWPrMbrOG+Xh0umUDd3VFIvsL3
kyBwzgcmHdxj+P+wwxlyywvegUbja17DkXCmKQ4FV94UisbyQWtQoSBXt5AcK1B88vRbPS2o9kBw
fw+hcZByPwhmSWHgTdqwQcfoalwjCMuJSiklVoPX+thOmkrlIW8FmYW2bjJ/V0n3FVErsJK4aZCc
ZJUt4u28Qw1z6O/o45Z0DTxh1J7oRX8EwNCQTjgUkODcUWEolxoGIyFo5cCHauV+cdFrh7TkURe/
fXsGpETnaAmdwWHiXQ47y4vBWQUnT1n76rlgRY8h/0GMgrbdlcAFtNErgYjfZBCNyFlzy8EJkG82
ismPTdMYkA2nd93ASFMA+6FttG2/+BalEft4OSNgJwHfjqO38zAX8/u7mQfkSFGolMUPq1NFQa9c
yxPDSLxSYiJL5zgNRa3Di8JjYGBNEMCQ7uf20jP4KSa+2mS3VmoOzDmCX0sgqEAbISbHVxsnKZy6
GItGYJnSyQwVgrb0DwCVYZvWqAnYpqGMw6AAP6Hs4Bg6ruL+FvPcfEumh6WchdQ3se6X1dxWq758
60EGIiUzQsMXZXBwdD/9lxLA+olze3A+e6voDKTMcWrIPo1OXKSNig3bThNKNP0Bs21xbfY8KHv1
sok8pgD0qIDaTDJHPbS6xCFZzAn8bKZHeEMjIUb4rgCLp6sNLuk2t75V8qZilSPSEzrUYlovA1Vg
32ik0SgxwyswIpmQcX/c2p+8Urniv22Pef2Otfrk8bVYAbKQXdKQfd0w+qHmjwjQLlXT7jwecxN1
xgcQVZKZcPMqx2bmuCmaporwOg9twY1S5+uQQ+JOPo6geKsOEVLF4Iw/aZiRY+wjtSaB2/+8YmIc
Mi5rKwXsOAO2jDDXwtnG/Uk8ku8LtnAZO/gSMmXSYiA60nFYOXyzP/titDJm4bsfJ9GdFeO9L/DX
7NGupla3KiIPpeDhG9HDLWgWsPu0CTG6i+yBhcjYN8IB/44GZPZTjzQrLVev8DDkgST0F2oQMLG0
yV9yX3XAb74mW2MTh/+hU9RNa6c2lIcA+YbgcnN7+2678mdVNV3idzP2G3sGcbEMoKr45MowLG64
BOSfyHJ2PrPGOPhwlMek/dcI/7Sg1YpVjAEt5obIMl1xSdMdws04EZ9icFx19DVDuAdyDeaHJ13x
cUDlaBUrbL0ZgqQ3i3oTf5GhTfdEFZ2NJXFC2WXln0UBQXAFLcvkXr35ohQ+ENpfvyO80W14JB+c
fKWQ3YvHmDhZhDj1Icsycpfj4yEfS9K3M9IvNS4O2hbu8CVQZ/nSwxB9P5d6FJyKK2HFRxxsvzbo
pcH1/7odRCqQyHMty+i1+1jkJP6n4iI/809lKQfVpS8YM2C05/NoTsfnWwnoRtpfXkb/eu0iaF/6
k6YW26ej+deL1i3kK7EaDIvvp2DyypvJL/JnBYM+uyuPaAtuin+630X/UR4q3Us08CA+ktFfHvev
ud0y/le8dL1cyPlqYnxJF2oX9U7nRQjIVdrKvOA+S2nW8LOitHocXcwTHj6XDGBy/mptFolr6MOQ
GIQElcBFNlSzpBwXGPMua7kv3qu15NPmr17++91BkocV95XyPC38/b4sQAnjt3+fxRxm8EfMGFLp
m00frN2tjEvWZbl+IgPfmITnQHowWVA3IeheCC4GOSoeqdk50jkSENOhD5YbG6XORz9wEmd1dwBt
K1pD86v6/mw8wNTm5mGpaxupQA270ypiTMxbl6we7hMHBOjQV2eZ1BcbK/IRlQytV/Mnp28GTgeK
tsfvEmCGaHOkauTp7pNKQWniEUqIJS6SG9VOzlSl5ot2y/y8DLQb2bLiuq5FeZryd8OdDSmX+/US
wkpUqBRORmbyZ+dzHGFVYQJRhj1g/no6Zh1NPG+kDCyTdJM/EMKf3d4Ev69Wjw+WBSSmmSQ7eoc7
UtsOffwLrRrVIXe3E+e7H9CNd1AuF0wu5utAZupmv66iN+7ZkuxaaZ77AnrdF/1vK2Ti0QRTYzKW
z5y4g21jkjt9Q+yoEyHMX0+PQyW9XWjeN1U1Uz+SJnKCGyqzr4FsJw2Kqx0SBZs3OHZ8/y3ItwUt
p2hl8Ktg8I9uMWXolnkHaXjIq5N9UbHlWHgxUvCHHclKB5FyRTNEkH+h61mVWJu6weqRcAITdCcg
2imZOlAV/RIrBvBzGadI+MTJIYXsbfjkn7QWTydFxxj1NyFqqwm2DVrg1GUrQKmwdsLlCFzGxW9v
HPsL5CKy+7+33Ee7vY1lrg1kDxJp8rTPxe1eVAfML63CRugSPyfKERQEAPsw1N4K6iFCx/0MiMKE
lwfk5bYKinysdHy25u2E7zDM3RvLGDrkVXv6z49+yvg7S5UeVcDdKXknjHvMUFtcd8kOZjXsgmvT
N5DjRkODWFxBIudhWgmXj2fJ5ZlCTozrexKSpCLgtIlRQ9mmDi91OZR/qIRAw/tgghtqEABgj0hk
wpB8ouGcPeX3JRh8xR88mKo5W87B8z0iv7L/cI9Ijz82AUWq+Xw/YlGWk/zBn36tDC84fMIo6kAF
gyS/EeUOJcvT1ZaFDz3stCYGkVzPgRKCvt23AM78+2DwIQhVdOrpkn4Lvbc2GikduMtGTXRIz/WS
goJPfHQ7HFMFgKte6TQacNsZxpPSwrKQ46w67qHTEqY63B3JgKO9j4QR7jYwfcXp4gsGdbRUyPcD
gAHxcAPwcMn7dqO49wqxbq+siWsOwL2lBp70v27igfjOXvKQx33P1CCk6fCMRrs5QpB5KsE/aHWP
Elb467roks4kehp/dV2BKuiH0bKi/iapVpv7WVCUsDYI4OyWJKJSNO7aZ3TMLgLUDSfjk533QonT
CAnR91KcU5Qz6IqFEYy3ZGjNMqkJNjJ3gqkYVWd7J+HcV5286FFaqejfQePac5hyDrr1TFwBxw3k
KOWOzUwV6hZREdu6SIyRGrDyqvh82JSg/GrhWipshossqfrILWg4rW5iiD3+14AqqPOANgto0h4S
sk43kDvJVRV/Abne3ca/zrce2uAzacNA3cssuuR79K04U3JTYR6eSQq959HGJQknohJ8hjulH1W4
Y3pl5ueJrqvfpbm6xSg7c3PslbV3xJZCQYEVvGr9tRvHGC0k/hoCWpzej/psJhtOP+Flkgi0W1Kk
4R06H675ht/DZbf73UH/KgLMKHxoomhTa4ZMsC9SJNaFmJGhx3Fp03T4Rdfr2FIVUw9hwmFdDREV
EgH7m3s8pE1VOl34LeCjiQDkCpswSpuDrk54R1lQSIKJ29rGcFN9aUkFx4077M/Qf1iJg00DEuNf
8Fla+Nef2K2wkSuIrij4uSuXaT7IXoWxegxvnVJi+l5FkLFddiCFH4f1jje6gFL0MBii6uzzTH3e
5DLsn3JyGdFs4zQ/lkeEsjmuCbP3qOfSnBqVxtGZ2PUtIv5XvgzzNEJ4TbPCdhijfjEz6ftxduNL
sJ1Rf+9BHxc5oJJo/CUg5FExhqHSSITMbu+aUwvYGuz5ag/WeM0nNS6uOsj3NPJ3M6o2yamB9bZw
76ORjbH0NGl07P3SIYtjxNxWeBFqt76gXpoarwICvdPpaEh0F8yBhihjSqsCpVjtsF0xOBpe2A37
0LiesCy/HFne78jCB6bJL8GVwggudPJ2N9W/dV46CbLFywFk/zrPka0aUvcyY0Hcl6Gs6/756/6Y
+vQjtqadAqMhJ4acQq/whI+vkzn8EFogo+SA+6jp1gvPOq4p46qHsWDUi3V7dAHnUPmy6EMc4Zw+
hlmyqefDlXHS84R1tyQZWna2FP1+7EK0w5wZHWsvsQUZkrWoYBNgwIH75/M/WHAeKowxd1HJ4+HE
ax5Kd2KSXWm+4srTuIFPYjscId1AThtFL7WnxG4i2bemzErCibU5zkBf3B8/tIBCJw+PxCPwSI63
DaTkBQcIIeYcYYFx0lSoiUtv5FuUZkCU/Y6/h6rMRgIFS7S2V5DiM6ru8aGub9v1Q5LxEdfzC/DI
eIy1UoCB6Lifz02gq3RiMfMDZppWbPuzZlqPH6dz1npmp2iEEN+giKH/zmMqYqOTzxrT0o4HDP1L
97DzF3HXUEWB0bfU9yH/bBJzoPBTkjS4z9sqOM162kGO7EYw+uPCe+76iWZYXGJKNySsqs+MTXTk
7LTsVM/N1LYdjMfIA98RCEWELbFIFFo+GLFASb4KuCTTNqYCqFfc4zvyzCLERLwVnpExO0NdTGyM
70qUqSdjV2gJngIw9TkEmMOCPdEYGFOGoFALNhg4ZGVjsFYPIaHITmmBcYoUu+BvLzIj3C5RumyQ
ct8N+F+QEg87IDbQdoEARdDZK8USczUyYC+Ojy2PtXpc3vUf66JCy0NU9Oie0+uAhu4rHbkkcj26
VcA+s088Wi3BSo14hZXmuD2HXRqoH0bJgOdGZHzF297cq/H2K5Asi8xZZ38bTzSes1f0FuSOIwT8
NHvuWUtvxwCBBVm/IcEceh2KSHBjC1ER+hUtN+INstyfLlbhQQ2y9GYd4p/QOUannukCjESfUw1e
hWN2edVcoE9XGkLpZQ+apsbVuPIpIwotodQypJh6KgCIKwGPByQ+3IkqeKML80vfYtMHaYU4SD7X
fCrPg59GE3wik5kXF0dTOLjRQtDVyhgW/DORXsgCeDVWQFCt6fiQ/0/h+U2bWZ7BuGtx+cU5tyuC
GNcisF2WaOFejTT9YODygt/aBhs2UBE2u/vEI9K0MywjHQQbwvd3bUfyFVIG7PD5YWRIf8Ge1pBr
PBVGJOzOwcZc++QbZf8z8siGkrvZGtlekzc3JbvU1JiPgx1YIOolSn+xF0XZUA0dkwXA/sOTr0b3
TBeV8g4T4gIKKoZzK9AN31B2qur0EP32cQx3RvVObe80iGGzdxseyq4xr19whhbS/NF3PAbU+Xho
qQqJlqaYF1C1t4xSohWQl4y2XlyCtdyTx0p+2UIkd2OmAYJoopMPK+VLMTkFKMSWmLk2mt3F2eJb
L4tSoqqtmiRHw6tt4lasWR7uitIg3BE5/73LorR/e3b4A8qpaTtmCl7yri7hwoPhAfSNV5HT67oz
7dkaH/uC0CWonWgq56EoQJa7j+uIDiqrL3I0EEHielm6ChQOxFB6ARiiuk4i1GT8dBhCVnNs4V56
cSmOQlCGKON//H5aMGagxpYpj5daku0E/HlyzwaQW9WcYp2TkacKLKULrtawaWIsbCN5E3w54KoI
LobbMKvx2NHRDn1K7m69URNDapnN1QO7f/GWATRyej46cY6duYxjid7l+gTEzL/OP7ovNNMa6DUT
onSOPcz6HEI+hRa3RT9wHPGSqOKDylRDyG1KVMp4MDrF7NUEKndo2VRW8MH36BO2j0Ouw9JiAS7O
CsyZgMz24wCdL3kT5UNyc3kO0I7pGNMd5KyrQO6Bd1ZFZRjT4pEJ5qhid3CoI8wK0jfXuU1SvRc+
uMPWNADa84wzcHjk8XY4iTF7E2V9viLen37l8ZihKnOH+eRAcMpww6n07JkZExrb5Ebo6Ffmz3Ny
HwI7hqi/X4qYoz+lsFePt71oujygmv2/zUCIwmu0QIxNQ2n57GXt+SGaUwZAKgVu1H6ZrnemV+Rl
HPN2XBNopcRQBRt0q9+L576p6eknpYUIoRAe37S9wDp68eyiaR7J+RB5WHdquU8xBScipdtBU9Qe
TNPOq3lAh0A+hWVxyb30xt7Mt118eMFKnxewIKcMzGZE32uj6ChqjX2RyexE4GldIy+hS2vowSSM
tto06abJRy2E0VMCkwQlGIdEtLJ3Nn26gUhKKCpmJ9KkvTIriHpA7SXxmcNuBUUgKy2A+301Dj76
SEdFgg7ZwFKAeNUcSvpnjof8v3BO+YqPa6t4lA7r1l2c2BuFp/abZgISgm8EzwqswkkOdNFNHH1a
ErOsoWDhN2f77piB9+BTTE6Ytre2Yp69HjmeEzLS4SHLRJiteGT0p9NEC8vjGh07TYnGcOsNp/Q/
T9VX9phwaR9jWCFA7kiDg6OfUaAo2yxd+Vbmq4Jk24ophyrgObJhF0M2IAqLHov8WtrowI2vwZtT
+SslfMgK4C9DPT7Dqk5SyhXidt8sNUBmPlz1nVDiKeHMfxg9U75+0trSszX4c/8usSv03vaexJp1
ZOjdKkwmJPrm0TIwdTzXlaYNx435BbDV4uADLdT2Sjyn5fvDvgBaolOrm4xitDWUlBB4ZqF5iczI
UcGTaUdvOV8+vowFXFNHjpTLHSIYsw4ZoDCmvGJMgIKRw+qNJDfrbubEFyYviiepC+xAMCXFUYBV
vwOlTrn+2W6aWcwbxlM+uv0EtpyUn4O8+yMrwwLApC2oOIOlx+gP2/U9CqH/tllGuNw7bEQgzRsm
sgAeIuMwGp9Ex6205lfQ6t2F/JZ0x3+xKtKPE51dkMLj/LCnNfFFLWtqTNgEQ1bzJrTUKKUv9yOb
M2K+Yv7MfEh5UXp/zYWN3mo363OefGucVSUSLsyqtGfFxoI7jN/9kPkESpww7JCXiUiBySyNgfQs
lKLwx6M4L90/filAuPrv3Tp4Wf5+psxl3yVsZbd20TUmt5ZlGYKwy79hjb3iUPBbXNMA3jILD0tP
IqLznzi/ffpfm8HbjFYEBbNhjZpFduYF0qXCAmUwLw81aATEXLTTpFBCwhxQzkilqvnyUPRNsuTn
MGEkOko0yjf0W0P7+hhwJeGhsUBHCrc8z9U4adRVZfvCayzzEvIse4IWOvtTNiaIGCSaO0RmaJGX
G++gXMOJKybRT8+cFzCOMekYzvHySGNkPqj+Exge48Gh9RE6qOdQjaLD3TriIYyPKSn0MXPUHNym
CvRJO2mfiAcWu2+zT/MTxxT6deQPdjkh9mkdzlR07kl/ywVseQ5bgeaazQqI/jis4ZG6kkTdUWM0
o0gHcNVoHVtgAGzgSM7DzIwV6jJ5KkXDuSsl24d4YJldXFv82rzlcGQBuRIqozki2UxcqsNHvhHf
doBgfsxeVRUBXdBsb5jl7wvpqUPypWw4lHNCE51qxI2acXBzPZYCi79hE1kvSaO2y5A9TwUriMuJ
feUlULHk/zI8UxIh1EvIpQwklCQE7JP7ZFJNN1P2Z+seAJRvQSXDFRite6t63p/mUItv14eiwo1N
Q95f/BewPJFRmR6k1dlI0otz6KvLSNxgAyEs+vQhjwWHTTnMag2gAZc8czpH/wRvyBlvgDIzSFql
27dpeQLHxzJimHbA79/eg7va0h/7WhG+An3Cax9P/koUKLjoN+I1/lMKXvYDValBLqTN5rMhTQe/
8QACJ8akmMiLrRayYy6/UeqgxihVSbnjWiNguF4hp4UUtZB/+Ku9ekHVvSzuRoUsoF2P26kl9ff9
xHIzYLrpv/IMdQveGAbQ8HBvAW2eaTmzTVRUcxrmfwAqECkyC4of2PNXqlyX09aSy4PY1r0StlPR
Ez11L7riKl7sfd3AVZLCySavxeJzJyffI+RXh9+S2rJWIgEUMuqr+paz69AU5/qlfRUr5iY+L6rs
Q1r5TM4jc1OasPYK2Y2/nUH2HmGh2NbkEpWJuefN8HEvwNzCuvU1d2xE5ppBeKzowqLxZhqQSbtY
DRDLL9nzeH6CP/RL+QteWtjj8meav8+uGbXmvfKkLwWz0GXFruImEa7cLF1/m2lHG36u968bI1mL
0bu1N7ZsR2jU2lQUa7ccxPd8FZ4ia6fJFVphtwRJ1Vlb7uQXCct/5h063edVvZRJmp3GJfFPmLgg
aUeRiLpv0l9X2NliiNxtCOvQrOxy97pQ7uBG60mpHEOHLDSt/KsCFdayH4MVUBS+/9UUxVBi5/xW
QDeVYUvKYbu86UCfbsqbmr4lAmh+Am57Bsxpg26+/u32ia5amI+iqa+mafyT8LQygd0oVIsCAWnH
MFVeaknpaS0J2Y5KKMKADg7ox9lM23zFgIRx9wT2r5zxVDD2Z/3bqQPE26P8n+5v/vvIRKMYSiVB
FlIhZBN4oNdPsrQYkva/9XRFa8ppqqovGs+tD/Tqa9TdiVU90T3nC5PZGItbyjxuWOyeVAWVFORx
pAJMOSPvinD30PwANZKwivi6YAEaWJ6KjbRgP3EtkaXOhXdlNC6mnJxcD2JB95ne3ipCWnTHh6mb
2eDlxVu3/FdDG3FbcTBkQ563jpcnDg3frlq0R7dUxLnztBlt/ZicBHYm9WHWfvdLsz5qtj3X60nl
z7OKnBvDWMHQyZ0JCt/1yTCmKPCbZQNMLGyAvNboIOTX6xvVQ4ppsAAqIlXgHmVOmQeuscmU9VWt
Q1i5n3hdsqSkMOBzBYgCQOfKLGjm6oxdyZySvTDDmHaNLOTOZnV2TLAYo8HGyS5HdoTa9WAeWFUe
9jXk7zSwfZENpZI4b4NVCMg/1ZCMKGULU1Lmzcoslj8OBFhYvTlvBYN2UdhpzdK0R2aMiuDn5Pul
YjGc206o8rpVvZ3NUr5sPPVTt/BStIdqyMoiO0PzvV/3DmfGI/w9gnYhhoLUjNdXZPQi7SaXc6ao
q4IP5l4F5FUczU4UF5wMLgDmhfGFcGcLrzn9YnOsRoWndbIbGuee9j/+qC9jadAmGz2fMkY67NrU
IEgLfhLd0S/BZ5hZ8FNqVgvDHssId3mgP8Lp8Vc0CC4N26vAARA33ilJ/yeK1kvSvL0cU1vmTib0
l46TwLU2WK3OCfevm1LOVkQTakxAQM1pf8AEcllFZvQ0/x4qz+hhrtgaPKaMIn1mk4vHCALJisDx
ZLgdNHf8dhGWM8js+DN8IUPkuNLCrMLSbDq7lP4dJVZ3G2vwyscIRFXvPMjMRm6qRsVKpfcB99wk
wK7mWJ6TDJKOhLZHv+haLFLU+UlJ97GdLLjPKXzC3cy7dpxJ9VS9XqpLPXDISnVjLlN18RjvlyVn
eMqkmbS9t5Bh4/ls3Fxm8F9r5S7IsrsepE0IopowXTbpAkM0BfNXM8IoPxMhJcMJKazvcqpVL5QE
s9rhcGIjOQSqhEsY/PMPaokq/M+Cz7KeBGyve8DDjdRsFk4QEuNFNZdmyPUEgCVpF7z6BCxyDydq
W1MvnD5Fh8czZG0DqrpGMb/I+fN7zZ3OL7BZArRZxR59SxK6xuOlKQ8XXrYPJqZQc5k7oOF/6P8l
lnbnO/zsXUOXyBGHVdJjemSdVVBqLprsYuAW2lvs68UfpDK4rbwf4NreCf+Hnzq0H2I57txvJbgb
wySuMbLoN9nQHSyLx8ustl3XhxE3nUBJdtb9Y67ZrzQmvF0nKGLRYKLdM0C5Pu4JCStpaF9JQihV
SMtUtKNOtW2SHnsbC9wp5h03qA3N9z3sCrkTPRAol4Sy39oq4ScRLvKY3hZJVZwd4KB17e4Yd8Xd
tX6jcr7fOON8gpb9k3TEY0rlWBbhsakmy42zH/xREY8jTvK/TlB3QiOYzp7bZ2QepFcEzAtOUkqI
nCiJpGh6WF4QM1jnT24gYkKQnu7TKjUtvhlFbuDGGshICtIl2PkMBD/wSMrcrK+I/HN3kRWUz8iI
xi2417rLgdqhmVcCvvznI9QNDAEA+ZFLnAktfBZr5gok+Bph3X2x8kNC7/v+tGc839aXyKGX4EP1
79yUqnS6C2yZT0poxol/cjJlT29Isi8Wr7WmdZ2TPPtTDZtIpmbAyJnFcGDaGmxJeMN1bf9aZUja
BwsL5kWMtjmEMXREUtQwbnwaSMTkNRsm2Y9LOxRMnGwqwFK4daONeTlMezc0/g7L7j8EVq6UBpEY
3GEDdhqxbHrhTLtxlXkVzy2QP9kczQtIP6M5qY3FMtJEwlonLBl7BU8i8c5GYI1ln5AyXsbLdeYx
xIrC07ywlH5fBuR4D4tfAy+TNHaTNVf76gDLEAM4lUCvuZxsDCNrhPZmJ5JywCqSxG8QIXFJEeLm
HUQ9Jh46VV/956ym3klrQtRzQ/LXSz3Lk4MpjRNylc0hfUNel5A5wf7WNTlQC3lE2tCzkptf0tfA
tJA1YWtQD1X4YuRw9YOxOVbPEztmWVV64afTYJkeqc3TWuL02ulQXwrBKqSVQXWmcWht3uCIoC2C
WoGD14vBV4HlVjx5diHsDmlNfuz8V1aGjwa0UnJdJoXFAycTdPpUHqpcNb7fUqvuTW517VCr2Kr9
7fvo9upTSYW3yBoE9KAT+Li41dc18fSzWdnbR6Z62PQKO0K3QSR65bY5IxAwHHCxY73bsrqJ9VlA
LQNQSWrEvlE/zq/x5uM15tuAHQuMJIZwaIucv0Hma3Nv8eKfI1mHV7pS/paOPN+JBaR6cDo/rPIl
Sbfex7mvZ+c2a2ZZlwLkMXrY4sFjleu+no4ALODbfJ5H9czvZhOpMGaOimwg5s8BJJiG8IpsEuN6
UQ/+tpfFWsXW8xsbUCJVviz3fLYSH/r3AsyWVYcqn17Z3dFaw9rGkvVRLfCGMRQ30alRfpkpLVLf
XOltfCiy+AEs9n3wRDeyxilVWB0X3hQZQxMzTnyu4sCEPcOTEeZXU4kFJoWfiT66GzNTUOgxiAf+
99uViRlG+QkeIXlAflLvNhrtHSUcPrG4sY0E00SqtJWAQJ9sM/qFa0NfOJcdgHWd6U3XbuxKOlPA
sZOjmFLC6EFc7uw3J4YBTRPn6lTGAoNFNAgDo+o1Rd4+sYMps2q/X9k0tChtHmUX2Q8o2xtIwfY7
Zbt5LMNmK49iRu0ebbo7s1w/2oXPC3r5+Ckp4NbZ01w4qCXvX2KErNcLspFk5TiBGLfst71dGR/l
4AedkNKWf+p7zOlz3y/7dIypXbkKig86gmjYIK1xTZBt+MShPsCopcgDEJ5QEnAeLKMoo0aN78pE
xRZhO1VJ3sEe4SwLLY3Bce6iyaE8dSxCf6yyFpLU4hnVgY9AUrKJGSwj8pgxzI9JCCkeAPgJkn1A
xta6H4q8Rlf4QGejh+4IgEsBMO9ol3AOmkbgUgXQjnjLJqPQmVQd3r06iSwE+fgyRed8Z72gZ8FE
O7gpy+FRs0RVoglc+aXxv/QHbVSkf5Tmzb1zi0VmWVXyLXYpg9ZBSOChPS46oD4ADOHxJBrO+EhE
qnmC+ohw4lRIC3ccLvQI8MNVQtxkjjx7yyAqevlhTOEhHVnZEmno7v++jdXnZSCFJy6HHxLA49YY
qgasyA1K78tMsXPXRyNVdaXyYrkpeCg2O1Q0eUPQE3RrxNmFeMBfKO5fJtghd3wwB/cetjHB8GfG
q18ORefmhfXvKxFBEPwFInhdm7SeCI/6uafDQ9fKl+N0kq6ibkq5pjyPuZbZ+xsKl62fWYGg3h89
Rb1e2jy7rso8UlhetHL93Iftj3siw/+0grIRhOoPNZlP8/IHgPXOZ37mRXte9SvlTXbYPAkXHfEY
fRr85PVZftmbUfvFD6rNZcEkGCSfj/E/Mm2M5MVkTr3yMRdSYi/pBUq6WJbC7M2eB+BoQ4qzzW+n
FvN62VPX6vxGuFKoepuaGuToNHrwk9+gmbQx1BCMUyD6AJ7GjZpQ9TC4Lde+4hGHgPKZUZXGHXCv
lR4duOS7efcMdBbCAUq8hWny4OGahd2pE65ovgtnOsjhfY+90/m2bCffswcbVDoJcDBDaXndO7Ov
Q0uNm8RkCBczFCnXqU/A9UEAkUf3fyfveR5Vb2xEtcxcDpI1nke/p7uUtRBRBW21T75URl1lAXqG
65MLKPTHGCNsTdWI8/g+Upmh76IcVxsJKtb+nI4Tav8DiZ1+LAkpBe8025j1JGXglkA3vPoKmuFc
4hjfDfgGS9O2aY6RJ0+tnA35XLgLjA1bb65rY2bsWxEzluBfV8b6Xl1lRNFRTAsQeJy167DO9rvK
p4+++XxxBYTvtGHjW5c/U31YXGQX0SCpfMt0LF9egJhO/R293hjeVlC6f3yhw05H832t4tzcTYAd
a+jHCT8x5Mjub8aJzt5/cioKea+a39snRwO3IPbFzGnSLH81iwxQ61mqiHbxu3x4Kw3BBc13ZZz2
DL1YBbwL6GT8nz6eDMGlL445sSLIP9/D9PhdMkGsmLIEHYHBI5TfPQppiz7xBYiSDPI73k+Mu1Gg
KFt4kGwvaxW3lgV3DK4MQ/SN9r+G9O3XURakIPS1sdDhIFn/Hv7gl6J7k36JX+8sueTr/gG1r29H
SvH6ogt5TSNHUrn4YN62GTjKbPvbMIzVY0u+HvPxcK90bpFIDbiv/DBs6oo8M9RWCAX91uoQQitt
nQruq2+zELHk5R0/NXRZOe0jNMMgTIuUBi3u9+RgWv6XgM32RvhvJ21qPVysFuMRlCZCmF713K8a
XsAvFO4CHcugouuG6GjV2i5Qv4ooV2rWt7JuS7JHemer6ntntmTAujBxxeeAKIIRjamgNzPoWVCM
Y1vsFpjMoKlOG+PDr+Eq1h8+PWJbw85VNe15Sjc+dm/CjqknNuTKLRv4ltbsexlOI3TLI9XeGdDk
FaL7JZ8LcgJCmQZpQ9r8qmtrYD51kibsouXsEK5Z3aQHL9gr2adZERD6Kkf1vXXax0epB3maky7v
TFqnzOgJHfFyVujPerQVVH0wxlGMDjPwxlrFnRXEM0P5aE7dn2V7GFDLfG9Z3zc4z4Ub+oVV9M2P
6h0BxRtV7scnczaUrY5hoY86sBpavZGT3lSXl2VOM8RekG8j93vRczOIWY3YntcmMdrUvgIjBTUH
Es2If6MM7nxpkoDIJut1FDnhbYpxabgkNvURywuHi0MkdUhvpgWsnDFyTFmM6TzIcOSzhEBNeVSz
99EHpw==
`pragma protect end_protected
