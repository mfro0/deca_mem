// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.2
// ALTERA_TIMESTAMP:Thu Jul 20 10:40:50 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C6K1vnnPezFnG673EDUDWW1Daq4QtfxleqdlDjSohIkOUuMv9hiTcfRbM488AO1s
JrwK/IRT01UGN3TvKX0wyJN0H+RztpWA9u9lXZycQSuPv85GpM5p6/eFY0ClwfY9
pFnHkAXcJ43xtvcGXSEsWhQ3EEtz1jxNhufynx44AIQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6016)
11FeBfYXVYWtVkCh+TR3wPUMX6DYJHeced3jse6CbCtE0nnCJ9FNsCrEn8uUHERD
awfZO9g3HOecPlPyI2ne1nP6tPwcijzJFSqfd4cxTuJbXFwbpVH2+lp7ViMS9h2E
LqWxlKEHbq42q6kpTtStYgHnpcDlqqTdu8pIHrqTM/m8gJwWzYawKfFgxHBPHwMB
Kp38ZaMAmvEeArrFIkIqbPGGRR0wbXkEoIsFG0zkH4ueup8GSEf92YaVfBQBlO/w
36CIry/N/5eWmtvCIdln/MAPAyFs5mAfClkXPNCUuognOdIQpC3NA5kCz6hW5QER
WYWksUW6Vs1dP678/M8qAa/SQSSvdJJASn47/CsjVOwCMoQw2eni+BFARl1svdBR
ACP7QDLllIAjXiOndC5gMx317+J6MvdMeBWQ/T72LSQAwpH1tYuqDJG1UQEJ3sAk
9J/wp8WrZJpup7kqFzOIN45aReErN74MZQ2NYpWceV828OwO+t3FXSceS1wVCgsi
n8U+6lZ50Nk/tI8KfIjx1OpOKlASH2Odg7AqbF5PPXjG39g8xOoRrB9lFm6hE+hg
fHsqac43GD3ETyl1O2r/oSggjS4wrnhX1pVcektwJpwWKRAqs052uQoWtkHyyLLn
EqdBi6sob1ymi3QbEpmKlTHdCBYKFtZbmurNA44DnebOK0s2qoSKLf+HCz7QMsPc
Xwhl+WRTPAr6v/AaTVnmO4P0D5+ZPAeumLEhL+T5h5n7INnansjk+k8Yqh5y8RJn
/IMvT1Tu9P/amzL9qBWlxT6czUlk2V0s/Tk3hgQ+hLFb/QeNBTkBojkfNzx8hNqz
3Clvj9VKwuGMDhtvhfdn7X0fSEtEq/2k3z9MJU8scLpVJ5Ve714ZwUBY8Q29FChY
9w8E2Uc0c83u4/aAOS0CvQgk4EgmEtOnLW2+k2hLIdMcoZmCtLuJ/fMI5xFlLYEY
alddS9QyXA/pv2buiOB4Hc3YA1frz8x9CF/KkJ6ziLDGOvUh88kMrRpQRSl5EDP2
MTt2kTjCslZSUo/3WvnbaJ1y/wT2p+47GJ3vbJmICm12OkMoKa6Ai5rDLG1AQ7Oj
8xwgdG/r2AowsZp08dPvc4xuube6rNLQiiZNe1p44VGbXalXvCZtAK/9uRsYqvg3
7hHI7c5b7NnzORkVywglUFQdGoolT4jrEUSxqbsfpAkuxe4eLCI6PxfAJ7EVhu8Z
0KFtVLWym5ngfJD24bR25fvq2JM/U11l6S33Sakm9BRwJ6GgWessm/Qe87eopU16
X2Iig0tM7qgh3c3BNKDBkPt2zynllttIcL/5kWyPgY/N2s/REVV/+DpvWUlnHJVK
g1M1PEY/6cqyrzsqkRluFYecKDTRssnIhDxMNclaTjCU6cCQCADhnvAgDZGFZFQh
N1EIkcDgvWMrGAa6wLTDEB1U1txhRp/dlW3tJQKDHBCdDE9UM+yBpz+h7TjSEhT6
mZ+RLffOiEjtoe6t2KNT4nsol1QRbzt9+SiID/YZ2ImQdrrqbpb2hEQYgpHClcGV
xucz1p8VFBhP45Ccy/4K70bx0TvOZNlRbcVsdjTdsI16/eJQHSR98zt4pgH9NYST
XBFh77Qeb8corinjypRcJjBHXWSDJVHO5kumnHq+S+Hxp9STqPVAwF2TpED2oLWH
72uuHydJWbasHoMxevnJ63kJmXhe7A9f+xCJyDdxQ13NFBjx6YEuCNVLPXHI2dkH
+5vv/44ilZvTzwz0PagC6zD8pl14g6gmFn4idHO2A6UsXgDcWvAFZfiSG5pT5CF2
Gp+ehlv2twbgamr4IHWrH8L47v2o1Kg7LBn3h426qW8AdmCTT0e4foKbCFb1tJE7
84lYNFu3Tstu1avz2Hv0Vwlwrcw+hbTSDJSkX3jNQB5p0HO7wOIQsza5D4yMZ3TP
84FwLdbMGBZ9j/SKTd8ed83fwvRyua+nl4ZEV2/YX57F1FNBTfDn4h1tTbyoXpt8
8nDaHFwVo3wOO0LdbBpayHXskI+pT9YdC8jLp5YN8p2kagkGSANJDP/L5p9odMEM
rKJCFyiVu9E9xd1/cxvK5UMUNt8XHQkocdbHS7FkXoZ/8n2swLBb/stxmBYnH08x
rL1pmmyRBqlJ7+zC1gwcgWcniY1nHdhEsuicYmyM64K1EGxnW6VPsJR7LVErWFzz
YlV4xGwUqwB0I94K/Bvm+4fyZi2dSO3sSCkT/G5mEvpIXGxDOMmGrx3teXM9B5wV
cBqWBRfE1QDelqFnq9xSGcoUXPerY799DyAZs5h2ne/wtBQakNvWGl5i3aIbsgmH
wXJ8/fbE5WxfM1KwsbXRVSrpGEJaIYBymVZeW4Lc5tmT45wJaQ/1mI94D/3SHoS3
8Dmu8pzm4ywg2v8BlXJ9zzrdaumxsuyu+0c+28xI5IBmYBByUAugprNCL6oMUvTh
PL1gMThaoAP8NbLkd8Sne524M3lJDhgbHUQgNa4c9GxfJPeLvc3mClO7r6zi3Oyq
Wu5gESdAEvUOVPDTbGauPAiNJHKqU/18ETjGFjbRc+ieX4ePvOs3VGLySI5qHG9Q
3h27/TC4hKLt9b707UcmZBd2qcWLebus46F4uz1GfHKU4HF0nJvDsZB2bsR0ZpXZ
6xwtrms/Q9s8QOmY3BI4jKaWeU7yf9hcHhza/gPba4inhEZcSe22ZxH581dZJ0Sy
7La9mEzK2E8Cg94ncyNc8gTeVlbdr1Mst8eQi8wERcz+ViRSFHm1HGNh9avrEpzI
0OR2kw4kLPXD6tgWZbnIsYyodt1pPVhHQEZYEO1bHmLUOivDtB1DWXXkhCCnVCJg
aZ/yYzViyK5MWFVxA8qwWFJq/PPOwWXW6XdPL3fo+q8iGsQ1ERHyUePEmo94OrzL
D/XbrxNY679efmAAfh57JSVWcmWPIAFwlL3vnJZRBazk9fyRb4w0YtdzwrqF+W7y
D3/SgWJFdXnuPi2vvEx6IHnnpmNLCuqixy5frkQXHYRLOrR7ddV0VB9k6bFTWPzm
oSp2UIhop/InHmIDEjTDyaOA9+KFlm3lqPpjbstF3ZiSD/kUB/WFpX+P5WiOO3AT
WJ1URpvK0AHj2MX6UWU1qs7E88VAOTl5Pl2RjgMZzveGdlG3bHCHYMk9KqIA49+Y
9ua+tl7711ZI7Xyu4migA53rj9yscCeLrMOkA4oKxfPndi1xBavQ5ihzgUAwCZe2
7C/4VMI6D8ByG++NsBv5HluLym1H1NWr6RCve+3XzN1oTv9Mu/30uM3uFvn9Fcbw
QLPnV0fa5NnnTKyzaFfi78ZcRdd/e1d6JHClIsZzWCx02YFjPOc8mkyVfR+2Gaq8
qPm7EVFgXM19gpkCZj2oreADVdQiE/bcobWcSctLBn523rNxvmj63I86C3FIZ2qc
SX5K6See0aJvIvfDIzt9Gz7Vx6HikjGojiwoOYPtC/6dlMUoY2qO4nhSt7EsSe4e
ISEX7COEMyKn3hrkr0PsxtK4s4OAPyJ3yeTFxlpikwusBACgG+IJfIejj+msMVC2
/QTOtzDcKpfiM+TDMKjqZK/R0ROlsVCyqHT2jSEUXIfFbzPHZ/7sqCHDMYIfLdfb
INTrce11ZTLMfPFr2H9Xf1q+vVaxd8CVmkWOka3zs2hM6i0dxUbKh6dqN/HFqcu8
bmnO7NS0Tt7ye4Agw/RajJMFULoHF+BqAM9drGTehJ/kv8ywVMQpvf7ndlq2+yd7
XXyckhaa2AWVbtBHu744ptvKJvxHj0KeD6hzJ7ZU2jWxZ6jYEOlVR6UuX+A81ZLa
3/BvA9UNWgobdf64uMsIAImy0ef6E9h1FDY+4Z3c5I919h4rcdzP2ASxQcIeV7n1
M+CZRjAqywntjQCbTw3wy6G46/oGcurRX9YZ1i8oNHN0XBOASUeZo6VqG9aOXu18
8zRvSIy8LAwmwaA4rYUl7OW5ABbE54jNg3lOySQXGtj0Q9MsO75PwdI+psAMaaoV
g+A/NGSZI53ZHS5uSL9QMCGlLOHKcq9r4K1LySm80Z4BRhPf5jYIrJLZN5LT38Cc
zOEiqJz6jeHY996rfauPkcbO9tujsHk5y1DdVpSfL11cc8IuxeWpdEAnolfm/IWh
tO3kz85gDUpjEPLCp5XdBMfFCmo1ZgPq9nNur4NkRgnFxt8yMxMIUtXVyDazBm37
SL3mFabIBC9++fnxDvono2RRGl8N/dpm0B48HO5mQDI3Yy9KKghV8DeNmK2FA7la
74NrCJ5hzOWBH2KHmchL+C0J0ZMgf9HXIzAlVH3FqRzh/4tTs9y3WQ2z8LFejI8s
W0vmK9OczrwF6jI4bvclcGNe0gf7YRDId+LrrXdI1jYjXEcOiKtHhHqG1hwMKIrQ
xpy8xe2LFSxFQsMRw28eiK/Wt8Qdwao1lZnmGF7PF7qL/qfIWUAkG0vvZrUpYwuD
J0PxEm7IX0UY7eEW/FDp6sJUlPv+RafZdhmJCpyQsbVHDNqY2b5JtFvsdpYD2+kz
sb+bSgmE6J99+mJf+Ywd6zK4lFuP2daYkufwdrN85JtXRQEu3+S5PjdaFR40s4KE
NU+k4hnyRHSkouDmF9YHxS7KDTtfnnsVFD0T0QyYSpIaX77fKaj3sH8LDqPcE605
75SchwAqDug57CywzplTiT6COwOG2n4Mj7S1YZ0FIgHOXMjqFtcEN6nzceYCh3Ny
rlS0qgCdOUfaajzjCHQvTz0SACdzcgm24dhaAFq4AAmB35bU7aiQ/Nyg0I11rBhf
4m/MgyyYxLE5LKJ7yhNm6Rcat8Tz3D3LJ/W3C5ZTxlzqOUATc8WPXGKXVVtvmuAb
0/74PoyYR1oLJm2fOzl7VfAHn2Dx8RQCa8PE2HNvs9HiZvTzznID2Thk8bsiIHuc
tIWAZHvJdMZj/7wX7q7sEzoqfpEhdZJjek0S/XdYiWBFO3F52r/HGYGRYJL+DrFI
D7dKePz7O+/+uejx8FkrvYUPphn32i4kpwAdjDxbHj69Kpwh2U03YYxkefgaoOrC
8joNcqZdvY0U/PN2Qh/J/iVaRab6xwjjZm5VvwcuENXpijeImZGaP9TNZISojhqA
N/lp8tMVoYqQTkvjiUkKmkQN7xWJ0jEuiid9wbHYMP7acD3riXC8GO/lPEIXSccb
uYI6XSRQHdk7JYLfGSpuwpDuaMMAqHo7oq4pcEbxgnDXOMzpbf9qpwF/dRIqN/HY
x5TYidhH9Q6lFVUTXN+jsbRg8iGj+sUq2GC76BtNCstjIqbcSqvQGE4Rr21LXy0P
QIwW/dt5H+Q41Z3My3Gc0BewKK2VgDRp9QQSB3caPa0dL/d0JeaSS6xacsKYtYOo
5E580qsUY/YkTBgMu5NBE4j7uGLOdUSTMgmn2pbZnU5rGyarornDGIr/ge8f00bY
GNGgMFvw3ky4pnP8YlyeugSHAunjtWmFtth0lwIYD5MAg9Pzv8nwADMrGUEZFPPW
fXpqWld8jZM77Q8dqGvwAM48juc9aTLSeT4XbFV+knCFmm3qtta9CuXNU/TeCv1Y
1jlZ4wc2s0RVbl2lcjtBiFtSvImyG8cSP2Aery4ChjUvsazhkPIb9NDvT6IosR4x
9tZOpKb2oe17zsV4qGs8KbRhaIobHuSZgPQ1qaBm/k4NWYDdx9brjK0HYRKZNMdj
ZKr9d48n+deeSCsl+TYT5a6aBrC7RqEFWy2kUNxEQOxLizKIEDKHEdNnbTjSpJWb
EzP0tGzcex9LrGjCUafPVV1cokOJn1Ik1sPUq1RdB6IkNTBWaEKt2XPIc7VeLzB8
emGDvFdXd3afjbsJWYmg7JzZaDaS1vSd83G4NxhCDgAkyDJT9wo7G23y3MXqa+13
8zcrKelrBXRgsYMzgioHlmWSfU1tLIgmIewCU19fWJxTkcrjSMlK1zZHOR/uYPIW
/QNtfYYfPbwpB+rqhjAUCMXdlSUp0QQgUFG7Ko6+EUbjZkW10Wa6Q641IwXyZFNO
u1bYCc2rB0siGogSVcACeH21dzd+q0r/wRHf54i4K79Siak2TuVCxh6NaKxBxEZl
jAoBtFy/7/wdfbFuKVJGpLbDqGuDUeQT45NTMcMdqBpGq7eww/qqDApUCrYXZoJK
jlW9cmdBTO+wBrSim6chayyfzHY4CzjRbBgP18XLu2wEfCL787cvKh6YteQMBuNv
sB1YyjHfx6Sx5GapEqZLhgfto+YKkBBjZHp2CZ+qwDvQtx6fvL6QSNgwb3IZ2xym
KHuzUFZMOdnKLuyX73UiXM3YVLiMmfo3Vfr8vxqtSNDElMlw8vvoANhwhhhxPbZe
LRVNQ2NXjzehEIah5zNfCag2rtCDPsPvihf8H5OJOO+1C1rTP8hXUKLIVJD90d/E
ff6L8z84db/H/lRsPmKldAi9NV7PGBD53IZdzw6lg1F+19wASzmKqEW8SDJw7Y5U
7WmOUBWY/eauSZKgE4hqzjNsoCDObedUslXZNlyv9q2OT3pfRG+vMzSgB28OtfND
EqYbTcv75764sSScqohdumj6RGxnCrlpkTDF3icJnVL7ed9sd9fgDyKHm1seraz3
aL6BO0s8IR9aAJ/jwo67XxLnv/566bqS4NVZZoy+zKx8OFv+e2z59I30Wc0/URoL
iqygdLRJbqUvHA8kz58YDs5DNLGuIPx6Je5PY0zSsFh4ffgI1Ld04kp+ptiYOay5
8eOYoi1IJnSBkP5Qy3kIZeCjamx5oyf4h9lKQ0+6S4UBDStU7+0USMsylFT+6eHx
81soZvzmK8g6OE4DevsNGjdMZWSzgd9QwZMWiZMGAmNvd0y34gALyD+XJd6rbiis
WQnv8DwBUm5r2OwQm38Hb6VycN9gLTH9PUL6UXRglhiWKfjqjSuhhbyyfSLmR4ui
OF0tX9l/xsoViH02qS/0LCQMilaFo/LdsaUaGTlhuItvCmJUGHHHXAlONcBUXoxo
UQgZ8mCBU8R5lFLpmB0OGPDQ6VADsOE00KGPIE8A0yJmyIJarQU6PXfVx8rQJYGR
AYmn1NIVWMFch6t7Q5odAum9sk0YOIWIn4nCMyy8XPvyXwtNT6NOFYvrvMXAGLaP
NUwiYzpKAfH4VkfHAlYkO+S2dgDUh+bFAjtHQnVNLgRy657qn4IerrmtGesqZ2Ry
NgzkMwTXOwfNfBDke+kq22Lc+7FPtOSQ0rYk6TpGXWQYaH+T364OFbWAiVEKqLQA
ntJX6W5c8Kc0i94ECc91mQGWEqPAi9BpsX88iajTJDREXFI2iyBVOhdgs/BdXyMl
m56qhKQhZ3sysMLYao6Rc4lXjV9hIJEdQYxTkZbPp7/A/CQeY3YaXgtk30MAPST6
gadnn17xT0b5IzzOfuqMtChcvsn79JrS5p6Vh5LhL6KG9LE4QMNidAgk+qMcixMN
cpEFy2xw2XnqIUcBbcm1D5bA/4iZnurd9LvTjNTrjBdJdAdF+wAxthasXJXLL21S
mDeriEB52bmd3CqaDub/f4AkiXtqAIOdmnzahNg9Pe9oLhMyqMBh1YBjfV/oXbtm
d6cPsC5L9dXw3Tl4n+0A1FYZh/K5EGIkASs+SPyFuVKY4LyJgnDf3rNHsg3k8SV5
t1v5lgbMXXEFJ0/yTNoihAWh2F3HHVBfan/cg3H9q+4J032E4QH4WIhic71Z7cuQ
LGKWCjhDMY+Ob18VZByhfeIT2D69dsoOzGIW8lFCCOTplDtSN1i+QYXc3cSHmtBr
3aQRug5T4/S0m5sLz84gl4smbYJwhvLCMUJ6m18hw8TwE3ClbZx57aq998Uqy0il
pcfsQYfhdCQnjzshGYiCN7VlU0xa+n1fGRaUlD/OG13V5+M9jqqaNetYi1LqR1n4
5qGOysnPYMYpuortg/iAILyE5YF4EdmGudQcyaXwbn6EiAgprljF7Co7gQP46KuT
px4POSXruZVA6cJKz7fODuX3Uew8YPfQ+9NUz9kOYj7lAaUIDsGji8GPJ4fE4kaS
FYeItsb/Ylmpm+/Igbt7xwmOs75uprfPleA2i/lfrSde9i5JT4YFNbjjFkg//fmj
tHueiyukywP6/h6OWQKSYA==
`pragma protect end_protected
