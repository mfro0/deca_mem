// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HH EA7C,U62EF9_HC&V74\R:AP*7:K1!<GC\RGQ22B #472C:&Y&=]   
H-J4/;**S0>X>=MQ8 ]$V8@):]KYB*:;,+$27E9&M:E*2%&#G8N9!1   
H#JVTEBO)/[ 4RA!-(1@3C*$_.KNM1R<-5/3Q9TM^+QK0.\'"_@JFD@  
H?A#*RZ^("L[!:8H%2KI>\03C(8KGA9D[C,()/WZ52&#AJ^:&_!L=7P  
H=6L>W2-P/[A6O3E(S6Z.DH%(I(:#([KVRTML0L2V^QB[PD2J,!>^A@  
`pragma protect encoding=(enctype="uuencode",bytes=6720        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@8JLCX?DV.?"(P8?%@^\<23MXAJ&N!JB97\I:#^\Q<BD 
@KV\44U,F'D(>H:4G0BZ<BIV>O;8-R)8,(UN8CM/POM0 
@T/V06Z* *N.@J"@0!8?1B8+;R^3P(V* B\,PZM0,>P\ 
@UM2&Z%"1PTN='@%OSFR6JA#@U^HVUDL..XDQV26>+7\ 
@K*0;>'D)&*D,/$(B0%@;?D5PTFOV"6?<,3VYV(Z,-98 
@(U%Y<U5 J"Q-D5'B4]EY O:6XE"#ZT=[T$%C< Y>M"8 
@GX9M622B%8(]C-_)\'@/[]&@O%KT7-2Y90>VC@Z<!L, 
@;H![ ?'S-YP"S,,]CF!SA+]<LU'-"E75_1Z;7$>63"D 
@$S8C:DF?^)YG>>=2UALJ!.7<J]*^W$G#C@D(VDE=$G8 
@1;%78<$\W\I"SXP@8]>[I*0%<G/8-I8)-&2-$ 2WKA@ 
@#WAA,4%7KN,ZNR2!?&2DX=)*@ RS#K3%J&2>\NA3)YH 
@WS.WG9KC.) AN7"&NNNF;,Q&\&ESAP-NZ%<?A"A[Y6( 
@^^T/AAU8KZ;%O8.$>J+WP2F SXH!B)P>#\^7X378([X 
@>J7ZW.3H//M,H['H\'2L1)5C)F(0"2W-)T*$7M=Q(A\ 
@)N,&I8<H%WO%F6DTM+']:Z%!UJGZM4%L\G#K<+;,&VH 
@#T@:3SDM$7E]P;9(\Q'EDL,:?7)1G\135X:P@4MG,&P 
@%JA]%% S-,+O*4.)8#X0 \U^(T_*:3A4\\<I A='@R\ 
@( -:\YJEE[J]6$1*5!6X9O,9( ;Y:F>-W=]%M=> =W8 
@VGY$B9D%[("1&^1WCU2]QH4;[@K%O  EE:N425WOCF0 
@%79C:P-HR,Z*M.66HQ]0RFQD_%_7#=0D_<;CU;?*L+X 
@HRD9(>T:^(KA%BL)1/=/X '"VF-^Q"+*\U?<5\ !.)\ 
@XCRV:G(]5FV20D+70T;["TDL6I(SWF+4;,KD]P&JJ/H 
@N+/!%U#S:92QM?_D8QGLAN10Y&]XHY0I,&UL:.W0HY@ 
@K&H_!>/G^N=_UQR<CNK_]_?MG3I5C_<VC9S>K'$_CR< 
@T%3!6?'^W3 0^JM+MQ@+LMY$AMZZ)9$VM;P[!W$N)7P 
@:,$X#G8Q,J0M(TR(LQ+>%F/;@-/X > F<#'?\&0.B%8 
@LV^$POF?GTV47=U,CR@9 O>+S9?GS6"5SPY\/!8!"0@ 
@0%!,XI9NIG$KB7O"OD1Z^LT3D^YG);8J5+/&_,ZEC)L 
@6)RF1?RPKB6>J!=]Q5AUKS7VERQNH-=!*:P ^!MC*O0 
@M(T)KZJL'&)?UYWE8ZB:Q:,(YM%1!8F0928!J0IK-T( 
@10NQ&\RX6M';<;C*QA'6SO9PDHAH'QJ_1_^W<18:+)< 
@ F\5!2.2HI-KQ1Y5.<N#K4</II2-CU7,"W$3>LE-M', 
@P?XSDH7XEJGL.BYU=5TZ'4@0DV/-IE*;;2+3@G4!:D  
@B8>>#V]0"FT8I;:T<GMF@20<#*T*+*_-+1?/<T5&0I  
@I29J]$Y+ _3MQ4Q5WX2<F1M@DOI9J6(%?1Q2R115!N8 
@2QQD3<D6-!!0WMD1O9 U$= XP12[A3^-$CZ-[AHS PH 
@1US-_\]U?(G!^OX0(<[0E>U<N,.,4/SGOL*<<1=N!-, 
@%:S\@":I4;1DVLFSH9._.<A3#>E,$3S-EU,4PKW'-8@ 
@S=$JZARM]@\XD9!O.!@!(S8#K9(E- 4;XG.>B#* @(0 
@>#0/[$EN$AM[0EAX'NP:OM$/C/G":*4QQDW9CGBB#!  
@+5FE43P'-ZW;S0,Y]Z/KX86JZ!<3+N08-T"TM7K;U+  
@TY4L8$IRI.$!35ZHN-:QHA3HKD7OIDY2RD>AL$XO0ZP 
@Z&=^PH,;"O87,->R/)IBV"*0<,WTMM%"Q:X@+%K/LO0 
@F)6$ZN%P=-D>40W]9Q6]L'P/L9?;PA+[.+WETWY\%6  
@34"[DFEE!7!3]YG@YO8[PYH#@-QA7G3-]:8RFSH]H]< 
@.?VO5V3-7.#-V>]110A$U09[=OP$?OV>=ACY.S#K N\ 
@-[D,^[YQVTNPX??.8L2>XI]6'VJC-4SW<-(SJHOJ-]T 
@@5\F)KTQ:R[^R.11)\"F"W?K%6YNR<=;G!6-;W;-I)T 
@T>B!QRJ^[U3+D\G'-U^E<PV%4O,I60A]:#)\=36%4VL 
@\L&639"_E=HFTE1 '):X04:2G\E\P)4K4/I#CU3MC.< 
@@2AGOS!E^1N<9%*VR]5K.#2+*4>3_44TN0L!BNSA U0 
@Y8&_R:W(IJKUX+2)$*K8F$[3J"UDX%$8Q/KK>/X,<:  
@%\&.&<U27;@R8IC&4QZ]N'-^"?-$0C5.-?<-OM6M<FT 
@N:BM0Y>RPW:XZ!P[9M9%&H>T+%S;N[N!J%PV._ZE7Z$ 
@_'$:J$D]  "23.3#DU+L)!URN,P56'XISY=7JN3B/"L 
@P.AU<1RH1:4>H__ZT1P^2<E*CG='-2 <K>>G6(@ ?U$ 
@>HI5'$LD5F4_26&WL9#38(V<)Y!+8H"KXX1QU2*7 Z< 
@)BR+)O3_N50<:!K%/HG' .XB#12_<GB2#7Q]+18W'4  
@H<4&4X:?<7&$_9G?AJ&('J&?0_.D4'9\F(4UO!:V-\4 
@S$ 44EL8\$M;GQQ%Q1RL:Y.CNGBP#.$>^!J3P@@'F]  
@?BAHIWRAH!4H;KB^<1;+E^%I:-A*0OUI50Z?;[0'['X 
@ *D*/IH"65.^O,M,GO3^O!4MK3D(]H3I9%Q@:"#+/L  
@N82IL^#ZTBT#_/+IIPKV?V]\D> &1_YJ>  +4U7^WE\ 
@.B_*(0!TYP7$98H%83X@O(=XUP+Q/M>7M_3@^FS*:XD 
@-#:-GQ[.%H;-+OR9T+:'@1AAF@\MQBSMU)Y59FA!H 4 
@=O6B7RRZ6:C$OVB&^'8P.P5-]\;U-^61)0..Z3BR#D0 
@CW6Z/T@RLA!ORYW.4R^4'@P<0AUI:]2P <MO=U)+VJ\ 
@*F+ K*+R0=,:9(ZV915O7,5D/8[Q/&5)#3(9P%=VCP< 
@.7G\&,JQ/N!A^W5T!60=I/JR%\%D/3:D\#KZ:=5LA1< 
@2I0!DV)&:V-]JQW*75$Y.R-=(:B'C&  26350#N?P5T 
@'\D7(C/%RUZJ!C*@[Q[4ZF,=RCU TK]5%$BR.'CJD_8 
@JWGT?5/[[J'YYZ6_&NX3X$+34T<D:-":[QX@?):)'&, 
@V((/^SVZ8<)>?H\W2F3"$16Y,HV= 8XSU4OA<$3HH0T 
@W!L\\F]"#Y26"H?>54\-:X8U<[IG9,Z<R!CNUKR*2#D 
@4W^Z?SQXXL^!+)B283<C)YX!-C%!U>[W9QW\D8:IZ[@ 
@VU2X#Z(FL-!1AM*5;J_$.6<_X04Q^O8=BQ,467U\QG< 
@VZI=:.]V=T9R9*HF24C'J@UA" ?PDEF-SK*'Y'I_6HD 
@!5")V$QO01P1)A+LE#C2$X95N"A_%O/^Q(RZ\]9[)ND 
@:H)$H(<#U-?\&EMYD?] &-6,\=J+P?&K'9P\0HEDQMX 
@Q/R.4*W3P.'@KX<LST=(:L2.:Q+BA_0W0 B3R>/N_4@ 
@@#!E[LDA4X.X;!=U@^87.,HN E'4C7%SUBWGULBN"*( 
@#:Z:\,F[(-[6?)&"!CA!&P'\*B&+S#LF%=-"+]VS?4L 
@A1K#Z8D'9*B4Q^JV^A&:"6.G_R*FT!'SO\^:T KPTR@ 
@JQU'86#K@H]FTG?ZZEJVDMK-L1[7V,'0R9#8ZYVK \P 
@V-*;[2KY6VSW=U#W0QL //#AK3V.OGZ%3X'8Q3Q5BG4 
@J2',*$ 9?"+^4;K,5%.I!W]8X\Z:0?D>\/*I^! A1+4 
@IW-T>[-UD%\1]H7FCJ1^,(O1,X"UD+RK62^-.6MRM7P 
@]?F%RF ^7C_8>Q61'1#HKTZ*P,@6AH/H%KL=0(\E>H  
@(7=C@_-A5Y?_;JYY&](KNJNY)5KA64%Z.'$3\,:FTQ< 
@F,TF@W-=H7#T(X)("'W)%I:82/8E:%JE. A_-5U=*SP 
@S?USYNSZ7$UHGJ7+X3"3,\>L&S1RP,')_FK+76Z1HA$ 
@6.E[S0;'8FI8!K9YK:YF#TL==7@-C4KL1ZD7_:-M.*0 
@6;]U8-&!E^<(T!;D>%,9J_RTJ:Y(V$TGYH.JIIUT::P 
@0\;OI%'B3%<B[D)W5@)>Z5M3G=)?>2SWHK5W*[T7 )< 
@#>/N[AS9:2;YWC<" ;5?QG?<4HFT+,+<0^!5(UI;2>D 
@9+/)?2-A;K<@?(UX<))'(3Z*>LZ_S>Q>NJ_Y^3#])EH 
@2SV:S77RPD+<KS^TR?S/&)-7D/%6;D%CS<:YA*>B^14 
@1?>W6K3>KN-G\C9UBB-)Z3(H"G*\GF7\3;1[RYGD#0D 
@<*V0 4%?9-JB)\HM0/M35@^,4O"0R>MP*;TR2DSM2IL 
@B-TO RA9)0@B7*%Z'H-H_49V2?97 W3F<-Y:CR=66O$ 
@FV$=5610H.:N!%WL;S)HH]4GE,3B9]_/QV&<L_U05E4 
@H[F1+_+=(O"RP3I@Q#;D&(>#HYP9#XZ:!$^8+ ?>-%L 
@7 V*KS9%+6J'B-01&40)(FO1VC/QLM"S,YK67(9]XX\ 
@6S"$,6.$:8US!DYRJ&_6J:\/X:D Q8Y=V\'",*DK'L< 
@K,/>13[/6E26<M/M*[H^4S?N]#]C[]'N7QA$O2#8X2, 
@B^PU@4?MY6G#U#8NH5:"]O';KD4T#CGPR'2R>IMI[^H 
@QYQ_OF*(4.;"ZVE7T%/]_1362?0IK)WF>IJA@*,V?ML 
@HNHKZ//.90DGEM[NG_S,6[NUNUL.W*PS? V>8L%0<_X 
@7-RWBO3O-L( >?-'DV=GJGO#Y',8N=W?/@R(VX_2NK  
@MC^%*M3G<1Z[?2[4HR@IM?4V()NWE0R^S3]=W*!3X9D 
@)JU;PON\*-;;/ZD92?G@Z=GBB_ZB-^^6>/N<2D54P%< 
@R,3\,\<38(8P9%CX5:%Y"HYRCH*/YSM!O35IFTE!-Z( 
@<X0[93!4[1Q%KXI_GM\@,?:MD]6G,CR_.0U9#4JYJ<X 
@U859P"6(795Z"ZO!$/+\)<OPQ<N3:E^ 7PHEO=\2X'0 
@)J*PE5=F.5XVGK<\0\$&1[=&*EB11*\6=X9TM3_EKL, 
@%\;,'A?5RS_^9YL(26Z]),S718JJ=[*[\,RS'>\:ALH 
@0=9J&0:?44\]E1'T/:EH,S%._N@ F>!PO+ADGD7P;8D 
@HS"7?N&624+(UO"GUV3X_F'A)G2__5E93'3^$,EFS^( 
@].RI=P]ETR\J)B"Y&/E'8 G:QHG>U@Y<%EH:E!X^$;  
@Y<GNTAHWBIC3];D+7<>B77BO]*0UV&J \_)R>=GG51@ 
@.S,2^WUFOH?>.IRQ&4$)N.$1R(;ESY59+/]M[(M0+R, 
@3E'PIGE-S:U>H%OCBN9,OYR0IK[ \DWOQ)P49C+OW(4 
@2UCO T^X<RQS76-^5%<RV^L(#]YD-[GMQ.#P1+R$I)P 
@TAL?:HIO(%@S:&G:2M<"[D,QL7PI=Q2A2.\QVMAO6X8 
@!H*27 O0N8- *&!YDM*=*-!6IVXCMY<>@V10)QKM8:0 
@ JF?&25?.IT#Q>QS9J77#FVOZH>%UV'D#>DCD0PGC64 
@G1#[9%A'-$PG4T(2_+"- CF_G%WA(Y=.-NOZ>EP&=[  
@LH9>6C;!5&>17: )8O75B,:]\[/27RA>'^TC,DNT\G0 
@O<J2-)FAKD>LU?U>E/F_ES7ZOV+X16[T2@%/96[%A/X 
@?2N$L\7.C[JOKMN74XOBH(>Q27G?HW]A7<XF:^I! $D 
@,S?T=\7TC(;6'5 &.VH7?Y FZSX]-*)S*.P_3^=Y] $ 
@[<0]P+@GM5$(1#;!0'JD7@;S-YQ(UL0FC0-;8NO!VXH 
@K.-6QX:O/=B:K7'S6[RZG_"DMX'N68U9HE$*CK6= *L 
@EW$1RL-19#K@ )'-LHH"_(&'!K!_F-W."@>O?X9J*[  
@^.$3[.I*;[Y$1;F2Z:S+'>U+8Q9RP>(2?W90L*MFGYP 
@.\\0A_S3N=ZZM"WZHS ;%L1,=;[J.Z'GWX9JQ&:S9(0 
@ 3T?9YY']J:/[ M/!\+E.I5&6,UQ5TUO:[8-!J4R"+T 
@#_PPV->ET#7?L3U;-XL>9^F9YF#TDXT05\SM<^2%",0 
@72+B'S2DG@&E"QDJ5SYQ[.UA'%A#>[Z0$GJ.,7 :-L$ 
@1]AKN-)1^I2(\3/926B%P$1YOD[!(*#05HWW<ZL2%\L 
@ H (V,+MV0VMT-B!#R2J\&C '0ZBGKPPO<C OQF/@ZL 
@NK#.AP4+J*1DHJ\LFEG9W[?<S$Z;LZ"U".W<X!;/)$@ 
@I6K##1EH@J]"65<$20<PA5E@$9%+B%0+DVW E>DTA#T 
@WR4K&W?%[[D8/=_M9L*W+^T5V[*N-?,3\EKR.2%A(*T 
@5>6^L%Q'$,#AV024X( W7EXEX*W&HZ]3')4:C_ _OE\ 
@9P6+=;-_ZV3[/:_!(BZ8" (2YZ&!%(L?BL14Y&3"Y?< 
@!0_+9E!)I$#ZD?BW0$R9J(:8M5GY?IH^+8-1"^E0/P, 
@5@;9^ZYQN*J>1J1LTJ7>;FH:W9GP^7R&U]V,YV6T>08 
@3.8#J,3J),<892HD0W?6%8F9#CNC-;ZH/DY&,>79#_( 
@/U' 8M=NL=_T!BO?ICY@P]I<NRDG_#.9X6MVC/D;9!  
@4AK :'=<0P>K*):.-WY%!N BK2&KD/]KLHK&S1K(%T0 
@WT_EF9>CX8=1QV^AV*]4X^R5,FDH5?A!YIZ\AG2%AXX 
@6RNGB?8,-D0R_,R=P(+/5_,'J..8"W:O69%R1J''[WH 
@'L\E:D4JP>ABK(?R;94]LA50WF@2AW6T=H$:@ ='GL8 
@5FBFSC-1:Y)_(5^RW;Z*I.BQ;?M>7@*8V0M=WM]/0_H 
@TQMF3;XA-802$)*;$XPXB@._(0[WHRUR[%RX,85C[+H 
@AZ)>9^@=&"N/8%INUV!NRA7D2DD?:H?0UF3,)ZF2ZKL 
@F<>!T%7H[XSBYA3P&D0PJ'=.A?6,*&#ZW[R8R;!$,>$ 
@/TO#GZ=ZE2^MSW)M[*AX.(&N,2</9;/J/^<R'8DN; D 
@Q]E.?N%^\07/.I?X>1;+U[<?G"TT?J:>!"-7VQ&F,&P 
@K^E2?L+XE%[?Q:E4F:S$,1F4]1?6#\9X#VXHSM&:2?\ 
@KG.0V>9>D'*+ QYSQI/&MS+ZL:HDHO*M4,OM=-%:]$$ 
@,]UBVO)759.G'D@*699EM_UIO4K7%.%/*:49 T((R(, 
@L97M$C//70;;!-[[O&\!4]@_X<JG?LL,\EN]2;#29>8 
@!GZ%T HF_8N.2Q;KTW*3)T$TSVUJGXQ$KS@L:,]*/5P 
@W<'!EU:KH=KC)>[X+^NXV_C<<Z:Q80WK@U;B$!=GMZ$ 
@45LCNZ<VEK,GH+*/R-$ <'1_0KV+'!2UJLKB1F$@R8< 
@,\<78V[;S#"]I!VS&87E^H48TJ(<Y*Q'%D#5 9T8_S  
@95QNJT7%-X]*F/?!PH4?5-,0Q"*9+_68S['%(?CVK:L 
@&R^ 3.\7:U3MLF,N4DU8G4V\Y8(5OJ'@;I="><LB;?P 
@?'@D^I#(/\B#&Y]J>A5')# ?N%:=FSLY"C4_+YN(O!@ 
@D:39<VTG?H46-NV/!SO8S]7]@-^FF=*YX5L5H[*\P4T 
@44B\ZRC'22^$$UZ4E:S)5YY7;2 WVJ-I8'JM[LFVF_@ 
@*2F*+QGMO:3=&%X5.1\^UR9-[$Y"MKSU?@,T@C**4^0 
@3+[H$OAX(HZ;"07..P1P25_XZHZ*C;DNN%#J3>6GAYL 
@DLJQ'UF \5%VIND&T=56@5;>*?>LA[<E:DY S^6: <T 
@BG@2F4'3ZW=0W"<YKZR3[1]%??U#F#:)LW]/HI<'RCH 
@ITO#!<CX(VSUXYF[DU<\SN/A&2UH!>6E8,)J*$7YRIX 
@<]#.17<VU5,[=D9L.V=6S3-\G]\GVQO #9,T[MD-WU$ 
@&XC)@$P9FJB[-<RQKW_E%0$/(^G8Q)$)'<#?*O$1@N\ 
@:CBBU9X7_J>10QRF8D%V0I7GE&!S3YN:J;=!HAT_*F< 
@?\VV$]*]^B/95[8NG#JEOX=%!1U9.L22WUQFB,2]ZKL 
@?KP@-Q;Q_3??+B>2^6^M'DO((9XU:8U^OS]_YSA]=O8 
@#*@84;:MB5#)J=(\T2,:TZJ=8F1[_!X^703[2::3Z8@ 
@9]>0)<X$4+,10:7P>]*-=O.GU:!S?7XOJ#9MWD=4!V@ 
@?KJ8JTFDP%7SZ!MAQ.2UEI27*;OF4 2A:/R-"UXQ7:0 
@8O2A:U_/E;QI1=?!S:GZT11'Y'$HN:3)ZZGCB(<-!W\ 
@);NC*E>(V:*2T)70T _2Z,R/_V-+);=1-B4 !"J7SL  
@:90X1M90F&%_ ID1WS 431@Y/3^N%:^<^I1!YTO2BQH 
@#CI$]04AS*;HZ#BR1L=\L]'.7RI6#XJ+4(I<\)OT(>0 
@]?G!PQ$5 :.R[UGML2%KX>_ +U?-Y9*["S1C3[((A_H 
@G.N'O7]:B*&XK?<VH8B:;C\"E@4<FC()Y'$G"XT4\?T 
@ @HQ@)R,A%%DIDR >U-%Y%D 7V*%ZH&JDU,->2T>V8, 
@1=Y)LM W2>!*.TN<M*O]'DQE^EQ3S>(51E$[#@CU$JH 
@8*RWQG:!A[QO>G%K_Z$^/6(8GX*_:7J^O6\.FP.+#J< 
@8W8M$F.PEB"T 23%).V('.=P)$AW19ASPE3N? EMYL@ 
@[YS^0Q13Z8J4#18;AG\DWZ%9!3J;:@:'8566W@/E.HT 
@$M)_V[2S=88<Q%*#/N,*G$DMH1^[UKH.H^"Q =0MPQL 
@1VCQ]D"*8 N,4ARN%(K]%6:/",:/\+N+LXE<4A"$!T  
@L@)'E;8OXFT+H@!RT5JF6BF8@!'W^(_G[3(1*W9;]\\ 
@%IG!0MSV%$#+US;,\D1&2[7M)6RZ58)$]K9:XK9N_NX 
@L14*E@-.BD 5D=5/BDEE@,'T(9EK[=2MS*"L_/W/I<< 
@0\A,9C  0C:J,"<O&/!B"TVS(=.3DZOE,M>7 @WYLV0 
@P)S7T^2O>IZLV6*H"\C^Z40U\O16L KX B(JN6KK>Y, 
@IZ5YW&$LNR=H(T(S.+1IE]:U2N:QW[MSY.,LX(V'PRL 
@)N>U ]RB:?GF2882_I_F)B=Q1;(=DWF?Z1WSO1=QJE@ 
@PYE"BHB"#R1 0"NI.FH''#$+)4"*UK=IV@PZ.%D\XKH 
@;S[JBDDQ5G? 4=/XTN_^;*^AB)>J[3Q2=N06JZ)_'<H 
@777,9#UYM(0PIC^_!Z#J-/U]GF3'MX"ZUZ\6J@6U$V0 
0[F I13W(>@ 'F.V8./:YU0  
0HV2J"HH<#R*RBGF-2Y'M'@  
`pragma protect end_protected
