// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H3 C;1%@2-8HK#_A'ABX4DU(\A+<^&,\9&H]<]4F\365M:QK;+NL7M0  
HX."_V7./6#\\N,SM5%1*N.W[G/I0F:>P3'#E[R39\$,2D_6,#AG!3P  
HJUEG!FR94./@/"@G?@VWT%A12UJ,A*!#]'.Q9A Q40\AO]4YZ=HJR@  
H<<YK5\=H49^E VL+G2=;Y& I[(.X$[C N*W.!Y,@C\2Y(5?X7C8WK@  
H1E_!(JDT$TOD$X92O-14-Y+I#GCCF5<+LCID^&-C7H/N\TS4Q5U6J@  
`pragma protect encoding=(enctype="uuencode",bytes=19536       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@8"EX[-B_19);TTS*KZF>JS<$3J<3HBA#?&4*#VP$*VH 
@1U]Z>PDO[0KX%"OLW:CXQSX\N;Q<@48)D1P_2+HEL8$ 
@^[E3=7>)1\4J=[SV3(-HEZ0@UT@5.IRO+I%-N+([FRH 
@#?FAT:%09X5&/^"MOA+1AL$9Q.$0P$'BN1X?0HRT7%, 
@ VL>MK);D_ F"U,YX=^B+B]N)%)47A *F52GJQYB7'D 
@.'.@^X)%9I@$[^G!3V>-8\ (Z5\B*?>]X+PEM%XH%&  
@QT!)NJ6=AHJ6PPT#_H):F2J/5F>2K0:V@O+#@,)F1/T 
@%\&Q9:F9\E!PH"CCXU8)6$XH=)*-!%]M>]AJI]0DE/, 
@O-HE0,W) %+K@%HU'OT3Y8NLNO#!;-^O0)D@!O4._2H 
@:3PW2/+09."U\!YX*6R=\O'W<-)K-OKXQ&DELXZU8+D 
@:2)_.^3\$TH*422\'N\KW/'' R<GR"S;BZH.$G\R"YX 
@.]-T'M9,P74D1#X/"F4Z(4]F'YT#@&80R5.*8=$G-QH 
@,I(=E:\;SHF1N?",>ZTF4"?W0DQ;Z(Z[53>);UF+(J8 
@G4$)%UB5R\OP(!;TBOJ)RJ>&A$O+U(;L\^&ZY+UW%FD 
@D69C@<&\\\(\TP/<254Q866E@J=SWB;&<9E,5H)VH]L 
@U>.C+("E#%&UP?X#DUD[<=B:7R3X%4*!NSAK]*@.6+H 
@H)$#Q+N+Z#L4\1*(MJV>]J]UIC$G+'$!OVT*3H^>,)\ 
@GG'GAW#&,:-5M2H576'X8DF<7S-W-Z5TS"BU05JF!$D 
@I?$,>3YLHD1_S#%5^&MK6@GY'UFKDLYX[X,4 SP$WDL 
@=)4;;[_D]4GQ$M.]BM=0(:^W -L]\W=!4%NGT+NOF;, 
@6W6>4IR+Y? ;_P31Z%C U0[-9YG8A 4S)SY8CG179W@ 
@N3:18ZFD,(= DUNQ=\/?42B+>M579RE0X\$TFJM\RP\ 
@=0OQKPUL:@#^U&"5B"V^Z)ODDWJ@T-O]DEV5$!/-&/L 
@?I0.NH9&E@Z$-D6Z>5JF/G4RB!6BNYS/<.!8H#AAK=$ 
@&A13?D3-F0I( P>M,"(NA55VSZ>%28YD @3>N"*O/J, 
@F"0/%"P3<B%J4J9V]JJ&2["<8HEM;<*U=08"]@VW0&( 
@V<\F*I_52L):5W>- TPUU:S-EMLZD_V#U1Z[6",W3'L 
@BUVJ9I/C^,CA&3BA=D9%U?]RDL<VEZ5WK1!/G"J%CT$ 
@!>01R:IN>9T(:]]93[RX^V>FY<L9?;$*M,$[.Z)EP]X 
@[3&F%RD:86<(R>L(;"M"?*HGJZ<4?B1.>6-&&40+UOD 
@$9!\UI^(%Y5CUJZAF_CE\]>B;B("HV:=*(L_S(Q*%W, 
@'\Q>:0B)./-"N\=E83215=4E[7RIAU$!0%M@P>L3IMP 
@P+L!G:<0NDCL)%A_7*-<G;E',!A$PRP(8\"G,50"2)$ 
@-IE\T%_9'YR#1$6-_*#TCL^\(( P & _7UUL1?(#.!4 
@E 7Z!+7E;] 830^/UFR$'K>6F=(-7>^^D4+7 2S@Z"< 
@BXH],UFO716YVK0O<ZL)XJ5^Z-]@! (70CH2ML8M?3P 
@%;Q"T>X  @^:_D6':BAUXJQK97T+C?#8.'V_W7/&L,T 
@H\^E#$3ZB4JH'5^5@@ZXF\X9)&E;B#(3N\)7#./TK.D 
@F:-^H8)-Z!H\&\2/>)FSZD'6$D#",521_CTY&)BS;W  
@G'#@J4UIXFP0V6/_P1&>YTV)$_'"8-2T6@FCU4:>&1  
@XKGW5XG#X\.HR31-W688H+@6X&4\9^S,&5<E]%0DHX< 
@6\JBZ$]UG,$A'^=6Z@>0GUAC:!PYW;^R3IV?L">L"-4 
@<&(%1!G)$,@^^&PUV9ZQ8W32?)%8];]&]7[\V]=0B;( 
@ 68A+:'[D(4T:'>8^_=UZBY ,5"KS*:+FE'DACE/H?\ 
@$L&&:\*Y$YUD47,MBNATJ;G7S<'68M7>=DK 7.@O4KP 
@!P/J<"Y0Y*#F7.#5P);JO/;.8Z+;..$R0)FA=?!X6FL 
@%27W*K+6D$]""F+0,;X!)()+MT\<^TO.U^'F/)M[+)0 
@(U*A]$,ON*MS$+[I9<+=N&GP@U4>/3RH%'OY);U3'/( 
@PH3W3;]UID7[D5-EQQ@3JXJ?^LP?E0,'$<H3\#XO_U< 
@DQ&;77ZA__)\DH%R6-O*CF5V3P1EI@A=1X86J!6T:#@ 
@%\TGC0WH%"ZLUME;7%\-B">E^5GZ-SYM+OC)<'0*]0P 
@]V(X\6 $2'CX>C %YR\#0OL1#;G>*PIP<P!O(1A_FR\ 
@%13)Y#K(9,'^NM4WDD>G9FK07VZ@*$L^2@+T^*-',8  
@XZY5-59^J',NCZZ" =PDR%0)11#Y?E["87 NZ(GFP+0 
@0 TS^0>(LY]?2%GQ.G9J1"M&ODYT:9$](VN(]).2RDL 
@3^P*'BXD!>H%2R9L>=5(2Y]RVZP<3_>5JL,.+?K\&_0 
@>OAOKP^%^A]TMN$3-#ACKW6&P(NTF4>Y:.V7QY<%%\H 
@O6>&;8YNG>;)@!4K!%EZ0!*G@@'S8Z%WSTE;+=_]&6@ 
@GRB6-OYI<GQD']ER6",W#=6:1'?T9WWY486B?$%SJZP 
@>Y "2L8'"L\):4@7ELTOJ"$95H208GDCUXHRJ"T(FNX 
@F\,,?F7$'AN(_Q+RQ+_PW+JMK MI=%" _WHYPYOR)X\ 
@BQ^E?CM8"D$9+C"I3QO6MITXM!?J4M[I77^-P>>B-)T 
@ #S/*ID1@2L.A; NUB:<>TY*H+*8I4/TOH_&PON 22\ 
@IU_7#G"3(^J2=?!>KRGG DO7<QBC@>7FV=ED:HSRYMH 
@?'V<55)Y##W(5S1R?B$>FDV?;M>2N=B@',=G0--1!X$ 
@)6U7U#)ASGK_XPTB@"\XB^(TQ2!/W[# _,@&0\.-^7, 
@VA!^=V=T=F?=Z)L[2B('E5OUX&DYGE3=.RNL(;P?M"< 
@4]1 4:+^0+.F32FO7B 1YTY$*9L&VDS)[4J'C>S1Y\< 
@=XG2W1A#'UFYH6UIM$=Q(*U3[) ?]%6-'*U8.V16!70 
@6OX^Z'#]>,7>;P3X?\C4C@0L.$P@@+D\G+)-EM7WF%@ 
@A^=[XH2AR!GU#983C8.9,1J#15+/2,O.@_JE-A=T!QD 
@FSD)KFORF<?J,?=%]!V@"561QO<4V'@'F:O2"O(81,4 
@DXT.IG$<N]S&3>5S!960D1+8\]'D5]=<*,EL.07P_U< 
@<.1&.1 HHG$Q[UD_6X\8DA.@H"F9 %;8=#FFDZ60W8H 
@RZ:<B0/KE4*[OEW_]K+C^@?1)O860]EDJD-M=63R*X4 
@P<2MZ)55<+!'0/MG+L(C.W_A'_L!6A$<O! [BS_--$\ 
@%6+6UT?Z*^+)T\4(#\*K]DWF$!7_  V3/S@QB"U]ZA4 
@I"?RSI9L&V?RS_1L8*71^6A:$S/K%=$4;PHRMSHM=Q( 
@:QI!<F_MF.B+0&N76M7P'V>!$\X91_/WQ#XL-VT$*/< 
@_\!<*S<73_NM>]""X=YXK:WDTIW&[UY8[&(':I&CHS\ 
@C =2Y"I7Y*ZNT&F2H)8*(=%.L6%<4TX#!^X7R&[GCJ, 
@OR"$"HIH/UMAG9O#^NIKA9(YM\2M%RRN<3-!!U13JEX 
@R_/&RDF6#%0(%A:V.3'\_^I$GV79YMPK#*N#1=L'M^4 
@O'3*[ZA09<E_:7U'==U1N:.-N9))-^W=4P(9[K0!F5P 
@]\'H;DPU%B%(.$GJMDQ-6'6'GSFMO=<Q$J2>Y["MDP, 
@,OX!S/2-HR<0E>B7O\>@/$OR?"NE#3+M:]Z.(XRJQ2X 
@EH8B>U#AO\\<#P#"AC(E[B*5N 5MZ94_5OP-^OD 8\8 
@K8$ :4?P*.V7HFUK/6#LP(<1MC$T0C(](?7E$V/L%/$ 
@?AX_71E"4W[I58'DJL3E#MZ4:< QCOSAIZZNG]0V<E( 
@=J%B&^!NZ5DR*/B[-)\]=[5(]GC"H,XH7XUZ+TW9" , 
@:*[0>BR>+L4OX<G!?GLRA3;$3^P+$&]''Q\V*LMVYC@ 
@Z0['0-_P&@<KT#X>Q;&WW<9P.]9KU<?V:M)GX]'U@', 
@;W0\!LW]))L3 \()\!ETC6'=-!*]Z"2,8))'O&OHYW8 
@F$[G+>RUN"\\F?33)SN6LM2YZ0ZA.YBT6?%G*)7I87@ 
@C#^_EBP9G+')YU(*T*?)*D9GI8V_WM"'P.(7?^PY>I( 
@6):@C('=UW^YVG)N+-Z8LIK9(@\8&&JR#%1[KNC4EP, 
@'CJ\LJI\\,H03G[CZ8]/WJSG?M@U9>-Y+X@GH?#L',8 
@=>_^N%AULK33QSOP<QLFN&7? Q_5[FY5M8%C+Q<)<L  
@_"7R;!1-9HG)=I+&F3&#OX*&T_\R'<;Z>[']Q,L]E)< 
@]VIVF"S6#+#U+2095P07=3RTW.1IU-W4;ZNXJ&DBRO@ 
@DY-!H0)L<\./2-.NB[\YOVX]7;P?HFVV2SSY+MF3JA8 
@X)3W+ &A,]!>+]WYF;OB=1@9GP81;3.?2OB=O#CG6), 
@6Y#WM7H93\4C-BS2BN34U1KY'Q*)RX!LI9(;<?CS_Q< 
@16WQ<TLM%M-53!D:5(*KN0R&R 9*:O5PBY:O,>FZ.Y$ 
@!C_[_EM"(*T=,X,.8\CSMNY8X:HNMP3Y--0CP/MOD4X 
@A2K!(P.4(A.'1@G%P@=.U\Q <#%14VYJC@K;F>_T?.< 
@7TT0EG<W'"87JI<P8QB2-Q#'IDQCIZ#G,,]_E3>/MAD 
@ALWC8_JOT&"WYT?SHHE):L//5@=<T>/O1YOX"*]#SKX 
@\'62^#3-UD$4HG U-@Q$UR(22C0U7$X&L_7M:QTT%0( 
@B0VVP]B&A'_^\)CVJ8.(+30N8<=(H-5&I*)7%Z6L-BL 
@-#@<0,.B1!E>GKKJL?/Q%\/GSQ,C>>?@7<_(T>)7JWT 
@:I*]K<H/8A13^KKNY:=  :C/?Z5H:41]^8 SB $IF'T 
@M(#1PZIPV-,X( N''=LU:.C%1N5(O%&8<I92.C:W<PX 
@UWKI0P9=QU!<'K.9_/IBKP;'Q4?R^AC=(;TG2YRMA8  
@F5YH]\H*3I[&#0CNHET,E$(B.SII6O$7FF/X!UPYJF8 
@OU?#9W5TX\8*:]?#!;'9PL3;E>0,%P&=E*25K43U47L 
@<]U+]YM-GFRC#% 5G;GUJ. #)OF.%9YJX<YB!:LQF=$ 
@[D.LS'&0!%I%CHFIW2HAY(BZ^KBA8UUX9$ !FA33M]P 
@O-V;W&"G(.9G6C:9>=3S)'K.\R8RO!:@K&$#/>!Z<\$ 
@Y5%#"RNW-D/GN3[F@OD.'1S<)ZXVP-\8ULR$F84A9^< 
@Z:M0[@QFE?>'Q+](Y#KC:3F&5-?<C4O= 0W!#P,!J$4 
@/M_I!V(>TN%E-F9R]Q?.QA0J7F8OOSU6HZI\C&8 G^$ 
@D62+"#?,I3V%9,Z2=AZ75*Z-6[J:5<R[_A6T@"01?7D 
@.=8R4T$F17N3)SS-^,:83.MZ?+M5/!M2CM\9@4U*5(, 
@H]+$GRD?_?$O3$R.SL>83GG7RC1[2V=ZUWKK, N:?+< 
@PLE+*U8^JZ8<6CX"S[(\6M8L"ESTC(8V"-7LGL$E'_0 
@T/5+D1-.C=?6-?]H>G_ID>NYF7O:00!JJ79$KTL#R/@ 
@$#(/P,X& &9WAM$QP=3>;A9B")A%3/UL1&(&)<F^L74 
@)AHGV)L,LBC#_/F[W=>E;:0J"*45E9 )"[;\O2%!$=T 
@(.3?4X/5.D1(2S&DS>]K9-E;=]/G7T@(+OLKNA0TY-\ 
@XW*^6C,5K2)Z;4E*5P#H4GW'SZ*/:$!_E#%5'+1$#(8 
@C:<2^G*M8&H$\C402':Q87_*44_@G^T(Q7K0(\!2 WH 
@T@\P9>\.8X?N4.:@O>*F9)+V!2J3#=?M\Z=Z?"!;)K\ 
@#Z@N7")NVU6)R4:2EPY1E38=K(^#,16B%3!%+#(@2N, 
@L? TU?> 4QFW%)&!'NBM[0!>:UTI,AT1&>[-9(F8[P( 
@\!1B6H)A:K,AWF,V14()S*"">VBC"D!,JMS_6W;$G4L 
@8><H9TC-,$5H)-X'5B.M$6WA79#(8>_'0#&'M/W#6-4 
@47(=I_V5(AO6=CJ4K])2U-I*/<5PBIO\W>C\W*8%MWX 
@_>X2V5AB= P[YX[D"X4%%QIY1 X9D@H-XM_6'?4O]@  
@87M=Q?K?TD^3'G*0_8G;!/KR)8?$B*!)0RR'50015.4 
@8H07DN" Z3.K*UH'6>%6XKL9Z3>-(;3#(V:P'+;0HN  
@2#I,1__""/B,^^2_7;/CL#=A;25,'R(/ZPJTA@NCEYT 
@#D+-38#S%H;;C"0/$ 7UVS=FK4QYVY6VMK+ FLQSI'X 
@84UUR?+^F##YNX3_%T2]$A,RD,_E*-W?DOFC>6A2Y!\ 
@CFAC,)=)LI>8M&.4#S[+&R40;L%RBQ<1I^A55,05Q^  
@:^TGTI+]^&V@CP9N\D)$-KU5<G22_5%2SY(&$\%,AN( 
@]*[Q!8?:RXLKMD=0RH=4>8WPK!63SH*K ^ K;3I'S/, 
@Z2J#WO 22OCL)I1&V.> G\A*ZFF+U)TF<V+A'BES[L@ 
@E\R_I*=$OM/J)[AI^!,O"H:G9U)8OD%.;F;*L(!"H<L 
@B"=/GV* .8_[<2C_U3$AX^XJQ;./2<=%2=% $P17!-, 
@E$\-$[NF8 -;=QL+9$KCQ [>:-(:B'I9W]<."EXW\*H 
@O^;^5F@(!<!1"?K )[A6H<X6#VIX L++G+#3[\=KX>< 
@6A-33];Q?\('-20G<D^A ):2W<CY.H0)/=^@6.=&]+( 
@ZVIQ75?&<,S>;<'*#2G\V4=$ 3=A&X%"J69,*=6VRSX 
@/=Y*/.4H+Z"/_R$S;[9"R#Y/D.T9A#(USUIQ.SG=T%4 
@5B74/U":)=[7:0K]4,EJ;N-88IPOQ@_ MURFW\T3+E  
@K#("^U:F(9Z\Z-=&OQ:+*<N-GMT6?0$*'D4[&&E$<&, 
@R.$-TYG)\Q4 3/JPUD/;XC'$$Q9L%8#RT6Z==R!B7WD 
@Z&)Z4JVP&9GW]9BXR3<;QBD;MV?>T_R?9XXOKLS1ME8 
@;JR,WKS+JYE!&8\CY['N-RQ<N$I;W]Y/N]8%9-T57PL 
@,3*=KNBG.4_SWLE!K@:Q3>0#2#%877X*@XH%V4_,FAD 
@3IE4T3MU*%MM<@^05)N.&ZT;.G"V3\<C-5?@2'6C]4@ 
@.%"P""4Y!B7\_-R<H,XM<]I*P$%](<O^%CA,L98GR4L 
@2+A2F-];P ($ML4S26O*8A/;:VN%@<E)^655,GDGON< 
@ET78%R,:_YA[ 4A1[UKO*GCMM0-6(HBQ"+;&3D)>QD4 
@;['4'8L1B0'T+%;'5Y/#W_/43\+G\#A9K<WQR)D"DP@ 
@Z8> N@%%;AJ<(7B/3M?;:1*^BET,XQYO':20%"X#IE\ 
@HE"I;+//:Z6')VZ7%]HP^#HS"F3TF!+>'89^6]]6!1@ 
@SB#$S-;],<M4)?&QBTXW8Y^5D)F]:TK^C(8$..X\F&\ 
@0T D[03O$:T3W$23BUSMW4JDYLB=U")KF)M', B'U=8 
@8316A#5PB[V*(J :?)"Q:8?'_EM"X<J!]#Q<XEC(/?H 
@1K#W]CH4!K0\,XV6-K5/$81.<4.I:)O6T%A9^'A["Q< 
@1.?;%<=)[Q"8*B4E47Z600S49T2L[A]/E$1B3&+(=5< 
@M2X.QO5BI8\[KK(2C^5KZ(+@",DI%I=FCPVV\JV:0Y0 
@+U[(<3T( YR\)T!)S)'*)W-:WK[5QL4T\7'P=BW/G^0 
@LP5F2B(3$JHF.SOJYK>F([+8SP0_3R=8I>Y$YCD2C)H 
@)Q9B>>E'\9<SC?!-;V_NW3 T_=9]W5E_JCB7I+!43NX 
@_ 1&CLO@>;^)V;XZTHX_ 4!B R%_X;%!;&8Y :[SG/@ 
@'!G9B[,M9,$$!"*0,]-.222UK04;)2%<85J'(%FI@QL 
@1DFH7_"KSL(-<)TB&+G0 J -JDY6Y-]2:L8"DP+C :X 
@AQ.1<%Y^OK<O+Y5<UF2QD"AI,\<SLP P8^-7SZ1:>)4 
@J_!@975_TQC-=8'>O)9APR"C_YBR9IOZ'4<(P.^1'-X 
@M#RSKQ7BQXC"C:!7<[A'N-)R^B&F$GPM'P<&8L)*;-@ 
@N*0&>DW]!$%3G@MN2&&QDVI$OMZ_2 2IWS'CL(%C-F  
@W5H]7Z3GNG-.H\P2:>J],FASFFP=JS9K]^^2T3$&"EL 
@7'4/,(LVV FW,EBOT\OHQ_(ODRA[:YL^LZ\)6EFKI/D 
@3G(C5SSAJPN@SK]3:5N$< @CAGF3+O!'5;;#DCL7G4H 
@+MC7RP4VWJHE9,7#M2P^U<8:YX!*?1J/)18]/[\P_1, 
@<(].OX!=4 DRGNZ H\DB-YR?3J7T],V<ZO/*M,3FZYH 
@8L-^4+.+C.0!1"9IXY)/KE_=_0GS1)E<&E&6WS/=P\$ 
@_HF2?FE43DADW(H(%6 Y4&$T<3RMQ" @9KV>W\>J6/\ 
@5PDY*^<S%4!4%R_?Q*)P3!W41MXU-8]TB\0PAP*"HK  
@2+@&!]GQ&6S"2N2"]M$"OH2?4#0Q-IPIK!0?!$:W/V$ 
@$R)B$G]! I)[>99)#?L(;=-)/$14V"*/5[H*D(T4S X 
@C\)7M!H2_$QMD2H_=QO(9@AV9J7:%DZ&_!=;D<4)F7H 
@HS#VY.LV;0[$6(%[ &L0X3&[QZ83F3X84?C $G)5M"L 
@K 4D4'D5H$!#:BJZJZ+ 2^<>D1&KY7C=8_M]PUXLG:X 
@Z7A2POSHUM!]6OI;ZBVNGN?^ DA9?L";O^<M3FIL&:, 
@3!68-,OMQ@Q\H8T,ED&/#V^!!;(F#:+3APJQ7_$VD0L 
@Q;OAU5<QJAV/1(YZ> /XRV@F0A)3KQQ ">V$;"&I>7, 
@BLXRX $.D;-'K/"C;='9'\&-Y0Z+OF*R-P/@OTQ=EAH 
@%S'M.DBA%;-VH",%D2N@5O,ZM76;=&WJ_[KOBCPS+TL 
@T2I%TFH[IR]PH3X/Y0[A2ZZ8RMQR<IE*6@F@LL.'.5( 
@=K^J'!=2PE,\$_D&A!52!SN;@)8" Z6G9NI,B69^.<@ 
@&O=4=@8J_68.;77H:(T\4('LQU(^V!E%]-",](EAGW4 
@R$/A87=:/N[4/T6+;]CZHKX?ZZPE1A@BY-L')'/I-$L 
@@B$#>Q-*=N 0'JB<[W<Y5\I *.P1[=?/K-1&(D^/ "$ 
@#A\G]R0;.>BL7+W1_?NK-Z!#479)T])B%6.7Z1:?N]0 
@%JI&<4^Q.E"8ZN6X R,+1F^5H N&()/D_X8Y]H9@P<\ 
@Y*61B.;T$U@G<FX0,90"2OWQ@A+,.':>12BXJ6,K#JL 
@#]I' :F0(E_4YHYR#M%#,*.J ITU6M+.7.64DJ#1MJ8 
@O58_.P[DB^N2(+T9L/8)K4A_U_GX,$VRQ"?K3,#H"=8 
@3M*,:8' IQ_ D+.S@MFH^VFI]Y0%C#GK":881H1'%4< 
@//6)91O**GF)#O@<HQMSF$7%83B<,:#]$N*C 0#A"ZT 
@(D8&E;FP,Q<1=0.]L?ET'&5Z3@WD&N+ELDI\>\?]+X0 
@G\F9V3^GED=.I_:#N#)'5'XV#B1<EJ]SMFN436A4@ @ 
@<2X[AD/_W#=#Q"&0 T&\&=\)!LQOT0E(^HI=)4)\V6X 
@\31:V3CHK',CJJX4+F %HF+"3WMMMNL'XK#N";I^EBL 
@<NZ-A]]%9\\_AS&>K@_?IZK4I(195J)T:8"4?U[,UNP 
@)KAMTTT<L?]L&MY83Y>'&>4$C_&(&>4=\/])4V^4@5X 
@=.^44TN*_Z=VX;/2IS?Q:OF2W&GD=6G?)U\S<81\Z?X 
@:(1: X-Y#BW]*$Z\./>N/:AI-SV<.:(86ZQF*L?][JL 
@-8S=X!MY>U1T%UR*2VF8DU/BLC;[>;KRK"THO1M+0/( 
@-@1M;':TO7($+H30^) X)^>@J#/)%A=']=&6K%GG/E0 
@ZS/OX?A[(_ *[!WERCP9V->T?>]?B06G6 [W='\<[W@ 
@,POZ@Q0GZ9,Y.;"#"\K>,,IIU.8F^9:VE_,<5/R* 3, 
@6L+16 )[16#E@7'+;X'GW:A9*QV;6NN)Y'*U#D3NQ   
@,43@SW_&O%&6(F8ZP94R8P84P9?%RYS+2EJ?GE3-&L( 
@Y6H^G8R#1[9I_6DQIRE=T'S<>KFO#V2=$=X("PV78(8 
@W_Y/@HR,)XX;IW63L#F9.V3V$SAA""P<N_,V<QL]"6, 
@"9U$TZXW 8C>:56@"D]EF3P%$(\,L2L.S06LFK<4.TL 
@H[@[_^A=J)M%&6T9HGI)")0-?"I;9PP(P+EB:O[2W=@ 
@P-G$A#BEWX@O=.G5V@R7Z<[J 3JP>\%&36$:[L,6VM@ 
@H(89:A2S]50>+R3M8:NBHE/8:&9)<#8/Z$^0I"AB \@ 
@'[>@4RP!S3DS30/@R,W@;.X"1(V"Y80X8$JZ8Q'&(DP 
@KQYTA_AR?AC!O]1<O0&?K9? @B?NQ.$(!D9+)K-@R6  
@OMYWO1<&5B]3,IFCT.JJ;+OU)2-@IKIVO@6SCE>%%(0 
@*#MN8)#^UP'(+L!9<@+!Z^FZ9T;#^DR0!'[+746_A6$ 
@5$.4;L;?H?ZJ4F-JCV? !0^EUHF.N5X+(=$:H R='IL 
@HB71F? >PTU,P5Y78%\5?JQ8^-='*1?)?Q+:D=Q$OCP 
@@8+&LQAS7UO,L(2N_[QZ*S(=C5$]+K=76"T P:X23E0 
@%M0D?"<N72U3PBD^B*$Q1DP+U6'HDE;"5: IV]VJ[VL 
@5:7(+\T.Q,'/<8):F8Z1&R<%XO.%MP'PX@%9; KR;[4 
@V]OD&LFBHK'T1=(NR;=<LLJ2 +?]+4QF0>W0-TV*\P4 
@'#^FTEB@?/M^4.+[.(.<GNI]TSP6/;1B929 \ *)PG  
@"]#$C396+%0"14M">[[!2V)(OJW/"PG Z38_/Y !S%P 
@GJ2&A$I_$-U*8QV7$!5FC,UG/6Z;9X^Z!*' <TMA.L@ 
@=04M9S\'!3HZ,0P14%QL@A<U;BGD'@U4^:^B%16&#?P 
@4JP,#\8@:5BSZP@#"M$ZS=4]"I;[^IDL4[-'ML(^"V, 
@"6$6X9X-!=K))OVDJ2D+E8]^;;A\<[#D!%,FTV.1[<@ 
@X\AIO%E6S*4IH*37:X_//F6V@H0;[N1SIM/4#R>RQGT 
@(R.)T3V!]K4IZ5!V4ND#IF&/H3B92FERRM&KJ>:_NZ0 
@-V0#1!Z>[IM-@6\F)SD->5BWA-E/S*>*0:2M5Y5%HD4 
@?YDM55]E>A,XG6"F%!UIE63@9)QJNROA5%#@T^*$D.8 
@H=.^ @<.X<5%[9\ C<5BO]KI*D#D9O48J_]\/ 5TTX0 
@5#CHW>D:AO49+B5*DL9"8=R]GW05.Z;2\HONR^?#%44 
@]KJ_LSX&TL^X:M]Y5E,G A%^JJWPB)01;P40Q.!9&-T 
@^^T'@1S<HS.&.<V/F?WO%)O .>&/[T19\^ZGC-R.RW8 
@+?'Q,C0V!(L2?@(ZX'SC[]_J2_A+3G/-KCES$VO!^@$ 
@RJT0IA'[XTV"A-9_@G<L?$,E@GAM^]JO0X/]S\Z<RZ< 
@TC3+JY=.Y:&,*T-,'>\%IF6R!7CBC>\^#H _\593P88 
@# IYV5,NX;194$ "(-L)3EX!.;U6)L,+;/SU# "]AH< 
@%^$_)6X(>.[Z7C:(<R5SOV,IPY?2I!>Q=RO)@BNT/XH 
@::P8%H%/]+A2V5\I=L^*K;' D.EK\[(G9-E.PU'553  
@S"66UP?=2VG:$?UPES9<>193V$K"R.U_"[]7M)] /I, 
@GZO!-'DSM/?^QHOW +8-C*8U9D HWPVY$78#Q (:E$< 
@/KSN@MCF:6(\CS6&>0WA1ZVCP)$31]/,,+8]$-;D-E0 
@2[@?L=^J@.O"<X&J!48ZEL>&+2"+3D@!W_Q0"EA@K9( 
@Q# _ZE0,V=RE-TO+?U/Q/*'9;R_-IGK..P1C(LRZ)N, 
@6BC1;/>7;&,SXYVY!W(9F4$U)[Q2-LRT"=<*Q.S\X24 
@H>FT /+[E*W3)"H+C LU6G'UIS*6VS:0J;VWPA5L--< 
@+,S<$O,R4JT4!'?7U%!NCMKION OGME^Q<5/T019X"$ 
@P8[->7I(^@?;=O34,&_9KZ+3X_3NC[N]W3/'0]JDNV\ 
@-II0$!&/PD9!3ORH3LZ,_Z:Z!VI:M&GNNGWC\$OF&8, 
@-U4FT1*Q $RN>L.<)$IRM=)NJE4Q''V8NY88\^-+\Q4 
@9FDB:=838NZ)7'X1]@@:JE_XD FU,&Y-[)?DXX+V/MH 
@_9K"AFK-$-B+)P($31+:V J]2OUOR1]C/@/G OL%.>4 
@LX#Z*_ M+1+E]MP>KG%QN9:KB5HK/W552'_QU?!L)#  
@(CROK47%ZY<?RU=4/47'1M8>;!)VH>)_7.;]64FG_Y, 
@F=>P$G#&#]">),K0L0O"]P\T8)H(9W7-DPMC+9^#E)  
@0E,M(Y.-CAC8TZ)OHS%*[CODCBW2P5^!O2?A_&MU$4L 
@=Q(Q=,7$&?>MD"71I4RSD( '@..=*8I)$:NZ)G&?*$P 
@BZ-@]U3C0-/2^GL-!4TV7?WF!&C^!IM=R!=Q85K@4:@ 
@U&EZ(T?-Z[L;]AYTF*JA)%^=R6QQ[R'/!1QV2!'S9Z( 
@[J#LLTV[I&BL2T3O,"D2D.?B+D@8-H9?V.EBPBX)Z3, 
@#*%=7I#0ZKO>LT;+T?@L&^R\H.8Y^4/>/&8R^&V<YD0 
@5A<ZG]*=%/N3&]A9+6<\JM)P0LX238.J:F7*6T>3W#$ 
@K8$PB%Q9,S$198-K2&XOG*1BFQP0\HYN[5/&O(@/0/T 
@Y$#[" ?7"*2Y@9,I7D)S_SN'%5J]11/^C&]U&\N;K)L 
@:1HH&#U-BS^CL>U2%_?'1 4BH$,%[!^JTSS.*>M#[_P 
@Q<-EN*)*I?![K;!T[)<2  V"8TA@]S)9+K7+/4H\:=4 
@!!';#RL#U3GH[I%'6>V+7$FZKS&Y1^>6=5SZ3:F99(  
@*L'-<]$'V48'UL;]4POWV/^1K1HULR(:[YW1-<[^*+4 
@MKG?JSI(;L70)2$9&EEZA+3FAO3;"=&[QEAQS<3<K', 
@<<-6?0"=<9P>!)5=,RMT4('M#S:A4S!M%B-=W;":7_T 
@_RO5>53E<*>3&@C7+ OOL^<6$[&^)B:AQ'S^9&QBE98 
@E#]\V\Q(XWX<NL?]D<E[63P@5GI\N&V0U;\:0[ZICO0 
@$)5&NF]8(T*K++5![/AR>%J00.VR?IM+ \A-B/ T&8( 
@>L_G"GWYJNVN;WYHD8!#(%X7H"RQUR33F*"AT!'S1,$ 
@%3U8/&W_$JACC/;H>W[#TMG;#[,;CWJTZH/O?D#HE3, 
@RX,XF=U*P.^?;RD,[->JN4)Z8180MI @U \?0UP9[&4 
@X/_7\G88D2!%ZXRGRD^&?FK3YF,P.50UF7Y-3Q6+F1@ 
@69G0(RN<!@RA#3][FV5S=A=X@T4SA20]IQ2_RJ;LW>< 
@\IE=)VC^3(!'56A9O@D2C%I"75>SG>>8V*0/5$,:\2< 
@()'R>2S-B]BHX,2Z+/N^S07,-CDM+#[&"&+"ZN&68VT 
@!/E>9'80:_3N6P4Y[73K">P+?@V0.SB HX8C\[DW^30 
@E07.&'-W:8^31^!U/P5'! QO\[=?..J(V$36)&>Z1ST 
@B<3K/Q;-&^'L4+Q'=#29%AB&S/YGW\79DQ*ZG+B34'  
@7K-S:+.\#P+.$R);6M4"V@ @Y4R6+"N]5W.6G];,4-P 
@?A!94>X:4@+"2Q=O[C8"P ":%_#6U)V7#O@K9:$R(BT 
@2G^YA]NS3LM\/7%_%3VP$VG*'9EH)+Y=(_'\NME*4WL 
@]M@9PR-I?OTPIZN7.>];ABZ@4W,U9RFAE8F+\+OJZ*D 
@I.EIT;!X'C29VS V7K1.$7Q]NV&2QIBN13Y-NR!UO^  
@M19LMQ&1B_\H$^-'9I9WP)-_H8HL;*JRZ%!OZ$.9#3T 
@K"KOTL]7GOP*-*K;&Q%"X"#P*7KI>H0&AWLPMQJ=E]T 
@?+3H1L6FE-S94VDT9M2Z=+U2U7L"*%?:1R"'-0$9VSP 
@*G9U0?1UZPW1H)?\\(;50U2$,*D *P6*#_&</:)=X"0 
@3ZRY3F1DI?]S&;BFY:2>Z.GY?']"E2:F._X"<X/$K*D 
@%X3OPQ1HIGGK(D=6'%5C\*T=PF'#.=$I)BXP,%#C!HL 
@JK=&_@,0ACNB@;Q!);:K]Z."EP-(#+T*ILT#AQ9XDB$ 
@TA-6*O#0X!A#@+FFV"TRFIX\?F>'YPJK+KA?PA'4A?L 
@4HX5V%K:DA^7W<H&L<%$L4F[P&5EBX=MB0]MNO/=ZZ4 
@; 9I9!96B4,M/4)&8&*O4+Q3S>,UE,N*B?5<N>Y(!]< 
@*K>+:J0#XZ-F0<9$H@(>6#DEYY[AN46K/J^-*_&"W?, 
@IR,<CSXLR]%I)ZNNR9M_O/Y1RS[[5JHOS*G-/MZH1/H 
@/P."9<G(379Z^-TX@$W^2EV=)$$\%7R5NV;C#.)=[>4 
@6.OQ<"N<Z)XRU_<CC][\$'CIU:/Z''X/5UNT>)T^=!< 
@(":"S:$WZH3_[G)\N30?#3?+5&ORBO"0M9-146+DE5$ 
@HGVD4L'I'T5* +4"%E_8V8WF>]7V1BI\>SGS_[C1-C< 
@2-A-86&JHHRK59>X^!,1-'$A1 3_;HF-B4$%14P_5<@ 
@AOJB] ^85X^9X)9+D.%U?'[@Y4X,T7GXGZQLI8<]6#< 
@45O#%[N. D57>W'6/@[(B_G: ,!K=;^M1S43P;K212H 
@.!@&-Q^Y[#-'LB8BF'\3,O[8C+T36R%1 T>YCA)C=D$ 
@QM%835-[_/.1%I:$'DV_<ZD$C."*2+HI6G'#3<O#IB$ 
@".<4OFW(^@U%DW3%&:$NG9,\USB3\K]'0*=0XWKVNDP 
@D8A1^+"*M)]FF*SY9K,PRP06UP*\O_'?;O*7!NK%<;( 
@H6\/O)S)Q)8F:[":\C)O,^TO#CY+37ETL0$YM!F3]P0 
@9#;O&Z>KHK;N<3U#Z5\V")QR,K_1$"0G/=:9:?HSB<L 
@\(9+<EU[-!\RB?[U,80LRZB!L%7-K]3676@?XGUN3G4 
@Z\Q%UB#<2![>Y)]WEE6TI,91IFAWE*87VGEIVDAV%\P 
@Y-Q3;?\0S\\9Q]+X'/F:8D @WTSEW_13W4[]/\GL_M  
@8=FBO^Y:WO3FC$'3A@IN5"*J@M9.(PNL$))HXGOF>P( 
@#DO#D#([$=!8<A4_J&G)<0_[$2@90&T<7+T[>6B*#2T 
@R8FBL?.H:*4=S4"=OM+#C"\W=JI77!N^1=B*O8<3A1< 
@XW$!GW=U&^7"';.#<8DN)WR"BBM IC1<[\60^80/5:P 
@N^RC20&35(&+5,3O$DZ3/I*8',/$8#TF-O2+((12'.$ 
@4H9_OM&A%Z2O>)>'%<"=!VLF2CX7VSQ]-0/!8,%%0\P 
@KJ#3'G!UOC&W'/4@*7+,C!19PO@R1=EYFK<)I]9*+%( 
@9MKTCO8$CAT+>JULZP]O9)#CFYBI\K\7XQD_S4U^<V$ 
@!\OAHKH+Q_&=L(%F!\IG2IJ((TZ$+ #4_@ FY\.M?28 
@X9;G>VH'G"4:=0VY114"19CN<:HN<""SS+@O /4;8S@ 
@&'W*Q!%<I>O\@\5KK6=]"<S4Z>?/6G!C;N6G6AC5&8\ 
@IA#O2RIA36%C*A"UU,LR%DOOFH+MX,-^-C$??Z?DY9X 
@C68UE&G%0) N[=T2N80%Q[Z>#FO/]"!E^9@@RG^L^W4 
@>QO[JF$YB5R^XG"Z&WG"X%D.N4J:%%K)GL$]6,UZUPL 
@.6$1N>YG9 RB=OY@A[$/!QTW,ROD'HLD"PR)G*(M'1, 
@9@!RLFY/ND'1%-JCP7<&1X\PU P-%B*^;2RJN7!:044 
@7C;O^@:J.SB\HQU(!@/L_'A356L35.X>2]9-.3Q0&#, 
@2@LJJ.^_S^BL$- MEARWIL_GX#?E%8#77@"+\0G$P\@ 
@K>DBJ23A6A%C18_'\=M!D)_?E8_/DECE#V0(-7L5<3< 
@M1+J4$LIU+/+Y#'U.P;AMG!%=P3+8+X\ \,-Q\HM+IH 
@:N/!C%(9(.PH3</Q$9ILIQ-^2_)SA"&"KQJ>AUT5 MP 
@-@S$%6%VAQ4$!"]$>AZ6M:!)27M 1MQS,2^\:%"9S=L 
@..@"&K$)#TP>2D.[RZ[K#HXQWN>,!2!P1OF,97WE0R$ 
@Z!;;.W-*@I H,;9\C2[0K'!(=PWJ3FG&S9YT6DCX5:\ 
@$7=T\/2!U(KFYQ96K^P&IP('K>,U.6$_IDF%L)H<K<8 
@D?\5\TU;KB+JUTX6G[)0YS\&00JE)R3 D54GY@*:/RP 
@HN"90\]F?[. H?8.Y=(^XE1-HMA;@7@Y7U+@ *6&PJ< 
@6WD@,4VESKA$TVYE++\3&HW6*_;J-_:%56D:,!;5>YT 
@M4^1!3>:Y'6FO$RZ@!YX;( 0#/[W<4/MXE5,%WBZZ>@ 
@@FH&E<2BMXTIJTIUJ*L(!#%4^*RQ/4C=Y[[J;DQ,VUL 
@4J="&@IO=WO,Z.P%B<K,F7N,&CN-&-0Z+$O5Y]_>2ST 
@ $26F"AI1T%(ZD$$Q^/9]VB^2_>$6Z-/:$?6H1E_^L8 
@PGP\&M!F>A)N<-^G8) 6Z1".*HAW3;V,]J!V;WWKH\T 
@&J>@U=Q0%^KX2<.GY4R(AK?*BTANDWB*@3+S$?$'3U  
@@)[,]+Y##,&/M<08_.!*4!YDL>0 $)1Y1^Z/Y7FF 1D 
@)N37%7$GS8";V#:4]YO1R$IY++ES87@TA^UT=__,USL 
@\$[0URN_T;K[;QJ+E[5+PL"NX^O9&99=0+M=6:[J0)4 
@*Y^/4[%8RC+./2="X4V:;*0?>+M=N(9_= JPR)" [8L 
@'8:#.K*E7A0$%S6[8W=5I''3OIVHAK>11'0UZPJIL"X 
@V?&65G5*(Q5BX)):ZS% -ER:Q0HX(6U:NY SW;-)-64 
@/U@<RL[1-+C)C;,M/.^\+77!V(1DC9IG7U2LWT=JB"0 
@Y008-YIJ"%$LA-X1_?.?4*_ \.$99S["--NT=_NGX8L 
@@[@&HF>@35%D*+Y<L4' '^FYR&G[='X\ Z Y#S:HHUH 
@FM>.!R;F:L/$7N2#BK)#,@T69]4[RS1DWD"F2.!YIS4 
@&:<-9(U,4W\7_,.,]N*<A^7?,SBC*8$L:<SIP/CP;C< 
@B#.1FT^B" B3-#TV;+W5RKL<'79;K!J!7^]F&D;^*B, 
@,S-HL/ZJ,[0#)4 [*M'4)+5)+BN^J/^^_N8TS.$XI&8 
@$@?.0AITYOV%N9)'*97$1#VK4'-@<W]@O*=X(\'.FBT 
@+MOF)(.EQA'"]1P$M Y(XNUFTV=8SZI$%KKO="E+0), 
@ELX.NH$-DBW,<#2IS;'ERYY_\21EXZ1,BS-G/^<&K6< 
@)RDO*][+XMP0D5Z-V=J=,#3=EKI<5Z0AL+_D820)\WH 
@;!=%4F9S@ :;YSR*,P>Y$ 8;,Z:CQ+POM$GK_.X)CZ, 
@-TA?6NV*M_V>AS^"<9!GF4;L8FFVPZIU;45[PIXQI08 
@#IM&F!6I2?&0RCDXKPQ?U4V [N]BJ_"2XN$UZNYHD8( 
@/\F4F/ENN$DT2IZ%U'HL*"PDKL$#J?PRS\G[>LE<><H 
@:Z5S/WBY]?#BS]A4VUN)_G=3*9Z_.LIU4CXJRV?/M^\ 
@?MFNVM"0U$YZ*H5R;KH\9B9R]&X [@/(&0RD<!S1KOD 
@U:]'C C]B7V&7UU1-=: "\?*Y\&')]9>AJS(0]#@J,P 
@TVOFJ-:\2/_;?,IH@-/<'8*S&E-97 <NUG_6)SA5XA( 
@\EV<!-R9];,Z!U!2":#UGXJ;&7L\HR<X%2-'E?EA2/\ 
@-FT@#"<]/+IPH0J2NL(H'L64A:II?M6'22%,1Q374I< 
@P"Y^7 S]R&R[&<ZF2@1IL.>TT!!>%D8ZVPY9[[PI-G8 
@#E3^['R\^)'O5URGV]:>1M&M++NEY/3,_7]<M0]-0D  
@2$2 9BT?BHGO5V(HT0TAY15V93L)UWJFW+PL3<.-,!T 
@,C'(V9;II[V:+PBT?*>G,TG[Y(4^'KAHS[^YO#A\G,, 
@7WW&L:ZO]AS]717BJ^2A17<E%:'8FST'WJW$.TDQK/< 
@<JB\H2<)2BV.&,WGG1\WKHZ^Y]UWE;D8H8L<L)()?G, 
@L&?$(4XY%7IR>-RX?BKP9;2&$0S(].K5?,O.L0TG>PT 
@D91EH'VHV CYC<SF<"GE"' 3"S'5^);.Q91!0/U0\\P 
@;)&A+GDJBN<K[().T>RF'QA5_^V:@%<P=3 #,4QEX), 
@'U!M(JSB,'M(O 16BWGKK9X *E;Z2NKBX/V;/@52#,L 
@#M9-T7>]LS2%14[L6#E[=-=+!9WO[:+95JOZE^Y?"?0 
@%,8".M$I3^5#J2$3T #VI%^0BP?WA:.3*TV-1RJ0 C( 
@9\!"R+2_B9Y3=3";_@@VW,;FN(HBP]=9-@^"#SU^%VL 
@D(<R;QN^@00@-JP,RXB;/S\8]9)6!'T556KWLG5E0#$ 
@T[GZ/N#)<!H7++[((9P45>XB(JB:.S<,+D!!S^+*IIP 
@R0%R^M946;W(@H.,#T?INDQ$6X5@2E%ICZ!ZY^( )L$ 
@-L: VRL>HR,PFHB>)6_YH_-FM6P?N][1L4#0YV<\3&P 
@>)#XNE7E!QBR^J4'%6D>;.SIXN8-DP>E<+K%& PY3P  
@R.[,(L7AEBL+.KHC]W("A<@4[)RS&J*[Y]9"=&<_VW@ 
@-$]B(V\U8&73@V:Q*WQ-F OLYOP--0Q>[AFP V"MQ9X 
@4$Z!:(A.$WSYTSR'2.[IJ#^,>A_GN;9_<; A03#CQY< 
@R6I^+ CFRA+\<$E*8 TER-'GML2C(Q<S^735-TO%WDT 
@_+ T'$.JV@MU-D]@.85CR%KA N7<4N=E<;!<6Y6B'C( 
@!L RX#7H_T,Z8SA\86(4&[\(\.C\+9PPR93IHQ0I)D$ 
@NL[GEB/X0*#S+8(J?3FQ7?$ZY&>%44SP$M-O5D_B.&H 
@$\+V#L#=BY</BKIJ1@Z^A LE:'?G>M8Z@54AG-I53YL 
@%-G!:*E^[-DNX(*\>S(WDVB.Z+3/#D!9.G"6\GD!5X\ 
@@./931DSE)Q=D%7CB-I1IUO._#7/$HEI1\W0T[32/TX 
@)$6+VQ/4)H1@$WK+05>F\MZ;Y5;2HA=75FN7\6#8>&< 
@;831=_W-ZU9U^NXE!^^WQ9F7H!Y, ?00N)A?,#(UH9T 
@"S-DK8_0=CF<4KBY?IZ,62 6R:YY54TO#U8"].LV/:< 
@O!?+Z'M-WY_UQ7*8QP(0HY\4SU3T0B?R<&B"=<;QT#( 
@,-%"D%M,1E';#^+P<>UP*;DXC'=X/:1% HG*)M-6VP( 
@3H+Z)?5IJAX">!1L, ].=B_-P->W.DG[2/(7Z_<R6LX 
@FR<JVY6K+ ^;[[0)?BV?*]CL;W'#=]2@CS!<%IBB[.$ 
@6.*:XB,.O[&\N'@^1\X1 8#SZ^J(=?I.R&E6G_UP@)< 
@9O@S*&W ]Y[.*L\38"S,B2&&;_%2C%9^^^J;?CSS!CT 
@1<))?V?DI67.BJ-W_U6)%3/*$<2.P&MJCOR .BY3)NX 
@?98HPH^;NGM\6CXQ'$#IL^@4,I)ET*C@NU?6!=KHZ-, 
@3>_(IQ-5W9)-_5;C:I12LZU'DU-(\F?% '%KL)7$"<P 
@2@B!DP[JOHR!;KM^4[Q/(TFTP6KW!3F###T*CC4>^OX 
@N[ 8+B;Y-$V9HDC.4ISAB9/P/S7+H/\ )"'!HFQ7/G4 
@N;P.]3X_MC<;6A?M@%Z;1C!9<Z2\Y+?'R?8>+B+L_&8 
@3U6\)V;E%@NP6F_.-@LRK'[))2<,YC7&2Z )":EK7Z  
@U^F2;)!?CYUEZSO)WFS00I_&<83<QC5UN*V^6SGBJ'T 
@!M*[,ZNQ ,*X<_009(O;/ZP410V[/][[D),<PZ?.Z   
@,/6*T#(?R.QQ8"GG9K2!Q6K=4LN:3M@S)^VLNF$;27@ 
@F;$F/%+**$'!=]Q>[0 +U.PGKFVL%])D6$$S!EY85B@ 
@[''4E<J&= ^AF7_6*NT21__1QV_<Q4!RM"5T;]B:W<X 
@&V$:E;45T?MQ@.U[4F--"-$W&)@9*J&0O&^X1%(@G#0 
@3";AL3.CE)0=%MVCC0QEZ'+70:CFG@YC[T:Q8L-D'D0 
@)?'%^ZF:1==7Y]_*7_3Z0T#+ Y',22*C\-@XV6#@GK, 
@<D;0,WM6-<6<(+R9#.L.R.8F*O8H"Z.B NR'Y9R/Y:  
@MY[*89T0 9?N3.S22GN91L9L/#4><\3/W_HP,-$.YL  
@=%]0V7N5G<"D'KD*&ENN%P<J1MP$,*#)H9,]JS;(NBD 
@791;V7^+))L;NES9H3+ ,0H;ZG:?*,>:7-2&9+'0TAL 
@3KZYXQ&P&O[.,>HM77X\D/YLY2B"]CD4:.T@V+E5 +D 
@P/L8JP,6_BM^O>UKV""5GRMW,YP40)8UICMN#8& =LD 
@E9=D@D8201QZT'Q6-:'G ^)NT;#TY.TE.![23!2D /( 
@B?.Q(R_&RI]CKV?@4\HW3%^ I]E.4--E2\7L=+5A48T 
@R=M?_-&S)\@&-X_L*-^*O Y,=PX"EZV.F>\3_P;Z7KT 
@1O(C0)7)+7 4$!IW?'4&6(J'RTF IVW5LV%/ ^JLT5D 
@> 4NO^(1I_3S/$AFUR#1I%J(B2&-_7A4^KT X8195A$ 
@ 7X+%#<I^."KT2?D-*/]:VXFRP7&"+!E-W.%!^\X1*L 
@<H&EF)/[F,[S4-K(U[90H'5+#!J.FS79:%F[:8.\^TD 
@US;V$?&Y(/39)D11V),UQZF0)69CK#\M M(&-3,!S(  
@+A!.7:]\*P_'4LD@5ZO0[SY9-^'WKW+8%75"+WTJZ*D 
@P==GZAQ[F[F^>9ZJK0=$X%85&F7(NQ]YOV:[P#0NH&  
@-EOKK:EX;@#)P,%?6/%IX=)L_?P"%2,7;S_UC%XOBN4 
@OGB&ZF:F29^VB?;SNE ,]-2YC6-LUK$3;M"1;8H?!N8 
@>Z2@:-E)%X[?I<4\>-YECFKS-%LY_>V=<0SV97J+KK0 
@RW<KNGZRA(^\8UZ->CNB;K6_IS'$W V2(G\I_24HHJ  
@FG07\B8I/I'F\H?3US -AG=&5FDD[IRQY]N?X0;\R)H 
@\NAI9)1&I&5O5@X>^2_%="^YNRM*KE;TT-''C-PK'BT 
@G>B1^"-T?>_EL<%Q?9)EA7[*QI^!U)F@7PW=#N753K( 
@8XP-L.)<,4G3;F&()4N%_Z5/I_E%)["#%>"'J%>]Q7$ 
@6!>3I"(;?X1W&?O<7?,G)/A+7=)-7LP#J7G7/Z.W)SL 
@96QRZ\;<XB.++!_LE91\>4WB :?6G&WSA'Z^\4+\Q?< 
@9%BWF8IE.@%R &G5GH_QYJNRH,H=;DKP6?'WD\TA;H\ 
@5MK" 8)$Y.W\]DW$ 0UGNV,1ML#:AYJ$(-EUVDK,?&\ 
@$[<KNT=SX19\@81\_63,7$"DMO6[N(&X!"V7Q?NLX[T 
@2[*EYW%(2/LCN.?9U_1I'="TM7MLY'#[*XZX6B6+R9( 
@,3,H,G+&]D*09>K"QU%:-_R]RIL/YP-H>R1-%^/DZ'8 
@_ 2(BH&TZ72F;R=E]O<E/Y-EO]%E=3L ^"G)6%-PF+D 
@:Z$V/]*(AU.I35,;V0]*T:PU9>4,F]L[)U:&)V+V]+D 
@'O\4\A.88T68H\"J&^,=F-O4O#/< I>1_?B.;Z//YD@ 
@!K^VD)RO.;U2^^WSND;CQ7J/(2N+ 5MA1K&8_W CO0D 
@,S&';$"FO3;4L/JQ2:*U-TEK\ \S)98#W63?TK'BRL@ 
@FH+$6>,?U J/UGDDW>B],G"[ZR1U(JR3[CO;<T5%P'4 
@'<+6$I7=1.01=["YD#L9+CA^C0BCY\"[X(\)MY\6=2$ 
@;-E<>$)0AZSVW>V8L<H^&K,&J?)0R_P) N9L'/RJ%T\ 
@,8[M%L10<.-D6E.6&)FY9*)7Q]$:_<&$/@@Z!^'^LKT 
@4OS!'9__)89B I2(^\4.7VW2(^4Q84>T"48,;,C7<5@ 
@$]9[,9I)ABYEC%B[<USHY""E04<=6*M@_1FZT@8O5&0 
@^DMX3V(YER8FDBKICW"MF=_K5?/8PJO[]9'S,+:77GH 
@Z.^S)?MSG,).C>9S*-O9G-.LB!T^-EU@9@N"WY&R[T( 
@*;-ZM[*:X! "'IJF\[2\"#S,YBO2ZT\U@OWD&Z- XO$ 
@X_0N;GZ(KT-_'\S/=KGJ$N/$E.B^R].,O+3,3[0D#XX 
@E8V7Z6:I92HZ-6[5P<6@<&Z]X'8O>.V =$LJ(8<XJRD 
@-^0S%Z..[8+US_R\D^"8MLJ2\^<:0_-9U_8>NH)T]RD 
@K=47A*=C,L(<%-3A@KK21U0Z?2E/LN'N?!PM;E4+(%\ 
@8"_4ATFUAQ+PJ.\/-;.G@,FF#%54 $M<Y32J>27!<PL 
@8UB3]/#KZ\!0705I3\ 7I9D,+(W1AZ&2IC$":GV#CFH 
@SBUG%Y':LF.6^$[S>(3<NU#$?V*W0]#:8&B$"^!2<OP 
@DH^H:)4E[)-G'2=#M]*&9!09_6M_L[GYA/T7(3:I[(X 
@5\0!4?-((D^THPCYSEZS&XQ$IWY);6O9U3F<5.:D>&@ 
@?";KY^]?L=3@EH#SRMT7G&# F3"**.]5C_1HL/@J<RX 
@R=2([H_W4W+\DF:."5XF7Y^7&^0);E/-*?I5\9&59G@ 
@H_Q"_5*TT#+N0A.OF$Z)AK9E/<XE_S<?O- AKIOUJ]4 
@/E_FG9'(FXK9&7K0E@W&42O3;!0!:YOJ.7,:;?>0*28 
@&T)TRXVOH!)"4:OQM?':<9F/W-J'"H'"!'5(/;"-+&@ 
@<R#YF^)04Q>A]&O5)]A5>\4L^%Q9<3='2M^[S%E[<&@ 
@N@SE4: N@GG!>+V,GU$#BPF=,3[T]HTC5I/ZN274.)L 
@,^N18L*7#V(DW!T;_=E-BF*_\-?C/\^P6,#_W05S:[\ 
@_EA5UE091Y]7K;='/#I)/BR8=&9_8%N,L]P2B@H@^LL 
@ [M$XPS[R/]FU-KVAM/!]0(WT[S;&SA\S?L4X!]+594 
@(J@[,DV6Y@@7N[WIC"[2YM$#\&^"E=__<.W>$CDKNAP 
@M(=#Z$QO<W.MYHO^@5A%*'8[=JQ0'5<6FC:<[F@6GFL 
@J6K-O<W1K69#DJ>J1MG6W>VN0TM/;RW\OS<4R:4,H]H 
@PZ#R@I/CI63=!QV6." 71I%18@6=D=OL6+S)* G-]/P 
@8=T1- #U9DG"=!+.6:\H"6(189X_G.VOF9'TQ15M!.@ 
@Z5N?%B&UT2E5-' =-)T>SX&"+P1EE;)I(?0(>/V)GVP 
@;,SN+-;;A>@+!7/AIXRM/##HY?COIA1W#.8D.J&:_QT 
@^),HD>.03KJ&*@F6;AO:>EOTZ]:G"@&Z3;'@=@M,F9< 
@. ?$TPSU2_MX1>F:S=3&K[6SKCVY<26CCWGDH7NHQ"P 
@\U *X--!!#EUX8T@38O]J84$,BWMRZ@.D"QUK90AI9< 
@,^[RGC\AJA['E2#)8BT(7X;><Q3A*)-EF\XT\)==#0< 
@M7AB@";K&G &RR[ ZK<E%#"+=GQ_0'0T+B^ITMB&\/$ 
@&BG12;NO8?F0$.WS_VDJ#N\^R*IO?0AD4L'#C6-7Q1< 
@ZQQ\)P/1+#&U?@ND_6U.A/#;?9?\H^XF*<>$WR5DMNX 
@19SRJD8O-["E4H #H&;!&"62@^]))C_/$ZST\8N#/^@ 
@V,SS^N;G'.2+\*J,-JFDDH/6_LJB9<S;\8$ .$BD!/0 
@/E"*0@14[<)%LA'1*\3)1HY'W^V?3<;Y 1/D]H&FPAP 
@,+)*;<XXLG%68E2DD>UI%L]6D=GR6* Y"49CW-@S :L 
@X,)M5,>F02:??;"W_6.Z*HX%C43PB:$POBL1,!#.;D\ 
@B\)\LM-%R<ZX]BQ#A?*0],);!&!.,9>_473^R["6MFL 
@M>E\2Y[.&-MO_=<9G@$%"I#K2UFA[:.1_E4,7H\CTU< 
@15-_2U1HWMW]E:JA?(VO>:GB'T]:GEFO)>Q !(]/>3$ 
@/81QI/?7D-!!CVD,6#L+G,_B7F(F/XTLO/VA2Y?&,A0 
@]++((34YC0S]C)EO(TK)&^',1L(W78;%;,RXU=^4J]  
@16X\-2>^>A29MQP,S.:I#T[&,["\Q9;>$:W]'D6EF3@ 
@P2?&ZF0=>D@7 RNL]N-I3RF5C@%7\K\IFVF"1GOS#1L 
@WKE7QM(.N8-\CK?^?NEC*5153R9O-/.A2*NE/./L%P@ 
@JQ!S;*FIQ ^;]/;0*);34W<R8\1>S^AD@I"<(CU%^W4 
@5M^FJ,HTNHG$/Y==[XK,,31H -94X!9!"VOE>&?6<ZL 
@;Z&>7#\T8Z0:6I#46<($T\AK "UR) SJ[@<(G^E,/:X 
@4&@/?,^0HF$F> K'(T.N5>X9*W^O)B8W#<-C_HM@!7< 
@!@7SLJ]"<'Z<TAFC&T\@<;@+8L?\_A18LF/*9>ZB558 
@^;'>W\D]/HPSC/]>ZKFCS]Y!]YBQY@?KQQ3PY\:-L[< 
@4R 3(!8&:8011A"Z?/,W",G!:TBX'-7+.1WG?>)N<P$ 
@NETM8QK;8GOGROTSFB&FKRCZ3X#T+;PD/&D2QLQ,ND$ 
@B8Y!VH=@T&D, M9Y8:Q<A+T>:97ZPH/H:\ 84P"KBV( 
@F?TE %PN+\$6 ?(E!^L9J#5!KPJ=B%8(DC)XW?0P-#$ 
@]WR;C8+SJ\^1U;9()8B,X9&69HFJKTYMW%T6B!-@!:0 
@8RCSV4'YUO2=":+/S*<'76G$MWL51>S5L)235"+K'9( 
@)(#-LGL/&"*M)308$0ME&V/899@?HIS3@A%RT@ DUYD 
@>D43Y&-[(?Y9>8#VO0HYLV;UC9W-ZA^WNU?'=4&*J.4 
@\[UB\;[B-D"Q.7 ;$>DC[Z-G P]0>]&U6!0D%1E(T(< 
@$Q/O[W:P5E&Y:Q3W]9V&\@$N^8E][%K^?.&%R=B7E,4 
@5<8X2&D;D'/58N/XAP2W&">@P@ P?E@L-'/#R8)Y#K8 
@D2$(DOI2))UP,?UD+(*I6"16EL$=>@R\O:# 0T5V58D 
@8*AOWPS-Q\F)OW(HKQXX//(-BMS0@^G=!]QEYP(O#UH 
@5+ O6?N.6@_.6C7F29S_'6VCJF!M2JPB;81$V"0 U@, 
@]J+:!E$ Z[WE"I$%R/" E$K7H.MUZ>PHA*]^Q#EH5P@ 
@*G=Q.JC7L3ZE2$\34V,YS_[G<<^,.-3@K**U5?SC _H 
@-(0H3BK 242D[Z\:CHS(:EATH-Q_*VVT)?7HJEZ72.4 
@^^,]639\SY'=S^^^9 5#O@ZA$@4YM@V5MN3XU$FO/<H 
@%=G0.VO3T"'B+MM=HS.>66F4854WQB,YR SN?6+UBJT 
@O[C*PW AOX67RQ)A[G,,5=%A[$*M08$_YC18(I,OQ-  
@ Q7J<E_VS[1M&VMWWT>0L<W3W9.F.Y"XYT[4P"\L>]< 
@G-)* Q;\ZV3"E-5EU4Z<./.J;GI<+F\J9@%7X/5@9(H 
@FDB_)RDA_>#@8$^\P9%2&F8J[GB>:%OZV ;+\SK27Q$ 
@;O;M .<0C26G?_F7GRW[R"C_4N#@\XOA=Y4+AV%\O>  
@4FTA?JCZ3]F=^P*?@DH/KNH^@XK\Y@NSY9;?IW6!'(H 
@GE!+8&#MH730(PBQV>%(/(KW*RTL543>0.?*]$P$JUL 
@E7M, ,A8X;=FK?),!VE']0^^GQKZ(N$NW@!8VAIY-FH 
@PYO<]-GD?E^->NSV5Y0L5F_7 WU\1WZKF*0HK]=K@.@ 
@S9 H6!=(=R?:>$3S#7Y,Q #*VLWG+YI\F!?N_J5&8]  
@==XJ$&*196KC,A*9K80P NW-NRNAQ/=&NB:<:[</\5P 
@/3X[[/@J5Z,&GGW9A@](<VX<5@D4_I4,OFM?6?NVNED 
@&S]0)S9C6D9 !%8] ?&*(]?Z\)+4K:LA;-;<(9+H#PT 
@GX$/;(N3M;MVC>A";")EZ<E)DRNVMG)<Q$[V=OSB+#L 
@H5(9W>VNZ$EHEM0;9L7Q*^<*G-O.RQ-E7K!O,V<Q8.< 
@3+W>2DQ 2;#VB%KI]C#5JK2Q*5+OUL6W\6[&A2M!R+0 
@._O%LLJ3=#:%1?0_S01$H828M;M/MPDQGFQZLBO4AX, 
@QZ# -B!89QFSBHR,:V#'P8OD_<#E)$0P/#];\4%8OL, 
@B^3T@9X".<<+DD>'%IA'0NTD5)4NC=SQ-:!SPVU [#$ 
@T@'B\Z^0[LVI!Q_TYDEZ@W$@[JG4$T"U^0%,XD0AFYD 
@.AW4V>JZ44U @F=LSX'P,928*&P%5XR[@"-TXN1C0!P 
@A3^)?(4M+MMT,:9FBB"FZCV1/8SH?R4K!D(QV9Z?#<T 
@^[C G;AKBW_^-?8!S\T*4\=@.PNUJ<+O.%U^HG75&#( 
@9SK>@P9M7W$<#3MKBM&]I7Q-5:Z8&^S\=E[;<M<S7TX 
@;QALR?"C4G3)#A70Y7KH2C=U;R4*@4)C/HEN(3*FDZD 
@"-)'OM(X\%"\>Y@&;-UNFNO"TV_>VJDF$X+;8PC<,SL 
@ZQ_L[UV;!H?+5_/*\:OZUZLG/V*VO?)Z P7:2:M==E$ 
@KYJCG@Y#J-WW2;L%LW@UU8P@_543=8Y7=R[%W"@$>,, 
@QI\(U. [2KDF!^7T<1C'7&2CGVQ*&AWG<L]D/6G8!4L 
@?&4VB*6VV?SDZYBFC@[*@G'%OU7%('0((E(TAWI=8/( 
@;5XF3L23&^ )"O.Z%C-!<P4]?5R!YFWE+'+"!;#Z*@@ 
@^LI4(\04# ;%2M%0[;680(':!2130A6B.78)BR*,+PX 
@R,SJNL-GPN/HD9?]#VQED2J\%_,#J7W:8D5KM1@3GZP 
@N9TJ;71LQJ]$#&\)JT8]9E+]E)6":I *"M/7&L#'N[4 
@9\43GT_ZJ@#2H/Q("@-G/7K,=S1.,=!JK?5D63LPLA4 
@HE6G\1'QZG3)JGU0Y7'AHTCV[O+R#(?G>F>Y7I2 _R  
@H8X@UV6NE7AHR'<-CF8#@?"^O]QS+VOW$N8F2]HP!#L 
@M\]&YP)JQ WO?@I^+B8HM/?,),%,@F[VAJS09@+@3@X 
@>DXBU/^& ]M7H^R&Q6*Q%KQCHB$$7S6,,Y9/_BT)/D( 
@Q*"UM:9'QW8BP)^,/O))E#;\"KVYL,!M0Y^[!/!SVK\ 
0%-JM)>KKC$;SZ64B)_!3JP  
`pragma protect end_protected
