// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
N0+wvSqPba2aiE1sKIrgG4ORlz7NvP4Egu7z6F7jZcEwuSrxQCThlYRLL3vXc3Cn/sUovz0e/r91
Qkd5sxguGUJEP/ySjeNB7T6chH23utRuNSYm6Pv4/sbTOY6idVyADlngXvRPU3LPPSnEvwukhB/H
pNFQS0KA9UA5FXhrqGXzY6KDP6SO3zfe1V+Qq/LbokqHSYG+d9X4qJDWI/uxmCTvqVxknxt5K5PT
6SzU/YxW4/zouT5uZA7yxKN1DEN0uF4RM1GVpcf5+MkBiV2EBRiVCXjQc3aDxZekzSqFOdYJlfKc
/ecYAj7LBiazTPu8s22Jaj+IO9vdphaFWg0MHQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16880)
pkbxSV/DU0ZcwBthJE6kLqPhgJMzhP1N+8gaMZUo32rfVakHZn3LX/F2i0mOGH9InCmMh4G+UD2U
F0cGuCEm17KkqHrRTwo9xcYamQnbDj29p2hjCfoNpug1aCwvXxsRaNheJi78HjyLAkR922Qs0wjY
e9qGpvxPiR3w5V+xXoCFLxVuD1Mly1EsNIhYQP4ZaO7uYqs0SdOXJ3rn7781vKTAPkbAtrxpn6nW
pR4oLTCJ8BIjVikS2isoI5vCKs2mrk8YkYSiy/F4e2PlZyU+2PGAUexPsUG1pJd23dGOUoFzYa63
HRok0B5BtvsCTeiqFTvs7ebBlT7zNczrAf1KuJ0xzVDTq7vNCfNblp4nsD4Fs6HqPBl6x/RNOyyI
/e+oGd8C9Y1zeuhdof05JvdM9KTVh80XhTLUmKH9DqHX0U5p+5UnvLarx+emhH1S+f8f5Hclh2/3
EQD1/B2bHgSGL2UPMmrlYffMHxpk2jeDRFurlX2WM7SOzHBuNKivprxxIlYkM3mkLZh66VePz/qF
qp17/wYIifR4fWSX5EIVFaC3QzrHPFO4eZPqLDGnf8+9krnVrPq6HC/CH8BQfoZpejONm51xlKfW
n5AqnXr6sGzj0QzUWhyGtFdCkAK9iBzQTwBQwpnvnDMTsvjG2xQBCGmWk10rXiPX/lyhEngcCvdO
cJNzSdz0G9IKkgBMVQb991VY8mX4i3oiDhFw0LOGjKprXVTLyqsaDwoFMmO15ihdpcMGv5U8id7/
ZE2kLCspO8D6ZWdPYLHmhcuA4MzsSY6Ynd1K2JY2WCNY6Zsjy3sMYAmcviKAXaf6BcSF9ZXI7/cd
noib5nCp25z3ohC8JnnS2jSNCxKMNhKqTpoR0wi0Il/5dTN0P56Y8DhUIFZcWtQaBcdyTo8iSC9y
WOPr2m84eUF5Iv3syrQes5XrdIJQlyyhWRja/Qlci0acJ1ZCmPWSppkxrb+L6TDBPO268Ki508lT
ieU5QH0gR9AYXLMAGom5vrqUozUje+351wME1RhLhCX+69gQjQM31BA7kN6YftCM35CmvdNqSvGv
3vZKMqXJcKJ6EYMBmB3Iq1pWt5bjK4xKUxQKLacSb7ZO9o2gfM4qneSvz9YSry9lcoJ4TsvO8Pnl
EAGkWSVvWcvd1qkTLG/IoVltvb7L3RkXtnLQeZ6Pd1O+Bx1ZIa2X7qG5AC9nGAvYgaTR7PXKz/5q
2ot+LaQ2yShhuEC+yrx7VOeWALQKtbCQRiYcG8TJlJ2mNrzGGZFUHU9Ci9r7y5/qEyNq7+lP7AVN
K5SwpGYPTF+UO74IPn1WE+9L1P0vYyZJe+SKcD+fxkz1T7KLy2qrZOPXhF4xqYz/C3l1gCdC5vWX
SZM4CfCUOlRs5Zp69BfFEVZYX7ka2yW184xS5EObk4oXD2xxv1Z1FKC1WNiBtOIau7KzMPbuxKeK
LEbRI1sLDhqQcwBlE/XFUrYqoG45uXdNAvm4/PUhtU6HwNY/ocE5Bc843Rsdt2SAapVSsaOwMYoV
0/pSSx9xGn330qdoegGivdkr2LgOONOj2kBH6kSyhrNomR9e223uNrVolNXR+5iC4f0W6suhvM9X
ynsHSUPIrPxKxIm9zdtc8P3qRNFmPZnuHIYMsgz4hktbgRZ1/pOlsJKxCdcu1H0EznMHsulLFPQ7
RhBFIHBIjxGC9cYIZ/MBv0jErdUPH/nkcQa47zk/QdaLb7vPk9yt/dtVF1V3DLh2qVhw4wc+r7Q5
sAyT0fgqKQ3odC/yENGsAtQEjh78Xuqdsm7s2VY1xQgDSYsttUIp5aE3wR3FWHfbE8AtDTSeBEMD
/8hMrUzz4e9n6sPp+8BqV8bTqpQYc365mL9S3ljv4Lj7/uIR/1gtLz6/mLjFPb43F5rxFWQHepR2
LvoFQbp4l+FOGRR735eSUCW2QU3RAXLGsRLA+WzC7NXg48ZpSz2reJyD0p1hHAMeG+v/z2EYXH8G
SQaH6z8hh+9a3osl+uRtt5QwNJrf+jQeZs/8ht4rGET7Yke+W7Ymj6pDBW9uN8hrT68NCgVtAFGs
G+1yOvQGV/l+xbUuuwJKwzYo8HTqDDGhJZ+oDMi/twUda1tBMUvVO8AskiFC5a7Bd0HLk26AvrA+
TYeuGV5fEe7RyDpbqcma9If5hGnZWc9BscnF3jDh2ZoleyWPCKI1NikyVklsDZSNEoxhFdxpxuc8
L1CWemKrNABKIbl55m5aoeQ0AFEDfC9kvdAGx6W4oqTT3FwFYzlSYSMiZ0FZcLa4pUcNb/t+AsXj
6/Gj7OjOMW3mcIn/NZ6eO6sdoN4kVMtfMe1bRlK5vdlyMLceAvA6i8S0Dd0aLM5d8kMOSv2J7q76
1eM5uKgOJBNKcmSYyu2NHfcFhmUjWbryg4yNkXIxmTkFHqS13KB+3PUSDhB/s7EQuiE2MFqYwRZC
3J19wQ6wnkcpVA5MrVNgWOiCIzfi1fVX5XwukV2sQZe333EITUKK1NhhAVTaUCov4n00pu7DhRle
VO5/7Ak1Dg8Gl4rjR2GIJMUTVGrHhC4ur0b9lbYZOsXZXglKb/aHe8H3WzWVs6qNq2Gw25ltn9ax
ZYwm2ED9Sk06DIV8OKPINPXUvphrxtsoxEfH7+Xp1J57gX8GJHFnMREVN4sgeXeFOsbU6wFVxO7f
U8sAYPACLx1lr7rkKtqLBiTki2wpf+e7oc3dcam7yn39L3B8mSvpaN9E2g1swIrHAEIBQZmDLP3s
jtqjrs9oAt+gQMFs4ScVJmlvBU68VatUeSDuWgxlUDgEGAh5ZEntOJu4DOe80p1P/06jr+YIT67k
kndCAExyvS5kcT8B/Pdwwvudm1KhFGtvS1XZWfl3gzBw+CA0yitOcQ5TbjIT9NkfEWIZ29Ljlwjx
yGgjWA3SQ2QpZAc8fCL7sChXsCCUzBQaW4GHvWDNoKjQqKV+UMATjfjcZV+GxpczgD7fXRN1bMRx
Uwm6zmXQXtXJMQFCYD0qzu8itiPDDuSDwCHw4siHgmfaDyophiP+axOXhMKnI9XlJaO1X5YgQfSa
PjYqSrU/10jRRntZYi2j+4VsTxucmOcrQn9o/pIW4B49gqTa+qhbllVMrSw51dzXumQzk4MIRIAq
EXjH4hAmZWa9WPW7Ui3AyhJ1DMVD2CYS811UXHqDl1ambmF6qpxct9A7BkUnbcYhzEJxSFRJR3rP
PRY6R4Q0P5BCIjMJFeVSWYQQzXgbEw/SXig8aafKJyJpLOiuRHmcHeYDrlq7A+aio/Eqh+QBSRCj
kEs6nQsrtgu/DESuLcMGBH7uQ5y5jjJGZCfbpmEcVNvZgvaF4BgtwVH9UdP8RTrSYCukqmw791UN
mwomsuZjJRYfKTGVqC6ud/T4Da6Fw5I/7QpBkSC94t5kDgJdUn5MORAm6a9kIfkcBDN063HLUOFX
FZUjgtqZHX0GRr/9DWUuZtnBININ3r4F4MZjk62ixp23JxkMaUDzjWtFxWAeO5F5mJR8dhLembAL
8DDNT0sBQwIJF3Qh71oEq02old8/AaOUV5oRxrJbkz9XqUvwnLH8GEAJIgVoknrX1/R4BSQGJKeS
54knEcpHIzLPWGd9EPCsKN8NJ32fOogXW6Pv0G50ShqUzmd2Lfwn5WDgkMcMT+sAgoTDhNaP67Lq
0sfnnFx1Lsi2S1PcooOwppAdwtj/E3XlCuG9GB7e2pQHoDineAFgmWL7O46cEpUpOI1+k32rschj
ZIlsIa2/UKI9HPBpXQ/Xdy5BtRMvBobvCp33ZBqbzIDeSQR//PdYGMb2knJh3PDEqgUi9y4jfiN/
KUplnJjsPPT80BlmKrTCHs6OeLldl9typMNnY608MsTx8pPUgGhCfUR4+ZGf2w8kmfaJOthdgU2J
bk3W1ubOT1bBeP78wzn0C6eib+s8f7yZxhmvrQPUSaFz+2elRVW5QwEl0SP3RfUsyN4f+FqIXpJ+
Hg+By+DSwuLV3jvaYzi47F03i2JyO4+a0zWD0FRkgzQLMjI9THke3e93QgPJx1vexasDOTMCfN+k
X11V9gqi7Hs0UwOgSa8ZLnKaaRThAJRezqwbAtwXc4JP/mBR3u7wgyCeoQdbaT6Tl+BF4dZfK4Tq
3VGeSSyCrJxb1E++uFTalrTst3ahQbzSYXj0fb0/PNTk53qfvyp+VBMpkv9l3C0OaakqJFkmBBFR
mP0mlNdtZEdpElfskxuRZ0Bksifm1nP66BykRpZzfCVg/1ZSfw20AAZN/Fg9ytIjeLBqTWAGVN0T
y88lTHhMGebkuayC81kUC0TPTccGDiOUMUJ9tK7mij5AJtzfF1N3TzRrt+wcL++dJSEu2d2n4h/I
ig4cOCVZUnocr0A9e7hRVQNNqpCmKofaZuUWaMZm2r82OdQsfGzObvKywaW4GDkEJBX9LJ6ccBDM
j8gwfBJRtfNFr1eiKD7hhQ/he1ULuoNS5fslDLUcGURr/FeRhaHE+csEGc60OEXb0K7DMFSslau5
LcP/Adfsj8WZY9EW3pPZE5FRJxsU4KVIJR9Palrcr9YO8Ah08kZ/U4Ruw8It8HRm4oGv8uVuxJtm
0Qj2PpY5S7xPQpjuLbwSFS8kC7tEuOjtxzxe0GlIa1Evf1t8E8UF2WDeDzOHl71o2boHdQejALyt
18oCV5HyLNuzfrXy69u5AgUKRZKUeY6Ey3Q1QN+b9tuvML2CJ8q1BTXLWMFpf8oSatz/E1qsr2bd
FOvOmqwKLeagEBsriCGzEKD7DAJQ1Xm+NRhKKBrqFhC3H6YFAF1ZEc8be5sD/vWJUbI/fL8sj+oM
IWGPnZ15wyZrPaj/9JWQ4dZXUGFQOl1DbSpHraKutUyn24j3Waxuln1aWe92zbHHj9wPWcc62KNW
XzWvXXxYOLaeOafcaMohwNanI6kxsoYo3ZWWX7/qUEZOog5hQdnfqFqQxvYNpU2064/z3IZNWV+B
t5sA59IJQ7Ndv4cBemuUz/b/0HMTWxX9JJkr0Ca6zJOY1OMKCARep2UPTtctbVxfd6GV98Y4/TBU
11Rv1MN5KpQFJ38lLsCaAVV2NIiL3PHhU1PlUDJNgqIJP9ABMzI19lH2Lak6YidjEVb/BJUamn0y
p6DsX/vtVZNsx/BwwtDUWP2pTu3IC5pPEcJHKfWdt+RQkn+NpHU+F4SXyk587blizTgB+NK6o4Nh
R4fK48hj1h6SL2AuGlD35PuVgSMA7s2eZC8OQdVs8XrMMC0Ei4oFmWwJua6lryqIyhdVuQFDRMuj
+vlqo/b9DFcsq+4gYkH/enKX4efsCMTqVuecbQxxdUhhMFuK87YGCF55MTIlVRlzUk3/T05lAr7j
JlnuGf/ce3c08A0uvzzVu5E90iwl8rCN29TpZGDylWLLvkwqoODKgDDnSahlAcLAsv4aKgPURpzo
xVK+dqQzFf1rl0kAcZ8i9oP0zpOzgG967PRST6BIO+966Y73GGfzph86ptj2uME0+m3tHMfs84jd
QHPmCkYOTHnmPLukEXWnDyq+4LtUAG9Ukf20uIvi1OhOo1NfiEvuUsnc062OZ1eqN0xmHm6834mn
cer3TMNpCiy5/1Zpme6DWczydOM4PVCxEqR/SlW4vgMhWxJip1Ed4OJzRbQPIRYeHVIFBJ8AM+tY
CjIuW9bEGho9aT3FgZtWksGfPJvFcAYyGJLFCQnV4kYoYzWS/21Q8OjbcPuKwtatsKzRnmpyifra
VSqG6y8ozvRh0SEU90u4BZ4KYuhAWqBLE0+qVniHt0uZnsUe7xSlGbzFkjCjLER3C3G7ngqfejo4
ZsvH1tU16lk9ruMBv3Sq06ngByTjUxZ6rQI6WY4Np7llWw1HHxZsh9ZiEeqRodSpNnsYGDGA284e
OqtGoIFfWy4M3TAL4Ow6E3ltg639nmBFq7ZXGgGHVAceAxrlXy/rhud5d7OCiRyLeYeEhpRB2eSZ
lDtA9pPahqrQLPM2InIZf2f95My3gx/ZESj2DqH0K3kanyLol6QTZmWy+MduD+exBxcRC57dMEd6
Qh1wV4pbSUaplxbr7DMkn9mSCE3wQNvzJu4GQBfvxALk/Sg++OezG/6OJyNkESVFlqMrqyXHJ6Fm
32zqS21YCQFURDnf9De8MVI+d7eqLxk2ApCU5jm+G+ca2YeDBytAvV3VPPDH9V2L63Qq7sUxKj6W
Bh6l6bUkXbmkhpvyxGUiPaMEu0n20dVDj+JR2ius2xsD+mFC21tiffTJQU+0iqDzTKeYVOpRGsZu
d7xh53wZFB1T6Ow6A0PYozfWXoTwdqlqYTq6Wi1/yVatXh6IU4QnbygganO2jgasB7xx9qw1sb3q
WPKRR5AR86xQJijThtZcZLEOd/sbe5w+FgP05X+sPm56XLUFNmHmITfA+GsFuEWKxdaBmJv1BjDX
+FAC0f9xEmGEwUeOHouViWxtVcu70makx+rLwwh07dimsGTxJEvu0sV0zvGm/2YZb/OhkqrOnbG9
5Ezx+HG9aVqPqazbfDIaGKZQ2A/R4Fnez1b8SeSPtQW1ez2El4WGgwLe3omlQEWtqKwb0C8kzGND
eyxc1qxyG/hKipbjaXCBE8OzgsoNJ6jvwiCYhrosBLMyN1NahSBaEq+Ava6ailNdCmz666nzSV4D
SqSrBJUsgw5txKzkxY56Pbwl9GMKoRyi0ya6ciEJzVoYiwaH9xk9KgeNZPRLW+bHyaYUl+AMw1z1
zwAiPgxymfyM+itK45k30sMHgJGC3sKpmOv4yol+DlobLGqvzLnKmIEfw+5++46sP01zv2Yw/bA1
nDL0zSVRjxucKa0yEvO/daiw6XRN9HsIz6+Xn+/hdlL7OcmbF9hP3/IFF6vXkreTep+bNIvytkCR
wRiZpGIp4F0WrGiYpmy1H4wu4W4AUZAePSi0/dGFj2FEEks/+7wDhFSpd5O2mkP1fEwszQwdkJ9R
b4duNBUGjog0RvmV5oQszyQeMnbWVn5iax63oKOYKIqnvpuldfQcDjp4lTqMr9P5+1CwoukY4x8D
g2uRsw4x6X34ROz5mjVi5/jb81JKBcl2lvMQ8+NaXZUVHn4B5h6kZtnMFFDE8vRkvoGmM9cYGcV9
lX/051cYf+DX1rTr3Zwkv2Vp3wc+tACs4/8Jwdx5d6SshQwKnMn/HoiflaaUKcLSijrlng+fGJGH
MSg5cTtScK054bfQnUcy4AYP0fs8lY2hQd4UNj2/1m6IHtYlCsIIPFTGw2XleBC2Q1Ri7K2zRwbz
HRdYy0+f2/yyIMEVZIAxLEQFFdMR7W/swxmTAPONmUTygzigqMpK5vzBuhJ0tzulv9Bga/W12cyl
9TBkcRzxGvlz0z2/T1B26KyeTiSzDB4jc6uaa3HFx9JoBAzFg7x4Nsj0UEzl6m9xebP56jxdoL4M
4dAq7lGLyx4vWZ23nrC5DI6uzns4cPDVf5KBZ0lRsUMYu/WhpeHhPWhc1+rn9Z2I5eRFVWP51ugH
pV3hBJydZSCoxw0UC3tDVpGYgmODZ8VQbeSKO3W3JYFkFCxn4VYaE8PK5GburEuFNjs8tnk/xcST
VRDbCOAJYb43gHPQrx7uuk9RsOKBkeA5gENBZ6PTZNdyYL4fxVF5I55uZ9Uw0wO96wIf6vRkYvUy
8mLA8brUS1Sv4+gz2MAv0Y8Oy0LePCqpt2E0fDgFG51kBE7tNdjNYgDmOK4cRHVAGGHp/YYIhy+4
uiNOR9pFCAYq3NmqGZW+kCt31MJeWmgFJnyNW2h8cG3FXj3Jqr2yLGmfko778ywr7derWB7g2wBe
nZqwL2f1F+zgMqyHBD9L5DRxcfe1fx5BFLdauuizGsfYBJuEMpLkE4HXdtNBOqt8I0w0fKE4nshB
jzQ0O4xxTWP2vc6NIpKbNnJrUVVBd7vT09b8l+kP1sTgVuX7SdE3rVi+6RnGeXlpedBpHec+nmKv
F7t9viLM07laT9qSBrIdYsn/kbaoRs9GWrqxhlmW7CY7TMfcfoGiLTF/Pf497YpUYkZFpbUUMnRo
pCBxUUPG+MnjP0S4JWgYBfiqB56dYY228A1drbyOInJ5i+uJ4RC2MOyoz31vfKGGBpcm3G3XSRLC
G9TBURa0NHlLcVSHFHmOaqOi+Hur4/kky0hGUy1lMVv4ZBvcf5LFWPY3AitpH0kxEuald6AEjLmA
q74hGmuMVkBR1w8RWWE11Fz35x22hkqbJ8TulFKj7BgbKPSiD3vmqvsl4nsB1YTHs1UQOYTjFabC
iG42axQwRCf3TZF1Mmn5FK63ZJPlizf8hMSuIQpvUCMT945sHxsocVMyuSXk4keyYnAPLlslk2+4
xgvp4aZBUn7v6ewwLhgpXBXhdvMULcPNxCcRQLo/qLtRVd4qZYl2tjJitui+4fxeyk0YHQdygJfp
i891SoruIWVbJBGr9+kGNCboTqg8YEiJ2sBidqib1Q3iCLJdbT9oAHYIv2TVswsLcT5kNoYLGeyN
nHsYrYqsCZq3K5MSAlL9O+P273WYZl9Q7soxB6A9ZYdDKuDy400TneCSikb9w5Z3fdv/BT7mvcsK
67DpcWKm3d1U/O1H9Oe7ObnA7wrGe4zcszSNS142yVPo8ChFWUBCboxDXkK2o16+4zRuUcV7Dhjl
FaW0yiwu1m8U+nMZLmZOS35ui00cz1AAgpliXLphno/OUr7lmwuMtK66jJDFL40oI1gd7c/OAZpU
0Az0iglPSRNyBdHjiuPQKqmvGR8bUUsk0/MGcDh3LUNPcaXA7DMlFf4N5OE2+lHUs42uvc4WAnA3
uSlfGPb7dsKxOwMX7Gs9B+ZfjSzA59al5IGm9KUCHMUWytfA8U5b25JijCzj4DzSVC1EVsV5FKwx
p05KLTFuziq5OJdChlcdKRJwjlC9ihwLyoZSEqdw0BbvHDQxVrxDyHedasZ2y3w1+W9OPIkR7zCt
1s8Jrz9/RszkdRPPOOenppYOvTAD6HFqFL3j99fQo/toXdfrc74X0D8MPkoVrN1NSc7t3nn/26XK
pltcNTx4LM+Q1Zkw8isMF8PLgEkIPWNw0JYK3eFmOBPrIhUSWfRfcUF7TNXhM9nznxrCcKeJM9VD
PhTXozD+l4eZD22d07jnRtPqvpBFiNI2a75doNENbKJT0yH+SplouWMSCq3idiN7iLV/V7fT6qTu
eSkL1kdwy22nqEkZM5Ypx/Jd7xbwTbNIeSedc499Y9cnHm9ib4jDbnI70Uxv9SZM60fP0jJgjoBH
u23v7m/YEKTq3BQZHarezPswjoKwylSE1hGez/GuuYdNm+AsTtuU4kKVYz/KDaQHIj9dJQouBqC3
mXs7PY4Br32DQwaJ+Mwz4Sj1eXitK0H1NHz3/k9ao4iNZ/cPPd21QVFI+iQmjZHkz5eraRDrSRKx
yDu7ZQmpOsaWvhSm47Wf1LWoEcK5NOI+nz/6OY78lWcYmvFVerRd4+XFhADOK93f09CvJcSm5Y+L
ujgHkrzH7lMaYZyIs3OeBptz7V4c2NJXfZ6nWlluCnRY1ekPKpGooZBeHAb5RWGjq08qqjvuDBUi
RyCPuQGuU5Hzskl1ovmgfsYJBdDBTZM2jOWlQ5Hml9rAS5mfMMumgqZeigRfqrPjjpbXWej6lptg
TY6E/cnn/AaxxuJF9BcyK3QGmZjqnxYTRJBTx23sJxMuhflH3e8yfkXfNn0X4VZYqp1Cn2GpGwcK
ydQsfkfku3V2xjFcFXKmaRujTIEkCePtdjG3w0ERvgct1CXPhNDSTtQ5Mz+l/FEIkFidvZK+J/u6
iOjtYFzp+2ZirVDvp+z8jXNTHK30cQBREnBtcRPA7SHdZ1/r4VJIvxHxapRBvw6ieE1sJscqLRxQ
woYmAQ0YTJCiD1CaWZVuy0cO4WulpYorCR7CJHP+VVjQqdJbxq2Tdp4avrWcZGYNfs4qhggy+OCh
quC9j3PUpWp3jGnbtxUvuyIsdQciArX/yPAqR9w9QDgpoe6zDYTRJ7Er7XqbeL/rbYIDDyokjcAa
19DC5Wq+a2n6zURtrUA1UYmcKt52wP3DyNnoxFXGRTDiWW2tDu6O2TzUjttlYNNewgvNlx0cFPaq
iWu6fcEbR+FCiuqzqz1J+1ICPWElvMUpY3nlRfBMnHSYs6QkWfO05gZttgL8RYgmztKifZJXNiJ7
AfgFcZmFj0VlAHei9/+bSltXiR2wqAC6gWDS0SnahNxbIrLwl3/jhAp8JGIT7Dt4lGhKWZdyjrQO
j8kNLbUfV4PyOST5RNIync1QDex8d+irPh+xJYXwbroByHaqaGOy3QOA8Ptb80lWj+tucRcU5O+q
snSQOWDvFDR5axo3bWFLveghJhbvqv+d2vPBvJRpYP7nzHoNlXnte65zuvukpLX/mFFPDDWdj/N7
QPtlRibOGND7qlvPzwiFwAe/oc7ObxkxBDZ1bR9QLhxy6PDTXFJ1imRcpvb/E4xRwHciX4/d+fCi
9+e22b6oflZ1mPwNbsFG41soEEPGPE3bZliNGjklXJPThwR2GpObVA2kTBsOBZQHU2VqdtfbOl0c
Vtd0gopsi6aY+TmmIGWNXdqSF9sr3yKGbzosJO0gavF2+pJ2gHqXqljDMzlu/wdbgjIDEfkccwSX
DLlla9oU9CBtUHjRKNBNcscFqxaRte8XcFJWu+v1eHx92qT556JXM6LeS2PGIXEXImFF4Xbw+b1h
HM7q6lgdWvKCKkxmrK5Vz4bNoRVDOfP77oMEXN7YwvXYBZL03bcpyEa3HV+I8wAJZj//sr9Wy+Cr
F5RcsKOe2WYzHUZkOHxxfERjfC7911QYRXBYPqblqoGmrVE0e3uTr3jxSme/LLqsl09SdPdGcHNU
tI00tieqchyzfvSQTz0FjjVMl4pvS0ohDzqqn8+cR+tvK0vT5JKEWxFgWIBoVXinBjP3Ud4VXT8y
fcJRlonRCqCYD8AEos6S3+tZWhllJ3/+7Q14zcBZWnQ1+0HX9JCSB3BZAYtGfNkxFFrKd4KBv2cS
sJVKLnqHYEdqYFCrKtBS/tJaywjSSppTWc00HKjD5Gl1492USgfyxz0BCFqUayB8w9ZCcEc6WDJi
VuwVJ5b09GT1cYqeCmOTSyYuM8xIDY+2Y2BSJ/LcRZSrs2D4SoBn0WQBse7nDhcPHqdfSs0wLGz6
pTzeFXiYZH3FCeOfBSEwaKO+x73fDrZlmZNcHduxeSFY3E2urfiVcgUFfxr803T6RIwd4YOPEHDk
iS6aIe2ogWNztv1Y1IRCiINAR3SxJPSHGlUww+djESJicFK5Aq3keS3kH1W4uvOob7vYck8Gk8K8
PeyKV1hpH5sijpznMoHAsM1qfuUhhvpJJq8ZhFCmUkrb+rH07AeloKQkAQ7YCv9ZSrlAZjZg1ce7
ElFa/yA9Wm4ktdKACR99MCrOwBXzTHItV/N1wbh22uqm150ZJHgTxoi6jSceEbuGYX2L3ZI1tc4u
Z5HIKKAQq5yxXr9y7EkHocmOK5N+h9ELfRhkZd0gH0LfxjEUK0znsko4Mo1yVFacvXKrXF2CHhYa
Vq+JoLq8V62DduDNA4MJ8XaBvCpa70J1FLhsDYNxfdux+Y1uXde/1oP3EnCx+mVzXB9/qQpiNc7w
PqZuxNfTkiwqxX/1WD0bNmQNsRFS9Nempq8Lrriq8c4pSeA68Qxwap6cZg7+FjUOLS0M/z7BGkwk
fidtfY2sqMh0bIDF+zisBp/J6qhLauLnFXxPkaCnxBcm+vpVeXr/BRjjPMQ1u878gQQvx/a4lpE3
c0k093VGk57CYU4fooENXdZNWLmG0Vn2V+v3pdOTYTHy62LJQ1Y0m2ylJnRBovulMD+XLScjOduh
+Yr9UnG0rRGFa41ip6JVqhtE9NAJ9guJzoFOQUWCUmXuZxZRuV+vkxxznIz3ijDTLMtwMGfDlLK2
98iqTQoDVQlFGuyF+ELLO2aWTi7wOrnw1dbqsIfBV9bdtTR3AEYi8HR5zb1dsbWT6XZbbKuRlyj6
2C6ojlzdhQ+Nh4kAGFYURP+rYleeRPyvMaJYxfQVeRxYvkWqhFP7maV6Mbr3Lhwgg3TaRqjypaaL
9Ie03b0ZUuDtEY4SGaTYGTjl3nUPpTZ7JEeNRn1T9BezEGA4zdiKZVZ1Ywst0lEhMAJ1hg2NRlo+
Xu/UgRbcBv+Bf1uG84KASCN3uJhHvOhaSHZ3rD6O79bJYaVM9COhIwvIlZ1+CyoFvyvO0gKIih6d
DkWQ/qiV7txDJOQY+p7cWND/ESL+fbII3VSfIWNySxZVJL+Ab2qNhrKEToO2WwKvPscoeWN2L4QU
XzZE5JTNw/Ko17C90Xb0uC8nbx9T7FInbNUx65QHdDmvCQpxZDYu6tfj3yb9423IW9U4Vu3Ywx5D
YUtaLfqIHQJ3/wBkzpDKxfhXhtak3Zry1Aix//nWdKH3JTb4VeOJ3xNKSfhLl007+kDp1YFz/Mmm
DR6LPsE6UdDL6ZXDmT6PTiywwCpOt0W1qKhcYCyAsDbQgnw5+ovKISA6V8t1ztcFuvDr4F2SW3/y
GGP7tvuyocNUlbfeoMzhmtcSUJeeDQLp+nqVCIdoBYIU94E0DtUKkEENjMbOD+7hqnS4Lp6SLnWS
hhDogkw0ggjIIPW7m6p3qSwozbCsiUAFvZZS+7S0DisLZjToJGI68Ki6W+6efqaLzAVQEW0wQHxG
UxL89sbY5kMecSrcOxq38PMFf4IcMTLuMgsMsQ0TCQSl2/Hj1Zd0dzPWVDtq+0j6zxPzPC8Z7HsE
9dHsRclR2AxFgRY94mi4y9DBEgWT8enRKcd4f8sIUcqsHVSOnd5N4/jYv3sXiNUzn3mt9hzGwSyD
3icSTia6IVzXarVE82O8+xcdzWhEkDtIz8twEGHyjaWtKaOCEPOxMvJMnK8WyDrIo5f6sB6gVyOD
JZdELAG5cVMPA58B+nOmDZGorBN8clRZxOqBZuZqzHV/SUpV0S7Rz/T3lBUFWp07UQRiM5kbD+38
Vffpig7OwCDhl0TAeY+5q5BCwV0NGWm+4KL52MTo0ht6FzS0QA3iPRcxa7ypgJcqZS4+Gcm/HWTt
FhLOXeWs1kXC89jVA0cz3dnT5N5Iihv/50qiWKsxINX6LlvoY7115g7uUFt+FNB0G1lswGrc/BNX
rhoes0h+fn/1DIjkLPIWEeOTmKurhGDoroYa2nocatnVIbYGEcnU+WLqZjJHQMKHfVwaC+R3xgxj
I8PPquAg1tQ/cgCwIyS4Zv63+f1HPVC4X5DZ5ntJW9XOPfMDQ3cHUFvo3Vut1wT3KqR4v9R1Dxgx
IJMxCFz7nUfuNBl5HylMmsfEHoQNrtC8SP3q+llq4fKRx74u2IdOBz21/uj4bR+Snuz6uL40eht2
7PcFplDbykd3nxT4lujxvNzaiLUyfPUTweM7mRmtRg73px/h2MIbotaOQIHwdzRtjaqcPIzh9A0X
inCUqzuNuEUyTxl8rcKUL14qdh4XU9wII9BHpaAYFoIcguNpehNzIVkUQsrEktuhxZexmJ2/+iIh
gn4VPeT8VIjrka8hzhXEZ/UljOueFU5VJ0XEAm8dMy+CPSSOZlcuPB17T7ag3qcgoh5NNKS5E703
X4zYmCmzh4o7RrkL2Myzsj/bWQhP4EiHtJGpmYFvLRnqELvQhZuDO97/SI+W50eRvdAkNjX8QyEP
4fwBAFoRvK326WQ65zhY5kajI3+97dKMNvHdwKDqINX/q1U163oMW4jdVdJ6WmqGhK8JpqIjZjd5
am/y6yEDPRzFR4G0btdcfxhLJEMS42MlZkDzUxLwRPDWzkDLMCU0tyVeR03FOHzh2NN4bU0/ZafK
wpHiHvFVO2LqVhliMNuX+W3f/hKacOyd2HSJbI+GrbnIpig5CLAlIjnQLGk3sWtagONQH7xHeCXH
BBZnL21dzwSJqgmH7cnKIGGBcyXDB5RfIBhURfhbJCfYN1VzX4nSMvIIApioFhXORvBNbpPT+8Hu
/ROktpRdTKYch1w/g1dPf47koCDYmhGD9yinGRQ/Kcez1Cc25jYRE/sA3QVa5d8xTrXHwc4qt1CZ
3KeXWZyLL8VDaJ78HMiCU0AoSrs+XUtlVWV9Ww+Ep7N2nqkJYQz6d8WFc4kZm0nKz2kLJkf0kZAL
/bBNRV1PVHVXBQ0F3nCsZZcWoF+EcNsdFREnSD0YUvc6bxFLrIm9BNwB/ULb8C6wbJXP9euzDR+0
10JURWmrCPCjp+sUCxGIlurgwCfc9g4eRMCXA1cVy6C5/RqjBEvr3K1bfMSA26yED+xqzm0OFJqw
vWJiMxeOpyZYliYqWD/kpkjoJzsvTphR9c/SMW7Ktpm0tc6TGAJaZ4KzDUmPEoVGqazm3P7awi0N
vpiT/IlNXElWBDu9C3aOswbGTS+W7OIPdxRfI8T0hOc2sc15or5IhGSFsiPpQSo+riTwSQiBC2G/
uNRpMdTaVpuuOgU0QaknIg89k1Byz4n9ncTugB0tj+tqj4wBYmMpeX9pp+eM8GvYETGlIgIwUzht
Q3sA0wJJmco4OmK2Iq23E7AZgf4eqGZwWb7dcPCYL7l/Gae2C5nx+D0iZifbCUAVqrHFH6/OAKlS
RqOAovBycz8nF752+nChOGRY3jeNGcGfa82mQ+6maG7y3SXJQhaQXrqdVRjI3OZeJ3eGE75tOdpR
NtWqeRw6M6KK5TQbv6XA1ipezP4EWu5s6VN377brcTb0vB2Ne/EDXZOYGo2I+2FqlTcmiScW2oU7
sCrvYI2mFQ2eVq7I0B9LxsuuRFZqV7SbqlfM+7auUFiXC9Rv1s2gTnn28op0vkg+unp6yGf8Uy7z
ajASWKVe9lM9dtk1qNDBYQir/aOyxBijNSx6AV8YJ4I8LOcdeX9QQMJ7c3zlpAXPWJOc04dWWZ8s
5lHVapCWti2+4ojcb1po6oYlVCg4XUOKywCIZ1ghvpAiVFYYPj370yQuwENZEh+SictZ4dedobES
KhTdxehLRfIDjnuZ4CpXAZn1acFnd/tdODryol2Irmnuj7r1tT2QlvHGLSQIeHUr8Gj6QDqLY7Py
EJyW8L/SdlkPknsjpMyqPwwe3zASHVBJP7SGbg4TBQlcflLaY237hFhULUoGiM7alqFhZ97GWRP2
hTHok5urcbWykzLj2qNdIpF9n9UxIU/YBBrX7CBxW3Ra0sb8SJStvaNdyIzzlkm7pkFDezaVMH9g
3vVR4DMuncq8O7Lw4uGvhc2YXIp6JcR6qL4+T4SKYAeHmf21d2AwbdbiLFNBJw41H8815c9y8ERn
dT7b48fZ+41nfDE2xYAvbGNDd6YqEw2b0pMZFgRh+lap0bepbBBwxYpk140+4jDVg56O57najYE6
sN0fUg29mhOPCDKDm46A13bWxd73CFe5Iw2z/OEsKFFYfBgQorDsTKN/KcDpFbigQs4oSJwAtwbw
5g/wV3Uzr3oXYT8I7cDEdxJd8/3oNJp+2Z635T34sh9OvXcIW0WjUhEYVv5d9XOjuN81KLKrHCXv
/sID4bY9fczsbArv4uFa4vN/rGq4Fqbzo4FT2Tq7M1/E3JpTFMJoyuovO3qnjrO85mrXSnkel2k5
btn4Iyb9uYPffVvyUYpD63lY+cv9zwFaDDn//kidwq3WKRP7zBo6tHrM0EX9ULXNg3XHt0hzCCfe
UrDAsXKg/WjxDtnN9PQGmaDMVoNz8yYVL3F4WBNoQyQShKtsJLecY83/yWAE5WHqXzbw/gptZBLW
Ml1mKRV0whHEhEqbmorl5sbAvCCi19xQnluHpOUGK74bLlaKmz+gDStaxeIi2NYqoB/TExZkWYre
R8zLSPMDAZtGnc83Tjfyq8gV3QY6Nxjbbf6hLsTuPu7O8EomypZ5CLzrTGmRBwc6+0dHYbVPRs8B
MV4bg3F+BShppGYeTOpEZ0VuOkrsKXaFxppSkZ5O36bC/BHNWMog6x004EvQ1qNw2da8EFdOePJ6
wD5ybd/w53YOrY70C7uBFPdl5m9JzfcPax9Rd7sgNWYUSQrGdycavcVEbghzIy3C9orsdlBe87yd
kalhl6dzgr7zXRc7Uz06jdbNalWI0zFKgqWGSiyWjMVPF9FUKOVcIVdayTweEe+1c09K7sZSe6Sj
8nMqHJQdYaX18eVulfAOA9YS6Q/z7YqufYgTpASnApiPqvP8nduCN1bpCY2UwA4i0DWEtqmRUn+U
dpBPqfAgQI4KLj+3zvfWYi+Wwt6EKSB/oNj3Jn7WYh+xfqB9mex3hZb23Z9heA+nbN0TH6ZL3sNT
tWEIXhhvpz+1xqv1xZ0aQbPJMkyrQGR7EUbHI2fI0APKhtJWVimqnlJtp7xX+MUndEEsLTBMdWIB
sjTpB73IzIa+i0lN9awASOe4PigMM7UweK0sxbgt4z7HXp1EoPPR9Tdw2t9TmiY0P+/BBUlHrkCq
2+RrUAZpU9ZEkwxWp0GR6YWRHXhpc/pfaIjOGnLb8TsiSyCq+TPKDGAtGx+3yV5NDGlTM30mBflE
7SgR6xEZObU8cfFG6Ak9ipqavJrvXhsve4IS0zIVDAXDTHkvmZ1Bxu2MfPl6sRXhiBWxG//t0pvX
9QRj83Px+5fe3QzRncSmvS8yuz4hUhAqOSR/hpUOCnH8qi74xaRy9GeINjApJs8ncCNO3LpJsEgM
dB3xQJ+PtEE35/OvC1JNlx53HwaLSzMz+ahYswvDoF6aE1ZWU4kaCDg0YNc3ZgEzNoFy605ekX9d
FNSkgreq9+njQ5qp+35rnmiyWIRN21RcXwvzvsIIh6yAIomCpGYLNLlUZ7FR0w5o131MfQThQUAo
DHJrrayGWDRhGazuFgTnyxBtctty/fA5zL8AcDFYjeB39IKSNjtYMrJQ0wZKD3YGdaZ/GtCUE3cJ
pblPV+lzLjRlpZLS3PtA/vRQd1O9G/pbm6jKWlfpm5fQFNF2V/dO/+mZ+eW4aRoZAEQz1jVg+v18
VZYqoYffJsNj1OHpvumKUsoZP5pymlA9kJRR9FzTc+e6HZkRjPy61MBzxQPW9IeuyJrgbmEp2ikG
CS+iIwapObfhorTsjGZOb4G6c0efSr49p0umWkb1cIlSnAB1T+bkEuP0YgzovM0zaS5242nK3gZo
my0trzkA69AvOKPwWkbhhjrDwKTZEnxyZ6KYw7CgQPtW703pURyZxQy65sew+bV5jZmHHbHbPJAT
I1ydNRjJVe676jtTxi6h8Mp5KzvPtQv/F3afAt3J0UnoAVgWMHdOJCN4nm2bwTwsy+by3FLOOXgr
IX2pN3lqvdLqZI4ozLcCGFvzx66x9mqQ+/3TGG+I+QGeElVhTGWgy9Xs0101zOo4KWvbUv8qwLsm
NeFHhbWgSTf/2vjcGoPdF50diicTNuiqlyySxW1UujOoFsEi8HPLAlweAr3L6eFDOk3czyReduHv
lxNEiUXwBebpWsRqUyPxwE0nO62TmzCeOi5xLK+nYIm1gQL8lT/OvFQyBLGfzFgsrdTDgR0wcoDI
dZRkM0jqBDXgcjFcDIfuWcoiyiqjoJDJL5yzFbvVhwRccyLsiGrQ2UswnnA5xJGHKOPfjTpvZxEd
pFCuZ+/QMzg0rabSD6YkNk5DGIG4o5Rrl/rm3si2kNQ3epvxHqe31OmHZwDOMXJFbxCY7IK1shOO
pmHaKDEH+9RBs+nGmledaiVqHMtyQz7gkX9QGYwH3Pghldm7qNiRyIKU1uzEoMvhjDG0727SJZy2
bm7gh5XUYuhqRtlFDcfqBjmpSwVwCwdvxBBuyNvXGPNHsihOnBOGbx1kqTPKfq0WUuk7hJIZFbJQ
Neuta7MvTbCAmw3Ig4Tz/JwZJlk6Mty3BrtG1p1/RJGiuxsmxWNNAICWK8D/U+PKzS423jLcNaZ/
Mm1HoSQfLxjj9NChxxCA4vsgzFQpTVpW3KWZ08IwPTaMMs9dp/BjvrLjGb0x0A/6ZPAl1V+gpU8/
hr7+2+5Aio1hpvg8njT0Gl8JCsTKcJoNcYqiONpN53elNyufFwCRdgFwAa15PbKC6To1XZRI9mhF
roTuOOPrwDZ5M9GE6Wpo+MOVsd9jEoVPsA/5PPy547sJLqd8YcmBA6m2D7d/NIILAUptbiMXPiK4
y/g52e5TxNKmOPqoFn1YX/chTI31uoVDGjT2/tmw8OAWzErqYJ+keiWNCLivj6DBSBd3Stkkjc6G
L9SEwH9t2S/myoY3YciFUfOj//brLu4TlhAL7+igaUitewNMosINDtwd+YHhV435o3wvPkGRB0sd
c3IiLgrrauRJufLUDa3umARESInV9DfCD7KR7QKrgAbdESRscRvRAGmolBIG5MIo0ym5Mb4H1hFd
XCaBADbVKb6RLuBcTbXOf6dXHDeT+Lt+KlW7eBEplHafLkv3z8nMQEYnX0diel9yybgFeXoQ7Qdm
PaWgRF+QCYTe31LosqtGhIbY2wDijIkpXVUhbzZYllH2hkNFe3/1u38YjypH3CoV0hwWoLeMN22/
IL+qEBBYDWjpplvbD2OdamX+zg7Fw/ESGR+J52xhmE4WROuJO0Ft9oKpTKQzQR+RDbkptb7nhMT0
Y1aJc4zz+CgchM8H3FHnYK6lvaGT4WcmMZtdpoy3noNR0JmSUI3Lpo6ghBenVu84y11jSive/c/r
QtGWYbJmudMoQ6psXFl1NEFvZFId4hWAi27FYBzWvXVhaNnnasnX80NqWNmsmj9FPTf8iFAeoIVK
H9vc8WqRaq/lxwOmz2Z7jaeM/f59Gjhu4vlpAN5HLKCCiF7fABwgIKaDqEXkjcNp7aP9uv1lmXOM
r2LQmv0TQmm1LuEMiFB386b+fRTIpr7UpIP5WG3swPvxif/CikpEA8WiDzk6PjqUEwvWqujI+LOz
e5kg4JBv+pDV5QOfnTS9AMPTiwnO9w2rTYJuz21x37AD8hsvYbZ3a2eJuwOUBHvGXbJNHs6u1xJk
U4CV0jFFcCH/7WUnOKPDPDQdnmW4e5zX5k8NCdrYUnl/NPbHUMELuJTGSeW4FurSEPMhu2fOCg/s
pngWyqAWVIAaiZfhNEeMQn+iSbcLr6wYzdvQJneLAmMSOzyFRXYb2jkV2cHnzE3zPEeH3UR/5+QG
BS+bTZW0HDezi84Yugq3+a4DHBlX/4Rwrrw4x3DyX0vrFQPQSPs3qJILXtZNYFYv2DofspNEwZfC
hgJLSq+Eh5lBF7lybr7Nz7GgCWYees6E2vHv3D+tCn2Ue067TzMX4xGuZ/NuwAxbhsfQUOCgboWw
Z3gjPTdjtPQi3ihLWEs0iUxbdgXNBfHffyFqVsN7adue5lCLrHw/6Oum1evNAsDyY9B2qtZDrbkz
wDtvKYgmG+M60PECNo3SekIpSoYLaI2cqhaUJR347InftY4pScVPmSXczRBuMjrmAku4dzG7FAFd
oynmjFOsRGwGKAWkgbNWNS9pd6RoIm9N3FZshU//PegqrqFbWmrXszX/WdK+jsKR/Q022NCeiTsL
Gy2vlPCvVECoqgbwrk4z7ur0b/Yod+uEDzCHjvAe3yn4CIG/JBxbGPb/gMIiRGnQgIvBtS8thSLP
8CEQvBb605hY+pO4tJKq5J7V7ahc+vvraKu5LSEiWKREWYpM9fMJQonE2JaPz7RddpWAxWrFG02a
riYHLrJgfWyjpxbMaI1YExib9j5i1BoWLWUl8P6N6jGafO8XaWNfujaE5y4I1uEjaT8Bl2ODPd1Y
/Qlh71Vt+fI5mB2PiIQP6JMr04LpsFRc94lHYI2fEDv9jipEXSX3p3gHVkPMqgHWBw3d0NVkGNRf
vQGzV9LfuT8M/kECLzwcOptVR6tyKf76iQAuyvx4nd7BRZSt35ikFFNj4QJX+/j3V5XsCswx7Eho
Q2JdtpwY84/OK4WrhOM15cA059ld1ilrkkVHAp40AJAbQEb0SNvDMI/eo+cMRgxzsmUypckOGuW7
dl4nYBRH3n+jXlLD5IL89fhPB00xpa+BO0oJ9n+yYAAxUZWuyozIDLj66AWceG+YDb+3E77RR+UQ
DDyoDhJAogtyLD25ymIuBcXJo5gQYc+LPbKucQOdNqjar8IWpnWXVZKKvum6qxHlnJwf7N4PYVrd
PfZIU2zLaoJBJmvQFYTbYze2cLQOv+Rk8QKdigAEZooxchoeFsBr2jOiWnWexBE/MMDchdyc2OqV
RL+RqJCTSUkwJuIbABVyHnXo/viVrDS18mShHns606sa5JaSh8pgounkOUHrmjosRtoTB0YkdrBk
Q6TP3+gXwWM0tqGxLL2AITw/D/am05Dgg6E+LQhlUMWrGKC3oa2KDk5/mXK1KYZHZMXon4T1A/sH
57SkfnIU3bJZbAf3GrJzCF5J6sHPh0GpSbuCZG+w00A2vMqIp5qdu4oV1UoP8QYxBFzmb739qKpn
OPkRzaTX5x9Hz6ndykeaF28noehC8E+P21rzHhkGVbjP68jMdNBEIUiwxibQmGGr2XAMowFVuKg7
xdocwEvS4pVx9j4igvunZjaSTx8Cdssf1ARWIBO1RJ6GLWOsIb+wn1+HXES+fnmpg1rHnw2VdB5z
qvm5zojvLnNWokLP+LmHEkw/y8qA4O3cJRVBqrDQcIYJVQkPmJ+mwr0X/Gk/XzXwS8ymk2M2ycWX
BKIS+ZsWdqcrpRMahH0o1reb2nWxDRy90lodx1cu9z+FaQv49st8/FZh3Uu1qFoVoRHKa/uztovB
lrsNuni7Q5AnWGprMVjzYbuHY+e6sHEZtAmccSCb2+7DxEEME6OfKHOljLdpNc0kxLIFEksm4RXh
ZjMB+HF/s/ubOVTk9DicJxOY7VEUFEmFcOs6r5PBbSiYTbJf478dGaC+1qGNcG8YtrefSgp1vmLG
CdPMWTv1so8yYlFSsB4xn9CcILLfmrZwzG5PyohPfdux91vlcK+HDHn7wE0uqPEweST1ei7PsVA7
Rxqf9lRNcW9z9qxbf9JO3kK4vbx8ogGvQYr2J9ptvj1r1CarQ9twHUAdvk8zDCELPfsLtmA50us9
7M850Iz33DV4lABo+DsK2Mj3HYcCa18L8FRIXfg/w6/liXwg2FhHaUJeS/8o0+NqcuePdgRHOdwL
VvX8aaf7fGFmuM8w9ZjhOx5FiIQgKwi+RwZ7vt7QQVPQ25QthWWG7KBH74/bVOavkzqFgUPKIp6F
MhGATltDc5vd45KEcyAguq4ppT1rYu9opw+8/FUCZO0QkFF9RByBrD9E1q4k6igciyUhJRBdz2O5
OgFhz1XMLeqt6VbZQcKaiQr2pyR8kKomMbuBYAdffAu7/Wrlt/sooUT7M5puLChc0VQ5t27L2TfE
MuyaUxFxB8S4e9jjxAk/KwFZXMJlTSjaS88ZfsJS4AXUsb9bVbVkXh/fq2r9fx57+ZLSlENioDsB
mJ1tLBIwvAUWigacZKjaSvN28tk5iypvj1TyBzEgoQLh1/qFMrArNNlXZDYleU/883dppW7WgQ21
k0KHGQUSacWPjNgwRi5d5Ie24VD6DcuOc+C05gmuKytyDUoWA/cnreXbUp9A9P9C36YTlNFM7/c5
U2ZOzDVJm9THPVtvGFQdR1ICwnuawE1gaSDhXMjfta6648gKTmFEL8R0sVwQ3SGFR8jK+bKC7/vD
sO0A+Kpp8GQxsmFmf7o92J8Q7A6p/ncsvinLcKhbX8H/lAfQFLRhSPAjE2gfcHURMvhObJNMlPlG
oTIDz7McqFOEhysDZbqaI2bPvlWP0qHG/y796kXhTFT2P4xQ1vgUXv8YXWO8eJn1tprjftPc7ncj
0JfGwtLAJVjsQbH/BbTzi1qEkxYhKGAltyIXAOuOhNnqNEYJHV2CeR1AKGbAR351jtc1RU9h2T+h
EVMgti+5Z/7pv2C1kFQZM5GSypHtLN+XLoafpUaOKQenwx5P9fs/3Zywxdu6lQa5kAOgW7odNQ9l
+oyBCn2KNkatnZTPKnGhJqBgZTrP6HMGmeyQySHdbXfPt2MMJ3emDJicgcBZ5/dFzorZr5JmPOKh
vo+wvXSpJ5CUMAH39i+ZjqTAAqxtSU00E+/EkJcew1itk+RpcbiGXXCYQQyciiXNjTSpfAJEfQom
oSn4iSEA0bLqUIdvvAMmXYpd8R7qTue4e/MCZgymKsTuVifk0XCmGaEhzMRfPfcxPGXQ5CMuyP32
4OycUzWT4L1fPVVMWTq+qsA4QNFgTMrMlWc7rWi1YnLo4FMC6ZTqSbdxYByI2al7D1yHprXxCOjk
kj458cVSTLsA/8QHgui+SOn/6gD9Kmk3r2HItumiRqESMyHg7hmwYa2dNCUz571U+5OYp9zA67J/
xXrk3LzKMcHsRbRNwufHM4OSW8y9j4d1RRbvBUv32pZZBNngo2MEJ5KavYlCmVKDVzLMtqu2etj7
RS90seKP0Tb9feMtJ+NPESGRMq3a6Mo8BAV2TrprusUMNx0oXWiWdTqNroro9TLq3VhB5i3NmCs/
VVpbNKljcsCulmm8fxnYziyfKtc14tiGCiaUeXc7Oy+wn7CAs93FT95lhrW00j08cE4ELTsPti1f
TxxafgcUZnXgTMbHvyVe61kopLuHSKpWlvueTesJrtT2SI58y05X8KhnXxR32ug5U9iIFkhD5YRy
AXu95Wj1mSQ=
`pragma protect end_protected
