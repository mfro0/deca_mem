// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
sjTb6nehcDtHrtqnn7cVDSfy39S30inK177dKWcwSnxNSI7AEVL3AGDjSgxP++DP
nYtbl2bWMW0iJLcwth/MvhXZkhV9SnSNdO4lsfLtYCpn02ZAW4jUysU2P3xoISI+
QHTttYCz0Qtz2rQsx+q6GdpitS9aZfKvKETvqvqJG6e21iB4YpodCQ==
//pragma protect end_key_block
//pragma protect digest_block
z4lWfT32vhVEHCYez3UoK4Yoeno=
//pragma protect end_digest_block
//pragma protect data_block
t65Qhmq5gH1CfhcAI7ntAxwNNaEUW5q147qYie4pKbwonAncSD9dFKRkF7iZ+loT
zxWYLlZ5fLp92GRRoERbDhbX1ylCQuC6irMOGNRE2yg3SOnVYfR3f1TqKPzEVOhz
5oJ6p+NHnio6M7ikjBo9POtLotweo3mgiLfD5nOz2uoM1IRsYl2l6xqurmjM8BZc
JdPrQcQkAMcHHLUEpKAirq1xltPUANMYM5VgruLl7C50dt1PmK5gkUTn31Wbr8cb
fFGi5x6aVudlVZ7+EQPaM1VZBm8gkP0Zh7ka+U3XjPfS7JrcPy7OJ4/CCdQmB1GY
6ZowA+ZcmoW2Hu6b0nkIkXuUgiumtciLcDMMeHVZYnB34WyZ/utevD43GFyiqm/W
imFinR3FQPjQHGin2hIXi4kH+uuzokrk6E7xpyzgUxygiljezN7u6Bb5pTAPacT1
Wy0IkyJjHGwnJQPkhHBeKbXmRt8zGSMrshEtdOzhtwemfXXTlgWmUo9ifLyDEAsH
lDbiSz1K6NsBJ3KnEVqiX/mjfQvZ4THNhojxOi8fsikRVzRS3O+TAXCmLXemFZpw
fROiah9Al4GrXI5dY9X0BambAI9DWZyhqDIZkrOQhbyjgt3Cb+FFzyvIEdxQtHm1
37p7wtoypRK9TBrPrKIRqvtuhn91sFfKX4h9BcKQ+0H0RKkmv6HiGPuKFNK4/lbR
ZLWJ17sMDiF3ru+iYQRDBGfm0piNJNvW9yVXp+ifW2IEYOgiMyK4prWBCYZBFy4k
wHlvsWiRpvrc42KmL+2UEaY0pMVkaLkzVfOzAF/PeorAmgboGZC27TDOAVaNZyGP
zQ/WzpxttOVELSa/yDSX662F871RDK8sH9zG1yYHjj3ITyyuJbjUgDGFX7xgG92g
YgnqQSLJGyj6kreVCVHUWFn2roPgreyeS0otVK1Uu4iTKCN1ayufBzaP7B+U2BjP
84tWB9utg7/KajzNudiXC2fa/NJqqFKtflxIcpaNHgU3tzq0qf2rBQk8qzyrwFLK
2q+wjscbIb+ZwOncDCg6vEg/OgJV/ok7op25ynWCGFhSMRlr+13G3WuE9gfwFDG5
+GR1qRwOfSI7vMZFZOyLPxLdBHuG0lt8sxjuFPZNhvujVj+3ehND0ijJO1FGtBv+
TdE0uhWzrOTQKYoN44hGaM4U4CDNPhq+LJG3G3IUrYiKd4dXPStUqfv05/ZnDAkJ
2GWCoa+PpaHZ7+0HAjXCQAsCZxcQj49zQytnHKKLPeQdmI7DMBPyEhl7q3ZieIKh
SHE3yDKr9Vr2y/6RahYY8VVJhW2vv3SklRpYyCz8ZY9hXI/kEqD1hY0IfBEsBlU6
3XxAtzxxwnKU+6LevWoDjUJjrCSeRda1KpnbGoOTnXBdaDtgQgKLaTVx9x4EIWlR
kUywsW0aeDASAeyqFjxljPocQ2BcR4cQug4lyQba2VqY1HL3oQLTJy8oWjoDWKY6
IuwJs6YruUJpc81LBdqBnitP842FiFUcC/JkFkA9BjFA0+zZFMMfQmq8SI1dta+b
AhYa2IeQqC2dDwpzeP71IdYZqYOL+Q/JUxnSkCeJQt9u7NAciAwtj2sBca9f2wuS
XQhlvqQaw2rBPddkcOQHctE7d3E/157PQLHeF621XdpytI2vW2Fv06wAl9a0upHi
ykdX+1EXV5uvz4g7ZEQG1w2BwAOQY2O5WrNmyIzzE3TSOaVak4itMMhjStW48FSH
zF/8+rkmujT86u3R9FJX/dvVew+jz4g4/KdsvyVJyiRzfn7N8f34KDXOqPwoCvMJ
34BjybnbE4eZeLtmrPOeggl6qW8y32MmOWLyZ2DHghQG1MEuS/5jT13vcmZmxmDB
KosTEUiOCshdvLbuX0cKk3H1iHavO+uoasoKUNu9hZv3XDx4WlKsIpSicHIBzSX6
YEkgiDq1TmG+j38n8eQ+ZUHW6blqwtA/VPdQ8joOm1R2U8/6ivbhQ+dpZJFAr8Sf
OgcIojvg+RidZ6ce0GHpSppzk/m9gsjKlLUhExnKz99M+L2nRvIwgUfGlZIU6osf
JPuuVcnNzKN3BqzlrRX0FeJUrjnuAOElf91fnbcGNwlHkji8ovJAe7ApK4kqFwLG
hyqgVjSei6UFTHj5iqRlCZDf+5wqTmH+AqpKc7A9+UXDUMtJ9LYOBcqwjDd/p00q
4yaGErmnX2Q/ygLETVUTnv++1BP6JRDlQnUyCeO5QFE1s6JKMc9bLUx3CSyL3nsj
VWioZz95lpahFQiwvbhCtYP1IIXh7V+QY1l35TKp+dFRGJY4XOVnLIyCUxp093YE
7Y7oFA1ZJfW6WuV61r7TkHqnfwjSdpqtlw5JQc1S3Zedq4x1OHT/hmiwgVOd0CQJ
n2fkw/IF/jnYbyiIQwR76p3plU/pJmISeX5IAiEK5S3/2cafXkO1q7Xr6XqEGaXQ
4XMiNUiw6lCjlfAnQnNwGDR9FOsxZiq3CThM7WEQ6IxO+vTPneBS8zWZOBPVtjzn
FFjecF5y7EdRCyuoX6AX5LysxBjfLnwHYKA7vCrujBGDaBWIvO5D6CTnv/VfGhrD
arL+1fM1g1buv6YTyIYzFODP+ScynKw106HgCjOVU309En/jOV409+Hk8yrGyD1A
3qhqPzLVECLmlh5+bNSOe4cabLh61HVi/0ttWxTlcGaXW4muPC0kspAhlOTtF6Ah
mefy+1QXr0eDsXpg9FSBuK79UCX5zfXuXu+FDjIRo95ujktUW1qv8sfNgO5AfT6W
gc45BdxJFVV4q7KKbn59V+coUHkmkvisRCpv+dNK4karvDio5fUYufXisc13sm9l
MeApJc/nKy+wD6wD+erQuPrCphwmFrHHD2a0aSIKXqTrluscZi73zfD41/ru20ex
XAGbmztigr2o7MQKCtK2cXrq32CrHn4A+UHuZ9uK7dGz/rQmKTQd6+gIVHi+VG88
vlWGmRVkxYhaaLR5wZCvCiQDT8kxLWiXd62cmgj6L5JqBTCQCGKM17jqS+KVlEpi
Y7DbWLa0K5RRJZ9/YgwuVz49wdzpKxeyyKbB51inXFqsgjiV1DMLPEPdT6ts/b+E
oB6Ll48HQS429aL8JpnUKf9fBKuedr/GUllmiS7pN5+Jrn9r2fgz/jtNCZh2TxpJ
+cbjHB5cbcTmNsXdoCJ5su7JvtJ5tSZ1NbX0zCuhRFRu/ECXRYRxi20Fiw4fjKOw
T5E3S6gK6LMytoCLmZdFVeud4SIWQQRtqUuIPzAEJH8w5DoeSeooNWTrRy1Y2Kej
jN6x8Iky57ommjrYMOD6GnrEOE5e0U5JL2/sANXpTfny+sQMEOYMJxdyXuSxmt7i
f5QJ8mzzknUI14LEopRKmUAtkujkfom45+ITKpfjqFIBjYZ4zVWJTjblCPCnxahu
+x3+WXvwubQWqHJuSGCloaUSofBpBixMlpPdW8RqWBeufH2p0GRdPLy5OMnRUOoq
jI/RS2wT2aVIXpSlG6pe9nApFCU5c9sbfSDI1d2eOgtK8SpGzCkmQPVE2MF0JH1p
o61lPUxtU/ezGRR5pG0Wfxq1TRHLjkdEPK13x11xVv++5jMN8aEJe+BAWLWmjcPN
56jgGmefxXlvhkLO/IBRFEZzJbeKsHQS9bVkFkZ1oIUkYgthht4UYOqJjXojv2Lg
StpDvJmbtY2Da+cqoGPu3cDfeYq6till3d2FqjbJ8d9o7DgrfNuER1nzS+516g7G
bpG1temY/5by3zMsAuX/F3oamTJ+En1GejFkxB94Yf+oAy09xS4eThvy1RXdLZPT
PFcDj1RtQXWbkjj9on9VayL+G2DO4MaXCMcMhRr1qL1wuRFB/Fr7Z/DROCJIxzVD
WPKeGJeBlIoOmIk2GS7sKwKVMCJZaX/8nCC7TWIhfOCFMXJt5em0cmLDxTWitKjY
gH1IkZ+X+Rh8iQ+BPqY+xWVJHee21rXOjeU33eaE5okHZj6k1ex7/2uC8F9Pdq65
OtHZtWOAFspJDJhBotR0+qO0IfDx0ZYycm8zAHsI8yjHbnh5X0XlpMzICpVhSEYX
zyz+QwmggRgTc/1/InjxClwsEWMFjkm+01HIvP/syZR2AilLg8fAl88QPzioEd2A
hvv52owK+rplaI4VWyfnKefi4B/ToWIoBBBhGlPh2yNRQo0XY5okF+qCwmfmnJux
tvSibuRLS4Lf+szgzXIgC+djo6b550rI3Lxuj6lzE2CS5l4uDEnRDJYPONvUO1mB
IQCOAUhAnqQUZg1FcLpK6gi5PKO6uIROipB13vewP+mM5Zw30RLFfou5V5qMllKv
0Ri/Fl9TJqFU5MWeOlaQ41YXHoAfn/EIsTbk88cSkIn/850Rf0B5fcgK0Wwgwi+h
HMcTVGG7vIT/h7SeVHp6tLX3Nv2rpeduOJ2R+BFop9CujOPDoXfNGVptIAXk7w2u
Q+F2dGkODPYyok8emUV6AL306+bqi8HHmYhLWTYoAYbsowBw+wlVMI5CwvFBLYos
2avS6DDvIp9XFlCG2gAgjv8PHCA7/bKSRFEkcwFenu/ip9uFeoyWT+KscD9Qi+4U
dVEtH+alRpno1cwL38Rw2+aNg8jZ+U38r5qlsGI8H/UNT1/WAk0TOF9c+bntzASr
oG8acDV5szSArU/NJKjSATwa6/4+tPKmpOaVxNvUXfyFzBYsAUoXcoKrw9YwwDgD
olHn4754M0jKBS97iu6FUdDzIWXaafuaCOwxDXTJYDmIQ5fZjxkXfIIDvQUlEI6h
ytAZy/ZdZ/2Yl5dQwa4o+8kSHbWdGajZwV6AAmbYJ7OMX8F/CxFLrGf4pk9K0+d3
YkKQoZuiPXn6X67mBWapqC1/9FfhnkD8ONvTrCfzPcaYN2gNHZB05Im8HTUxtUSq
4dmLBrn3UHhSuA04WHIEMkcBTchuQhce0Um5znRx/9PwDrFpHxdrka7wY+hVMdIc
7NSVMi06E1imBmRzOha7TBNSmFp/mLXE1bYziui5MzExrQEbrmkGS2qjTh+lhC/G
HGUE4DZ/I3+PSbcycmLhJP215qUzm899Q5iaHo+sWd5UN9EbcXn1MIPktJoybHVd
zBSOlEVZ7cTzO6SuQzler7E/Ariu2dmKgh+avGYcYMX96yrGyBSmuMH9fZCKyyN6
QZWk3mwBCm4EcBpBg2ZA/EKCd/5KowOE8BPxIZzNa3skSYD9UYgS65cEqyIhFlWz
Jb7TXo/M+wl172/kNIp8GzuC0/DASvgVXCcKcq+aMKlTOMNER0YdlGX1hOBQ1BcX
EpE63iP0lFqq7V3m9EMIbl7QoCWMjVib8JnkS6oY97iiWylhg4Ajs3/WzEEExquc
w+DNXlGRNJs3UZ3HQUSGiQrOWgfi7dUm+Fnu1IPcX1m0yWe9axM/uVo68UU7Hcng
PQn8jXSRMtFvKINXmT5xY0mOUm8EYxj//UziMP4E31VDLPneWcYmL9BLFfa4HhbL
8tUPqvZoMKLMDb7tTDpFhCYUgLKR2DeW67LemDxGXvawQtv6IYqka869cuBaUshK
h+JWUsLWytIM1NTvi0pBfKm6+Vpkzwyo4n2WBx3mTsps51Gr3ZoQBbgfnzUVZU/d
Iro9rqrxFcCqFoYuj8u4hYVnIXfLFZwmkswxbwvjDjIWSdTNEojiAgDhnbsEf+7C
jlhL+fRFWN5pusqriBbmcpm/3PXZ4RZMt5Cf1AdzTYQ3Uds4XOiA9eCukl/zV75f
TlS2gylKt3HJhwa+X1K++VfT/4TK4ni43wfj7dn/Uromt/AKbyrNDqKn/ceUqIZq
SEz58eA2R0kXcNtFIphgpgt94Mq6x8/+9P8naMKgm2X9NxC6eTwosxWqj/1DGa/r
SMREuuzhK99IZW/lUfreCX03h5ajweGBx8gHfev4uAz4xTiSd0RZzXVKP/wYw9ok
wNXnTA366t3BYRusbWTQ3Vk+M7VAnVRNtEbL5TjA/GsWeyvkJMCrN/Iye6Klxf4m
5Pwq1yKXiY9/ZKqdRWiUYfeNRLGcJ1l9tw4kPQ1pWRNEIam56PxXuU/9SoUdammn
Pc1AZqTxYDbjJNDMCK3gGGtNUthE1TvROHwheTd3UVBiA+S0tQPxpWwYE6vpJxo1
FQBhUW7VY9HHTRr80ZuXXBH03TkQa+yqs3CnfFEZsIsGjcEjZRWL1R3HE64GUT1K
Mu5xHlt6G2RmLIw+Sa1OOVdEdk9fv05SpVWnarffOu3rhJnOYktL5fkpfPBOnGOM
UCQ8MHlRIPNAdzlysLIvVtDOyC9/tSYd42Vlt8CMmOFFB5CeV+KwUAXpYKjWEwV4
tHk9nv67rQ4U2mRk1VflgT+BLxV0qwSLCaxS+t3xwr5iqRXCZDP6ksUWnDTjB1km
dwzxcvbQxjVtmc/AHD1aDL+fPwI3hwPD4/ZEdM4tB7Axa8lPyJn1pbK7GphUsCx1
O7+PWz/Wxdrw/DdRYHLKOErYTwZu4vbfoEwDiG54nvE/9gk/zMudrvfmsc7VyN8/
1MpXjLQ2AXSMW3Fszbre75c0lYjumi7WAO78CZc7EjrJqh4Al6z6HmM+smDj2hNR
YfBNh2H1WrjX3fg9/Ta9712Nk96glrmnotTEWsjoGEIXEHeITMpMBzkg0nONhS1N
OWbe4gPwmFBsLg3ajnMGrmdgp/y6cnEeSUC8lW7EallSD3OaGkePCHhmyyWCmbKX
RtS/pW1maUOvsr36LX5Gw6HKCQWfaj028syv6fdOZhlEZkQ+tJEbkt1h7ubkAxDV
gZfgsDL9ntu9BQfqDEkKG+w/lbaCcxD2H5+niAT0aZZZTwPXu1yyL/pbJkFluqBf
F+Dc2RAO5SbvPBnaJMLpvuxLpQJt+4BYoFIKtyX3+//JoKlkQKsSqZIvD4lz02Ux
n7WObsTFQejaXMTO3xaiDfxaI58lqK8PzsQ/EJmc/9xM9McJIN6yq6PuXiP5SOpm
dJnRd/hIDmp56dBwbzf6bCn6e1Tv0x3wztcy2pNpUMZTKSqX6tOB35Rc1LH8nEhe
1Q/dNQAhdFHrk7hvfrtBknnB37kaWlUwJGdFdFWfCuqZ6FJkp0ZZmU1Y7qhuvEoR
WHxubpv1VjVHYdhHAY0uBF2AiLTq1HfLXeSIrKrWeVYKNwkQfLtb+a4oOkZqvk62
HNAVodqV6XuL1GvP0H/nfVdi7sa/rSpAB/9tROKesDL/PGZxadiaD25K9C2mjMPi
4wZzABqsfKcWD6eM0WZSwSdEzS3gFvqOLlHdofuFtj8lbuFVqLHWCbPqDcCSe/yr
WJifEe5cradLffdzemaLm/rffzK8HcAquEwadFhwvXjMsAw+MVSFJuec5Ufzg8N7
NaX89YP+GznfbY4WX8EEWnLcIW9MHwO7w1TOpfrbFUwApCeNdvNX3BkBozoqkLC1
zU85vQUzUmthGYZTwuXM2Q/Oy2xjAivpZpBR7TxeAJuLKob1+hXVTnEoe7iK6LRZ
RG+MxqbScHR/XMN+sEqXqyuhaklJvZEgoao56OFfhAWCSZz6oHuxi4lHtPpP3HUB
JjsyqdBIxJ2BPNykflHUFnotOW9XHjiDSHIpQF4MlPDR24tgwL7YhKgrIR+ejdW6
izhE5YpLcSr7N379kVZ4b0AImYt7yAy4+FHRVLr8rpIx5E0srGNV1A/aWM5nEHXw
JznDrk2x7gX7UzOzlaKf3TgGGt0z1w21qFQfN+bPEI0En/br5faVojCMgBj4+Tcj
9zOqpOm2UbuJOJtS/ZXlqdWKvtdmAe5q4kT+TIvWTO+JoTP3Uo3mojM1SXyhx7kI
Am9qIRZbcPibhEPRFp1jYqWzlkEAXAKSbuNuzDjNtOPPs4nyK6Yd82n5e5zycoyi
SieyDdd/yJPvDx3wdc7aG3hTugo+oJBAXqulBo3oE3FOb/6XXcxafGVc7IAP1Ds7
9cHbxTtlW43pSv0So8VCIjFlhwEzjhLeWp5r1c/YD35KabEyRqCiwpewffp0+Xlc
KKAW/+UCppdO+CbUnxDuQ3ERwxb/7fX32PGk6hbC2IVzbtujTkftl+JoE2o4FFYf
vYhD5we03fM9vwkhKQU8hFCgzG8hHrkiNWL9SQ3nFr1SFvivcxOPDI+MJMFjqlfh
iNExL8UQxZOJmeFJn+xtmgmpVg2QSj160Oar+lSWg0YhJQBxXJG1IKqW1f5B/PIP
/76bopyXsS7pQU/DDGh9oFlKcHQKbrf6GJHKiRKYSZj77SjQ9g82vQBeeUOuRaus
MX4hkbUD1MQrqE/wpl1tWh3A30Bc2Fptqhvr8ViMj8YEhOIDEBjdpwIZjbhydDjC
EfNmXaKbC3PpYeASMIQOj/zBKXSMarCTT0s6V8Sut3Qu9WrOtZYysLoFO4D/gz5m
h/Tfzr1JItGN8PuMqxmjp1XsWDTH8rcFd0ijAZzfjocdOuMCs7dTHqR8Qgkg15q7
S0gfxsSaBpPNAmJV9iJzo/GZoBU6nqQ0sANULiko/d8uDMY56bbLpmwjiD+1b8gZ
SfCJv6WUDptxOvjWE5DO/mK4KG98o+1UYqedo7OC8iZMoDKaalAeQBMgPGstXZe6
jpRDHbAtt80RaPVTV0okBQ6Lxj/ORaAiYtykf8w5KscPAVRNwfUmTsGhMq3Uy4W3
bX4nK5UIWyiqpLlWkYRLeVST/yVMSCitZMj6n2p+7hHe1h15vTKffi7RSDxkxHq0
M/spmIw/vEbD6pHsj5z/db7d/+j2T0FX+20fySvRR2rwpyn2MzFE+35dH9XFFm+Q
3QZCM9H3P/aDUs/OsEqXRRDJrdfASLcMZ0E8sid4j7iLojY4bympyVn8HZ9urtix
CiGhX3IUsEwVGbGFmanEs+OSk4CaWQz8NtZnXPHSxuASyxL8vdAHjJl+XCQKGRuo
T5d0UlQN12sPUCZ6AURc6HTAUuiRPZkwmcRrd1vPprMkgw11mFVfTuEyXtn6swvu
XDJQz03GH4RzERS8fR84NCs3jwzaOaQq9fMpD8RbKcq8U97HHCEYEbaDnggkQU/5
X9fsk9izjJuvLhW64ufyhZS66PIpbM/TJrlj28N3lI02EzDOjUTryIYSli2D7pjP
JpChGbv/1D915n0Af7aGzf9jN4qBTeIMcgVLC0hYjdktI2gZoKBLAkHpkcvVMZuE
0kerdecqQiVYuFBcZbwql1jzqRKPxwZi965KpYdKxcteixC4xwEA1J51ubL1XF+d
a5hZEbSrbYu6aEKASJRyGDp+lh4zPLyOoG/+eOV7r5C4BVUhxDMk3ci/wrn75Ahp
1CmLovJiJtIwbtDYrBJ0ZOenCszQvfUo8IksCJbR24UVe24OeO3X+Q1qQcgAdloh
1xJ7DAgs9+nEgO3MoHKvOrh82A6QDDpSONI3c43pf4BiIcrBIPJywp5+FlaCYLOw
R3wqVDDLyGMnhUR8jIQ0+0conPN8qJ9Hn1bOhvFA33yTAA5A0c/5vQP9Pa5wIL5g
XVfV7ol+idPsEpprlhHt5U6Aw6YdX2utvr0qAz43t630VfdmZDTYsQ7rXLK5bBFh
mPvxQPKxQmNXzzgIWzYI2foE8jw9/IhxhQ9m2D1CRo++X5UtcPX6Cbw2EElbcQ2W
2kSBl8WBSgn3hpyf5EwFNUdvCx0b/HHMOvv+tO65nwaLHXPfWeK52iYn7eestSmL
GVOJ5UPd6KMfJxGsdGuW1ivdX7htiQZ3XHCOoB6SgIuA/blUZNrEJHLPqkzD5VVi
wah9cyrLkJXZe8VEKIJoWRu/Iq+96CQfMbw1n/zx5Kts7sdEIuMSntkM6vbzakbY
Lzc2RbDJ7+jmXIMNvsNCVOffC/Pi7GVwRq7r991GSRflimTp3tjPKihXNsotoQUm
pUI4Mgs+rr7B3k4ilQJ59N3AyUkvD4oC2sJd6TFN0bMI1HQlVJQ87WPg5NQY04wI
3NhlYmEnTD9uc4U3GyrzoJjhmUiue+pF6ZnWlrMtn/pLuahv0DHgQdkWhxqNj4uP
iGz7DGCKoO6JVkyzErFSAYSnawcBEl1uPEsMMwBzq9zj+4HEhP41FM6cI8VBVg3s
F1tw9wUllZeu2VUhM/lURr4kr6zj1rXEDLiwTvz0dNYM8NWwyhdTTK83pMQo37Mm
/OlK/3G9H6mJ5/j79YZasZodKokg3fREk56ABpo0Tc4Bk0+ojPSuz21yqQ212ZFg
aaK1Ax71aXjSkqtbFNi3hitwa21ozT5u7EGIBNYvux5ukmdy2P9stMI5nlxcP1s0
Y2EUwGVcEiS9Q3m27ok2r+TT40ODXGcPdoFot8cTaBxVVYDRLtSNjNVcZ8ZGH3OC
JVpLMdnsU2zeE7qDSSx4sAR9GiPmI1mOHxm8cC/MO6EzCh/U+Z+WsLrylm+JM/j4
ro2bGZ2FpGWbKDhD/8GsYsuLJ0jOmGU67ZQjkKC7SNFhY23+U2PT9kOon2R3JwTK
DiSBtUynpmjyvgLsYWD/DtlsSZ6LxDrDe5wUXleWvQfYlqyAPsjqWBVLJulNeL5l
8ID2HQRkCH5zDufZMNYOlc+qyLqZO5CMoZPiESF1JUHRKIw1BKWTEnFQZsLSxcwp
3YVTELsZj89T88WMelIQXTMH64pSJiSMtcse2EE8EVjZKFQMQ4Xop5aQouExmEpz
6PWd+bAobqdyHypNNQBczNwy/SBiafzWBelyEtgftsVbSwLONwaFtA8D1zRGGaxl
XeM0Ejo/nLP0QgBLBTniXAvp0WDS/XUcUFKHprTtaDr2TBIyKRirebqz7wYtSzLx
q/m9cFMbpyAmGzZDR+8SBuY/N7/6Eu+mE8SPBOn0pXfEzciNuTgp8daT6F0HmjuH
F4iPR8S/pIJcBNfnkYKLOaxruYgMyQXTeRaAICbhjFv3b0vIDNSN1r6XrlJ6OUPg
IrE/Y4j4n8NQlx0/mfC4VQVRsY0CbOL+7PtH/yUNl32fbEENSnlv5n9MnodmTjSs
HBUFRRr+2o7epelJ9gAMLzXGTKlwzOASvVcPKyCgSZ1BygzHp4T4k8soFB/SfbTz
achTbmtp9TWX3fti47sZZ6Mv0wNKkTULJyUnoToY2IxApZfJluKg9dYW8O7YYwli
ClOhIxD/BQiIo4E/3qOakhda/9guJnjqEdW419TFY2y5IfnjRPQngmeNplbTgDeq
f8PAOaDIja8lmjgp+R5W9F/kySIo5TwlEqtV/n6FpV9E4JGsFpEtfBgmQWekJ9Vc
yOmVkWHPkOnjT4Vj9VMa2yCO8CNHbDfJGKU1ZbiL9KkVXVWzU5WhKlrgMKw0apZE
Xvpc1rDPhmUgOw/iGVHYxFSR6gFmRK8iF9fX2yjGoejPXeu4AqTGAe4sWNgQFh8j
mAfHq+ctiZHGog3ZspJ5I0bfLqlEgmcPF+zY5w3ZydhydHWmT5vm0viEm38Csy5R
lYD0c46cOtdd0C/rME/WTENAND1P+PEo9Tr+ujbEctk32dSqHiTp3StahKlk/ooT
m53F6ajkj0XW5fzyHxvkodmvVRaTh/g9cyhniHqv1yYpMgU/bHdYnYwSoiQslwQ+
SIpbZlVMSLJWGpfWAIZnS684l1ruNkWMzdv53hI7XAVd4MeCALqJy3TOgwy+apCT
1yLhiWBru1tRmE9iwNZ1VKmqNFiPKWS9p5mMCmX9j0KE8sz0TMgY7o5iCIgbIntr
G0kMboXADWrAIfgkwAvhdZikn5r4aqcldRWnO7b9XJMwwmiMEGXJytCvVkY9uWXS
U1ccat4O1XWd0SsnowmTVjQE/toyOLpIgU+w/RXTy2R+u/49RH3pNeG/Q9g6IfIT
pJRzoZD3oqi//1IGrHsRUKrtsxpxM5Va8Qn/YWaB0H+GNhrNBbL3RPSMd3qMIxIO
uH6c2jt/FNE0gJn16npjEajTha5dhV2IYWHCtbHL9S6wC/3kVjZQUQuhmHcWcdnD
9cvX2DsEbFBFIaCjBQ1QVzNBL2b235H9DPkllckwKMYrXz870xguWI+Eo2ECmiIN
Yd3FIoFzaVZ7Rai3kDyLs+2AXJ7bWc9rGBC3retKsuYh57aYe76ikzBHxzpEc1Rn
r0OElymtDVAbG5/N5xhjCfocAYdzQDxbAN19qHS3WBV2yCpFyU/xjqz5xBEKPt71
fyTbPGub0I0paApANc0F3EZurSLqzprP3BXX2tj3Nr6i8KtALNm9YMuHsWC/khOt
1M41E2qf8Q2qdrmxzAhuiuQUjl0UiMhcDUPxYg5rwiqPyydeTphj9cZ/JkQmT2Q4
ahDJp3+XfmrYs1V/s9gR3BGSzn1pGXFfl+vGceV1SjfGqG7zGSUe73uaYeW6ppx8
PZg1wN0S9wg+w/+1JoJHFVibribJG/paESnBrzr5gC2r3N9upXHDIrOO3aIWDbiq
fgalXFxkxnBfpLMcfxKbnj63HfINjgwhVm66ZRmkPk2PzNS8lS/qT7jesIPnAx0A
tBRgv+vgTPK3hYLA7Va320s0p/KFnLozI2E9N5KTrxLhh5JqJlD1DNDhmF6yowMO
K+BGXGjsU/vbE7skXGI43CI0EVZVx06mFgsvHczdqHpArdIy9vvG9mJu9gL3isee
Bzfm7IhBCm3eGbbHfNRoA9kQ74f4bs6EM9Ev3S8NBY4D9Kl5HHfMBQ+7c4phi7e5
sY8UV2eJIzZp5KRkHQmiZUEgXs3Xfj/jWFxOp2ii0vy21Pa3kh3XJxHT1POWlY0M
13XIIDFR80VF9C2Y7lxJCR5VuF9V4dBEXL8g5gdVBbmvhmxkxfvM21ADCfgN+vIt
MD7VzQzUUaUfCqVSj0cmV4hoKKp84DS7R93mC2bpwGy4kSy8ukuVknz/h2BOGZ4U
YDKtKrZfwMWyq6sv73l6lxZTZQgBSVpV2Odvqmb5IUY5AKcA4KoEjBZna/Aly1CA
K/7AogaMdUbMGwY7QzvatUkz2LOMB+BdbD/1T2JAkWcOYevs44sYztP+aT3QKpSU
mluQtchvLJrOzcbJGx/NFcSgiKYkaLoD5i5CF6jcCLb3uYM3M+F32W1luNmQc5oL
lPLzGMspjj7rMQIPDa+Nt0CiwxgAkZdKMUt2kf9/SQEM88SIHGJc4Z1ZtogTh49N
L4IoIzNJhCfnwiUCig7pnKZalPtxsm56gjOsXDNxaqXK9ami5HrwP9iUNcDsaZ4u
cskRGMN5INrqLASsyRtGylC1Bffm0C7t6ciFob39/uii2J18uad9dXVKICd/64R7
RbotT/SfvCN4lNMVmd5t3qcCEmEeNhpktz4xQccCgCpMUU7RtO1huOjXoAmh1FtC
LmFrBDPRCHuIkxItUCiUUQE9d4tQ5mF47otqp6BpGw55j6paSr8bN8Jhc0W+7SBF
rLCfiqpNUIBWpLwNIPQYSAQV3LJhrcnp2PP7OBy+DxbXw4HDtIUpjh5lGJ8onSyF
/WkhFhMS/xxlJXMA+Gf8D9fbaYtz5EBZxz0ZdGig9i6jOi+udeYVn1N5qN9zg2VQ
KLh5z7qRzlM/1/a+ekLXiu7+D5YQkAv9INM3TMZpH8ZD20PZ41uWrdgluYthtStd
kpalJHFEaT6We6Z7HXxsabWNYynRmSQMdbrgGkCT4Y4NRwQwhfOsQfmBknlJog29
dAVaebRlk9CtCLThArxHJsAxSwsVIANuunGsxKRiDzgWI9OlXIdH5Kg8pXWX9Jho
OFVGqvUpcpUiseJ5y3uz9Ym0KWIwgiqjPGPzdy147A5xGnz1vSxu42Oyw6fEA8vU
91k5e6R4fwyK6b/zC8I3ZheJvG26vS7g+93rHDlJXhhxBSUzRirDshnnQD9BM0dM
WCSPcqairdY/2KqmV2rEAbpZxkfvVm7ONzrzdJYz3hV2a2jl8iR7+9sV3arypiFM
wy91ayXci9v01eDzT+pNnOYr0RkqGvs1M/zhXFL4Obacw1WkpdYbSra5eKMTSi+Y
Zsxyr9NxTBasIQVQ0rnt3hPnbTKU09VNI6R/AX7Om+Oj3O79l2W0R40CJcYfY2fY
39TAHpFfx9lNgzXhQMTNHvWcEHQIl6169ERdzmMteRsxP3WObcD4tZt/CJ1N87+Z
qUUgMmZodvi7ikMbtVPSKi6IkikM5DFw9+83zg+EqaeN1I1BEJXn0ZBPsjneIrWY
qx3x1yv2ag2wE+e4fcnvzTqknGUEh2vSLj1bH6ea5JZnsitX3HXJ7Ex3f5coNnkM
YUQ5GyLBnZfrB/C0pbzgIzwe9HEzdYyctNVdZztcoRL47TS4+GmK38bYh0z1fyTH
nKZ/z0VOH243dPmlWHLDmHqPOMbvt0ofTB808iG7iM7tnOdf0KJbp7JcamXD36QK
wdJkQTyMth5BymXFaKLYJ/w7lCneWdtCQ6dpd9upoCZrqODF1xJJSNMkfc1aJPAq
MRxVDjsHg7H1i3j3EL0rXcWFumkaR7jL7VrAZxawdIYxG5LYWiW41MPqorHlB7mX
cTm9HBhy/HZqXpQROPuiFcCCC4yESCs7mZxR2cAzz06Ce4UFGGW7IiDSl0TTI3ix
GAQyNvYTg+XHhTabfKPaiq5OOKA2sCIOzMV+JvJjzaSQk1+K/qbY+4PijLQ40FNo
D9MsVXDKQg40pFjdVqguFKv8+Y6qkCJue1OYqb3QoFJM5xNQu3zOUriLFp46DdXd
N+qwxMklfIbmDNCFZltLYgteGuAQVIIa/eQc7yYzeV1+/28EM/Ms1UEwTf5p3WsF
PR4tl+W+gMo7ODgOuFVj+a/aXdIrPUDg3B4ZcshbZHK1zU/aFObbXxSmR3EXZ+Yx
1GVvkX1S34tzMdHnnsRavob8xfJTIolw2EE3RvWuhGn9XEq7ON+1fRbmML3I/7tt
d3sOi9R4eXZwX4ElImcPNcKrubgsu5e1XiswfeWCnm6TJ1IHjhC94eH7N95ZMMcM
36qUoLXLn1Vz5Oljd12Xdqjz4s9G0RFLJxI5h6l3WjYx+h2Ylm3JMEzO7vvLiiXC
N9UCDMFNa7z30/ysKqsoaLU+AEBWWlpYANtZy4rLElaQ4Vj5a7GC/y2Z8kdhVJqy
CFZdPl07rRDQlyCqF0tbt3fXiedzy1anHKjS/y+TKrvZqcMPc9ZIWmCZVuyQA6gl
cLeyGEeGWWMtDXuJScifzNeuoUsXZby3Dw21zq7H98gcLzPc8xgzJbpwTVdnoiJy
7KQOT/WEl7dnTr8P9sCFf7fHGpk3m2nwNCxpryvzSallBmNZKOhgw/7EJgUaJLFf
eepTs19/5WakPajEs6V2BAdXOeEYiCTrsEvrf1CmP6FORO9vdAivWF+8bvUMIELo
89rSG72kwuUl7mmr7x7iGu+kNSCv3665bbluRBWc4WdXQUOw2DgELCosO3oGZfYM
WRmFlnU+403EZ3ih+PlJ0J1ppqKDqnkzn12TS9Yhmdlbl6C/oehTA31CMCUUbM/8
HWe1nM0hduj97/9od432OFG+T/OqUi0kkd5C3e8UZH5zGC/DhCzeJ0Hr85GgdDso
EOTWXC/EA0R9Nbj7GphHnTv07OkiVC4Hkn2WqaNYthvfN4I21LFagtvGV87WgysM
jIcz8ERa6lUOH4lcRi9/K97uAdr21qs+eEL8pQQEtzBONs2Gh+JaX8u589blav7v
eJh+gAtm2pgF3ZLLpTCz91/zFaCV6BZVxX2RIAKcxIiXhwlqj9djsA1NJ93KqPm+
tG2RXOr6kDNiNeZDOYejlyuWiLWrKRaPjSvSsL8dj3cBapwwkb0bPNFYC3IcNZGT
g7zn08pJ+3uruNkLvzy99ApfiOlhXNDO5gD8gBzTO3LPoXVzbwn6dQ8vnqpSl0uZ
BwZS4okJTkW+L023260R1zNtE5np+iuYmNDbWWrhqI5ayZy7+wxvewoSrpUIxiwH
UpQaKYOPSbQEIf7ApTZ9WTQUDqfLDeuIV9R69R4BoWezAbN2S5XHTBJBr4H+lFlo
/31N8q3P0zQf5y8pmY9EbUdZHjbm7bZabTjGoAwKO7JeVnhFZflZFZx7EQ6UaIk/
kLlgXUHqmLyLJlpx8DY1ysbYgtx/VNh9EobyU3No+t3vcti7Y4emkG4DkuGicIOq
4VAH/ZBa8ZEHyuXnDq/TPp6nlDypsOI1tS+IE7rRJZLln/w7PjVudHHyCF+on4at
HO3tWNNRpFzh/FOhyqXmzPECddpRhNDdSaD6jNM2Au+pmh39HE0cqvAl36cPSoY4
ic8i6K6MZLYfZsy9QhuplO+erp+2vBpXMCBgpjWZl8U1tvQIx9iZrN1Uo8WNSiXO
aMf4QiYxLCzg6Z26STCM0aeOHdi2jGBztC85Jfa3AtYqms4lXmv8F/ujAdObIx42
y554SVVP2eOjZ0eCPpGNp9VEpJPT5sdTIsmMt9CFwggoGri1HKKE1/CE6mTlb5M2
YkwF7yIwYPkMlkDvzmjFmZDqOj8JwbBj1+C1PHe0zUddwKvzW+sz6IrEag1RhMJN
JY45fNcZHqQsltchYO/6Zs5XzNnoIFjxr6GTzR/MoFnK7VLeJspOAS4IJA7RfdGt
XZq9EzKpZ1KWaSIO6XNEKwOK6OC8vBhbc93V8ZcOMAMzPJ3Fuf7HZese7ZtQnApU
CFWIbLDn9DH1hoPs5RbccyRxtyEdxqtMXC0V5jm6JO2+oFUMGmTvx2SUR+tXsQC5
6o9y1C5V1gm7FGspYIfmm46IwJ3owXr7ttiQGURyjLgszq8Cq44Dd0dFU/9Oriir
ysZiwYe5jtIuffLTGknQE6JEMlRk1/b6kpN2rJTgTNXeOlVMFgolWjAd7vOUMMuJ
QkBhsumO1evjKLLm9tcqX+V23DMySKAoGcMXjJzl+2miro/CwegF7UawNoDkcDpr
l/3lq/Dr5Xiy+OsfR9l7//fp//dgAahadKSoKe3YYpEdGXau3/yFpWQ5sBZCZrJR
E+0TwTlsL0R0OGOEOdRQZXv5GV1rZbFEuywzJERl12cTVcBJbhTtQ5vJp9kifnn2
zdJIoepYUCwOPqThtR4KktlwKmzx1sHFiKGF8qcQaWYEgI7Ea054f715NP+DQ8/P
8B8FaoPPkA66FaEpEUI7B3s8cG2IIcr5OnPPk9aCmm8uapj32fBRP3sMgtiktMPn
DbRHdgSHCHmgR7ue64rl09m44AfOoYeos8bUj7jxCXjBGk7FMv7LsV7M0BVYV/lA
ZQ6MRsdO4rr/PxQzJuhNiwdATfq6M0RLFk6b6mBDJIo3c3HR5AJ2cN96mYKV+4UE
h0gxNp1xjL6+uSo+hxRY4Kg+ivfbOjquc6qXPb3P4HjjJd2m5QJD2DAF9ARrfHPE
Om1nKZsNNh1yTSlO5rdlYYyNSAoE2T3FhNVWhbv/0GtruELnfQxRUvok7Ou+/OP0
Fit6Qc0HuZMD9D0GiuLfBGdTPhsiBiLz8TAzqpUovXDM6ySHXELItuIlzDqC/ghK
YDRlVZDTpuYtc8n6kOtg0L+MoxlVpIPEdHuhvEDNDx085Dnu4FluCIXVy5j9z9qT
7uy83mWrmTBSG7vo90PH6NJqMhYDyVgml7vL7/sumMRzOsICwoNJgysjBA6+7TSx
w/NhUCIcvMjCEP9v7Whnisb1jIoVjXDF4iSzeCZLwHdaHdGxOrT+Krc/KdSO6q0g
P4bKegUUqg0gPVEDzwaT/9kqdDokWrOlMR9pGOV2SXwP1RCLbTAKAVyOeZ6iypoI
wACubZVtKhmXicVHegpPaY7/wRz2yY1z5YTj4ez8xJBBy8Xas1ph3GiN0rBktp7A
YK/yGkRRKP+0Htfe7N10WQLTBSi4Cgyl8LogmmV0aPjTNa9L4W6YFm5e14KGOs6W
4fuyaSwVQFWBzzkaGd8XCNSvgAz8aZMeAHReTw+U0xv/CaFKdsrXHnFp6LYnFeCt
aF2EDAcV/xAPhsJKPcIFcu4AwMfR0Pli/vWgN9at5bFM3jMvOHpFZ7etebho5rK3
p4r8Fc805kvmfCwsO2IXBcJHoYqFyptI+K/eSR5G8k7/XgQAfLU7d5ZAIKlz56zz
e+ok0tHNYo/GLcqsOZNN8K+tnC7TZTbGYuiQTMxTMH21tntfcanmG6aTmuoV5uHA
LyVuRvgNDwF9qQNWuMA6UgXA0tUeph1W3/GwOTg+ewx5tvMXuUsGA2PV1PEga0tV
4tKGEM991MEQMaQ7IIaV04rpcqs1suKGzbVYXHDkQq6CPKJh2h04Kc1qTB3Kv5Cr
zEP1HnXuSgNr1HAXQRmK8+AdyGaF4KO096kuN8LLKQP6ZatN/MxFQbMeF9rW3Zyb
YmIKJgxUgJVeeqiUrENzHlRqrv8y95zjel1P5dWy3iGIiICmYf9/KfSohqAFbEAt
DCJiSMOzsJvZLD6mPDLagUXwUwxeBZPjtWypzWsb4L3QUMMD7P/rPNjxNZ1oy2kZ
xjX57LTXvD/GGpkNlFokgZ6nl8nI2/89Vfwgb/bRnbTT24+oXmxV4Jz8RnS+wvHA
O0aTbh1sxiIq/6PESloEkFkMmtvJolqFqYwpA+5/22zgIOwT4WGGnaZMtd0AZpV/
yTOhFi5WDRzSO+R4IaWxXRC4CnsI3COmtedG8GZidPR12uNt0DRPenuL2vzYQJ5D
5D4daH96KB1KwYcHz16JuGZURdodj2/4mnOpphzLbPDhSySWSsCyZiAclDvbyuDT
EL2BLp1/1XKosSb2O3vbhLQhn72elbnmAWUWaxZ/T34hL02D5bEw1AFQqVU3PeTD
wM79bLOmIVRGF4M3Ee78WhOwDKkBWDKtK1S7SikGYvXxyv/a4265xvBFIvQJ57gB
uF5zRjHgwfpCdOgtMgXhpu2BK64/xENS1XZEeIEDhPkmTVv9oIk4BtxKNybwv0z0
RcAgld74Jy2qIhuzYCtPDroVSzma7xRZ/40r9pYkL5NeDcyfxjkhWJeRUUw7COfU
ncaPBGKA/6RtCXldYnyWRtrpR7TWZAg87FizRmdb+1PMZPKPjUAQFB5G/lW2OqaN
DxxiL6d6IF21aVgv4aZCsTs7FfJbVmXe9PQH6pZQ+hFfwx0HKa4tbozKozXwKnVx
MG+O9riUxm8EJ+DMuR0entqX4cZZG7VQBTcP83oH3rYcKogXUl3qMX9N5hVgtX4O
hUHwReJ+fsdSQOjdD6MegH1XZq8ZrTbcXHrEyEHRZ+Xf/arYuJG+Ja7+iKS2LT60
1Q8qq6KPr9sMQzPzvhZt7zXgzsjn/8j/wx56scbpNhnm/l/N2UuCZnxhNVrzXdvA
5GUebFIVfhaqHlNPUoQ08Y+771yoSZXBuzpt/c1Mg8y3JY4D1qHxVelEv8QSG2Ey
UUDbpMfG5yYRBEGwxtILrzzgms/oCZoGtOYSycE1RFjn1V/g8bmERI2Jzvw1AOjn
qstP8gZ2TMisFjv8UPZossfc9G2bkl5vNy9FdIzk4bVsZaKU2Wasc3jp7zFQkTeA
vCD+sqdGB+9qlQSiOubs5E+fheQ+Y80rGr/wSeXJ98fmiFYkWBx08/eOhUm3O5Lw
pzqDE1d+xLTzUlWMBpFf9n0z6ZK1OrcTw+3sRb8xNx0rbY1TcxgldDZQEnOy+RNI
LZpAzMzo760EiIoWMeDvGROiPy8Z5eopZrZMmS2nm4Ho1aGJWdF5FIWYjfD1PFOx
JIbZ8PJHP9VFcGYDMEobRwSs5oUrILNdrBNTYzBSbUroD50yN80ODvQGO9thFJke
mPNKQLocxOMd3dGr/rMk4jLN5Dx7D5z35qnmXUNLKlxTWox3VW8+SehPQARAFqKI
US2mFVPF390seujI8xFJ5CQl2tOPDuZAJRlVvXVkUhIYmnZbjJxR/gPYvByp0M/r
11aR5dPkYT5RUWaOi5c1ie+B1EfHlR1Fav1c0rfuThg8pSfbnLWRa/uES00iQQAQ
jQMakkNOrj+O2Z6JGaqWPEfLKiMtxRyZn3/jveu3I61ksYCOkX/EuTt2ge6WFVuj
QMs87VGP7xoGBeNMRzDjUrmycHPmEVKxwqfWVqCg51na9gVE2zGWTfE4kBkTF/8m
lUeRtHfEPKjRU2IgXToyA8ejiwosa5d2FJHGAuMhiirKbgilf/k7Zsl+wZPLV0JZ
lg15gLHI1CljUQmSQbRnM0Zi23/Xu/f76fSnUZ0eZ7fSyUPVVGn71YbmIBpsktql
Vnikhpb7hvjquE30VisXsBNBrLQx6T80R9UrcN47CEwCR94s5rfF0WYzey5N+d7d
4ioqdZNNrJJEHmc/stbezKsUsBCEP+BuOO2Tn3n2YI5UXQhejC6IWsn1WU56vvEf
YhW7iv6SFzZacaGv6FRB+NIg+RqtmBTWYuVCO6duJHSr4kN3/gFd8ZA/IJSrA3d/
dJ/BaqAIbpy8h4ZWA1aAEeKS7Z/VlLFtmjxJFPK6+OSWt8HoT4paJCAjjyvgfBOX
+QmZSnBtEyi8L82nj0Kw6tveWmGucplHzK9p8myiwP6s2hliaL8F67jtHEnhgXCN
NkvZvZM1oaze+dVFKmxMGZWL+/Ygj+oQoDB6Bqtmawm+N7DxQ7DRd9SOem/PuZ56
cpm4irLJ8PTDH4S0z/LnjXG5mw8L2itVWnvs1nz2LZu4O8wLpoUFUHcO1nnuMh2a
ffQxhtA4dpMOKkj90RKoN/elsLiore1hosdP+ELk73gILDClt5cLqnKAYV8LE9va
EGxTPIUtiR4K3pl98VidGIfh21ajeKCJNW8ec0UMoDkPdAxTiApMzLcI4T2KGxsg
z3Lfs6+KKd4z4C2Pr1yphJEi6SPMCqyiX30UheWlc1LL7Tu+Iaona4TDQ4jTIroE
F8XbjLlz+vFWffmNNSOHw8eyAclOuLbM00waPLeWzsJCPfm4NiCOMFt7nPWwFZly
VXlQytYQ/Nyiqyu903nUh6CsXCDhlpqF55rTPSSLmQQeyBRFW1XuOgDdMK0KG1//
t3VVMYAPCMtKxm9vFUlg2Fq0zEYS2Lwt+hCAeaz0Zi9FgbbjUI940eas4itn54Uz
JLkjByz6QTWWzH6VzOKD1fdKKKpFNvHdOjIJrfQwkrVHvx3mck4EnHeBoioy5gGk
kED7jw9ldvR32zxJjLcmhu/RyVuOwqsR7cYrSSSPhjrV5gUuVyPzIsQ7nA44KPlB
+Lz5N+5jQ/Cde2+CHp9OVw8XszWCNBF0FuVxIVgEvG70qrNY2RQtgHEQXHRagA9G
IghJ65w7C68rA8dhXmoDz5bBFt/y8kl7wyV0a3bXcGwyR5mgZWhS5axuq0ze/X8t
NWm9TCWpasC12SyYg6fe0zzRxNAWMVmBA/qM+apCqwsz6KuvwNfkMPcs+MC3O7xm
c7soGymzQEG1Z6Ei0KwqCdGmDsLbU9I7aEbhwe+KAkfioIx86T4iWiMbgp9yEnSm
qdyuPwlmAPHNUghVnxgDmvVUw+KoUuOq7r39rm79u3vv94Qa9Rjw2hElHnL2bS1+
PAoYv2BDx5zUcIwp0V6xr1Ri3l6Uinns4pharPqspHiGymX8DQb45ytf6xBESOt+
OJALB2Hx+os7Rj0tPH8w2crdEjMn9KnzMRtXHWoc09Y4tIFvZXDW2mOouF7BV3cZ
QcjMMkeLA3B+rUbPlWz1oBJLy+ewwLfBL+lPme/+b3k8HfMMVkg/H8D4F+gA4toR
BszKGpSgST6JeSejGryOU5LGuTHh3+gGZWJYAJF5kAxicH/ug6hlaHDY7HjqCw31
VAoUzFIQuynmAA/SQfeEuVRNA/4zMq2/uVxjXl1w6al1bLVUlHrKzG1JQ8A08pjc
KEFuZvbXcwdm2EjmmKbo9JkHlxk45QL6HZaZusTRHMPQA39bMQ7VhCuILXBhd6Eg
MLKybRV9L0eZ+slg8DbouZwgCtrWC6cN4hKDDFIR5A2YvdHkZIeYWUxtIPJNQZNO
RwQ5UqmKmrf4qdS+t/qPZ13DB7TJjQCTmZfdkJN7H0t6aA15MzREnTJ9DoimqQdl
FKbrqjKvsBtUQciVTWtEv7mPCHsC5S5xKsywbwiDkz7kfjkLIprPiLPXdO+eeTdX
jfb4Q66Aq6KaTN00Pewo5ihPx4y6PLzynpOiRja7cK/x0K6gTMsWhTbDYiy+U/tT
CXfn9ifvUW0p06sVnl96qPw8kXfB3IsQx11BxSrJvMXSCtfwy0VsqybyrFZtxpG0
GUs8m+lmHsrJ4kB61UGGgOxhAcULZZvIfw2hDmLG2O4C/Z8E3NbL3D0UFvgSgjv/
PalljoVRCf28/bWgSKWU/PJ3ZrE5FBdqlKfEdUsXXaq54uE66G0uRdlBPmnA5tdu
Y7fm6Qk+WiFsGNZzgRQPmDbyEBElAfZV3oGNzPM3AxiWt7iZ/YRTEoQAAA4SdAZa
2DHBmYVU9Fnku9YlxEk3/4+WVlds04Bjjaf8FG9Z8eruwDAvbcZcyl7rkAae+0DY
w+mAqKXNu++q6d2VviQTH/8zGFh8iGt7PnS6pAleRzCKxhXAxKXEyP7SbVKPkruH
sbmjTW8ku5jZ76cbIEb7XSbz+N6cCuJ+rVu+x3fR5ues7Uvu9Sw6RusnpayinA/z
0FfhQZvJuU5b61AeV5UWezabyuBUOcdmn443Wwyl9ybj6Ucve7B8SFv6jNCUiY+w
Beoeu1e3MLxrYuMErs0rQ/dICdcIG0Bx8x0kb30rNVD3kfTOn1nlXWjUQYbpZTEv
PndZ7UGVFwa0NTXf+QHq0HttwQHKC4nzPSOvfGyDwXJAZL5D2urbuZbtyeweKLZj
hFwRP1Y70lVKrLnpxQiVZx4byQ+RYeFlzbRsAvhQWjlhd21dCUIuAzBeDafV4lNV
nP87o+YwGOnTFiBLwDr7m81sEqVyQiaH3PISw3cEdi8/CSCyGsta/wUE6WGnhjGN
EdAAQIhCY2l+4ohEFj2QpesV8uGjWzhPRWYMjqS/WXLhgIIyvDtpJ3pmz5SgY4cE
OTVIyjmWtXMJCFpAC779J8+tRpnuh13tJNRCvoVWKeXWcUcMMsnFYomXR9hW6G+N
12QloiCKtP7NMjc7WNm9xmaCZDFf7SYmHKOHuR+hRpA=
//pragma protect end_data_block
//pragma protect digest_block
vRI9UKiSROqR8q3DTR7FEatKmPk=
//pragma protect end_digest_block
//pragma protect end_protected
