// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H=9MZ6^ ;;%EOWT-F\;TOUG^MO'KELB*F:BNWMK1*Z,1^_OP7Z*/%1P  
HOG"A,TAPH]H#GB,-)%82I,PAVLZ>^5!DD8&2P_T#T7YSR!2FX;X7/P  
H2Z^4 =(#926_R"@]:$1!=$ROG>$O3J]WO&K1T=@/06W79#"@_@D?/@  
HOE\QE#Q 'TJ>KBMW^YW5HA5<T8296GA9TV5C:X]=N%L76R,Z]P@_/   
HZ+8:3<.%G%4%Q[U.2[_GE3TYZ/2W$);\ZU!8*YF$MD729UX%*S]]+P  
`pragma protect encoding=(enctype="uuencode",bytes=8672        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@[U1Y[0^2EAB'1YP11"N%Z**,O]L.HE5<0QP8C?:8BED 
@(Z UG0(N4Q<H;!IPGKXTRO0GT[/ATA_!**D#8;@V<R< 
@@&KA<IE@S/,Q1)!G5(DT,/IZ?=_4K^R-0-&%$:O-+0\ 
@@)CO("BQ5.<_76P4<XM*GN<*/Y,W4CDN=%EEK ]>_$X 
@PWD/SE4X\CQN*08BBK4?LM5,-__59;:JTPO[U?8TRD$ 
@\(ZGE?42<:?[(KBA4:CM6FUPWNC5KH?7RFV(@XV"AK< 
@QZ-H*GD5!5$E?IR>])O"*RL6NN *R2+21#55GV L?-\ 
@-G$E8O&*.XW<W'5-Y'ICVES6.9$PRB^UQ#OL-A[9TK8 
@W)@%\.9)35;/[@.SV?N[>E#\V(O2X_?CLXUF+0@KWT8 
@RA'T-AE<YKET)0UV(-IBDERJIOU]?+K^ 6NO,*6&TR\ 
@ @/ZH4S9ZKAU0G)?*NHOS_4,L?/2KPU^+SR\)!JW%VX 
@#I7RL-Z-;\=/V 1'_>E <)A,1O_,9FU[UCAH"FA-LJ, 
@ -$Q.3*9#5XC.M5O%%K+!>E*UEOGUDA4U!T.%!S]RY0 
@]WR&$3.5M8PXNL6Q4.[ 2PHWOT$_70L?\)(!(87/XX\ 
@!V4F;,@SKG8O%]/54Q05P=N9>'V:AUO>;)H!0DQXV,0 
@O@VLY&EXO01$9WGL<0E*!NW!U:SA8*[K+'\]:#A!9'@ 
@\T3AUE7P7R"5\%DHF/[>>]D:(*>?26JFE&<]CGO(; \ 
@(P7K4^3S0JAB(5.Q(-FP>==TYWKLA0A97&%T1 7;QKT 
@#23@&8RD)&P(E[\>LNV5:]7O P?EX!HZL\^XEN.A9+0 
@;&M(/>+PS6,=0E$>MKRE!==2P/M18V<;,7#%_*5;4U8 
@%W@-@,XFB.L8N&4%.* ^8+;:YL2!<K)-&%G+J5U#'1L 
@X[=]'RV*F$I$(K @A;=O9?%",[I85%H2>\%&#+83I&T 
@$^2^@GARG?CLKT)RYVUHUK36SVI1Z;#LWF+A]Z1DN-D 
@H,:)<1L4D^DT"!T-6NJA_XRP+NWO^$_<>2/RZ1\4X0P 
@/,VP+SYX?R3./TS, &VR&@<OFHF8'K6A^(>WV9F:/I( 
@68GAW-R5E[-(=@ED6EFBZ,%$U:W+&OOZ=[%:,B%,?_, 
@! =3^L8K6FW&R' >KOSX#3PM4C?^VX#KW;Q6L @L#'( 
@[WB92O09*6Q)Y4ZZ_?IPFOKF#TS/M9D"+KJ=(+.>&<, 
@%TGE\DU9/=61K>0VF/\L9 A*\ S9X>UH=N&ORLG!D4L 
@$*E2$Q:\W4U#Q)'*X9/4+4.7_%-:+;CLM"[UYX)U1X@ 
@@X *(X'OT,<X^N :N=(M<YDK.$KK4(9"KJ>XX4C>^\4 
@RLAE1G,2NR!$0%:?IPE@$Z9\!WOZ.K^BE=4QWV&\&QD 
@D;:' 7]*(C>/-9L^7@C;R!)UL9BW>BH!M\)4,-IAG<L 
@T2<KLOKPJM4*U=7B'GX_45I6'RESM[(>F6XG4?A15M< 
@NUS?UOC_;=*5W922433"GV8I^X=ZR:R!Y+U+OB0 _O@ 
@1V?/]QP!7_?N5#OD_F@CY!2_%2XJ388M96N&0(1Q8JT 
@Z(@<FO#?L@_$JV!8Z9JI:3/Z.'NTAS>=Y3XKXTUD9J( 
@6@[G"0.3\^&3VG,MRLYA%#ET MUTU4Q)SA/FV@GV-,P 
@73E48B6DON 0K 5W^@I#+@+I1.,X2RRB?,1#"4,ZN^8 
@ :J?_.5,KP]R<6S,196=*V]N,"(\C/6]!-BIC>G-S*P 
@(Y$!-W8DUAR]SNZ3Z93%@^0K*&0%KWA5=&*$(]Y=BZ, 
@V-LYL'SL(5D^"V'&Z1K+)C*O\^FV1-1F#>)-&.]EZ1T 
@@XB+!_T=\U=-&]QZ6-N7__Y/<#P%WF*-V<M87+_4 4( 
@CAG89_CH)NU%E@>R9Z/LZ6'$7A+'TYF7$,)'D]O/?-\ 
@;WILR%;9S9A0#ZY(3*!3]"5RRM6?D2/R]ORK-N1#6F8 
@LY>H@;K?A"M(YX9YT)7C4:5N "0HL3F^VGK%N,E# [@ 
@NC:6SB.#&A."@^^GG+G@[C:I^14^4$2X_106*Y_149T 
@@1N>R6;=@46PIH#2T,+UX9/R4SVY0 8"<1=H?&-C3_$ 
@0'GM)>R<XF\+A4CNVXSW\A_W"@8L;W[*K>!N<@ 6P%H 
@W'=FNGK<H+=82/?-?FO(&8-XGM,WPZ)HU<X% %#]_U4 
@ZI,8OZTF,(630^4+HD-FW'+6HJD@77J4/)ONCNRP/ \ 
@1O'2@F>$)]*OS.8J?KBW=!8X!LD H7(70X1F%H=/N+X 
@N;XA,N<K-;0DL46L]>%" 4P>8!A/E/H=<#V6RUL>8T  
@CCY4,LJMJ"7G+[<DD,ZAQ\;O2_GA;8:P'BCJ!0):IVH 
@N/.*:.@A MSG*H>OR2S@([:K(Q5_A!?@.>X*!@Z<$'8 
@_"8.WO1<3KQ9]]Y4>1B=4:4_AJ$ S;'S!D/5_W2PY!$ 
@Y(0='"+%%^>-OE$0;J"D4 'KPB71^]CX \5B9;3&^6L 
@8[34>Z]\'#>TU'MB]QX?\*O#23X'Y->AH\,R-3"CO$  
@';%6;K;</QDL2"ZXUP5.,ZI!'K0TG'0@Y#.XS+8P2=0 
@&541]##^*P'*S5['7=1N[$V*3[@[2?:Y"V;U)MB8-P, 
@ ?\MV:ZG+.P_!J"2NCDL2]R_J -Y$/]Q1!J+3!0-M%$ 
@38O./ZO6#)1NWF56TI#87 E@Y^H2$'_0KGR[3=/U+4\ 
@BQ6+#V<P/=C\<[<Z8WI+U9CYJV8<.CE%*]ZNGYPL]6D 
@\\@08Y*Z=*((M4FNW];N]G#:R> _THXNR+$!:HXY/R$ 
@N,[3!.I?RV\H]'XL?\WYSREU)P1\*VN'K>$&XD%>C)( 
@6H"HDS.L(XQ6@LDQE0J&L'CT?-&_)1I/KJ-;W,QCZ6D 
@6TKAAJ9@L>X/R6M+RO%OTP>&!1U9.X34R6Q)"5#JB!H 
@0QX#-,*\.>O@8&!Y?1JVXB"A(?(;VQH]00JP9XI7>9  
@#L*KWJ%<U%1BF_F/Z'QU_N3,\U; ?S-U_JR?:HF@=>L 
@ _3TC1.36.BST@N#*!O-3,609#U?[9@?NF72 2ZEXY\ 
@D< 8\!FM3M\J%Y=UC_EK9\(O'2P9Z@UI%2)R]N_C0$  
@C(L,(Y[3<!)8Y/UDK'DT =>1%"DVV*@:]=<K>X!HEF$ 
@5B0;2VO.S!P9##'$4>GRYHW\(9Y++,H$K<!^FJI[:8X 
@N N[;W(;X_R7!U&?XY&Q#4Q*!',=W9,)@GT[Y,*"K/X 
@?GGXX)C3'&L1BZ +#'TFV-CEA$^P2FZPGJ7CL0=%3D( 
@$N[3Y[3Z0"CB<(D9/^'X,R;I@@(@T0@^N?*8D O_U.$ 
@F571H%SJAQXX7"JI\,],J$I$6G%T8(_T"Z@KI,L& R\ 
@3:Y,$H_OI0=2/PNU6@S(<]@0J0;0' ,%.7XDLRO6V(T 
@>HQI!9]2BZ<);:?ME-+/8IQ&BH'-CA9D,=28L@C/=)< 
@9QB[;[,F41JVXT?.]1H36Y'HY%G\(UKIG.RB<*J!.=0 
@P(U*AQ1C"\3L>U/D;&!P+(Y<O>?9ZOS5I*=5R QH!8$ 
@3.[=PP(UGGG\62!?<&13_WCY.44ZO%L7T[(425#LH5L 
@"V6:[P+G;>O+%=H/R6^E]&T-DF4(2G?."AAOHV&DPLH 
@B:NAABHJQL!:GRW##,B6B!2)3NT&PL7R!7H'CY7W[?0 
@?7VH@O9DO%34W!%M4>CNZ(Y^]00.S\T\;8/%E74FN2H 
@>=#RH&/OB#VT]P=.@)H"RG9PR\DX4C?^4?(7<K?NNL( 
@OWZIX#HU*>,3/NJMW5U+]"W+"U'F"!^VI611K/IS@<0 
@G:Z.#?I K'3'9*>WAJ=WCVI=PB4??59:/FB:3DT,V=D 
@*P)E@OR=)-_'+*P-#+'E6T/ZGAVUC",W)H4[1+K^R,8 
@C,H!#X'[Z?;%<X'6$8&I*A"44P>M_B#.O@/>_A!]$Z@ 
@/PDO43@W@<_:/VZO35.^ +EH^2!,]/!4I/'(VI>N>VX 
@J/J+X_=BRQCN'+G"I(8Y@L9K->VV6?M[%,N-GMBS-4X 
@(0OR'XY\2311KR;YS8&&' $C$LC6J#-AL-->)<2^' H 
@<K'J5TT-,#VS#N0_Q03^-8,T%H>Z2)RWXP:4(JJV2/H 
@$6H%Y_;)_[%>UX+5,\+Y419;9&%ID\1'L-3]%QCM]4H 
@U?")A!*+25L]?+.J9Z6^'E/P?1,<4L:H=]SSEGOI.X0 
@HRM7DS]<\NUO_.EJO>5HYL4,YTP@L>E()/R2OF?.&G8 
@R#71?JFN=]/P6B)]GF5U;48TU*W2,:FK!G!C+&S4=DL 
@3)E_7G?PA50]<5:!+<_R)J!7)C"A_-RKZ\'Z2 5M7EX 
@([Q@>R#N,G5<U:@I^ZN.W:-=[,"#A.IT<IZNN1A_RM\ 
@*3?!0=W'43"LF;F=HJD_ <^XU9]U+QZ6Y,^ETC*0$;X 
@'1ER5"$,Z3QI#XA$E_M?YNK9<8>'*?=F"69 6"?Y6R  
@6QR\4D,<G[8G*?JBY!6)W/[[=K!WON TWXWSIXF:7M, 
@K0)Z(>;LY%K.%PF"P.VHF1EM;^89,7@ A&UU$VIVI$< 
@)RP&7?U?K V\)D-@K;_(6NRH :H=C,XDU3@I/ZBX@I0 
@_QRMU3FCQGFT$(!^JL 6'C#$VN#;Y!^-T-XX%6)_N[( 
@LUH0^M]4+RZD^-?]\P%9?"R DSO["*9B"!]E)H).GST 
@4/9H92>&U"VG/[120#C6#I%[+;DT<3 4QB::8O2(DS4 
@!2&YC)SU.&0*F'R?2]^H$.XU@I<4;YP>'NY)>TPE*P@ 
@MP%_S0>5P>3#I9^;QS?+R;H8/4[[6A326I P[HW$G4@ 
@SIR:9UN&EI$5X72:(U1IJ)<S=)6^5-_\DD=_P 0B=_  
@DIY3)7:_Q.9"4?.8H\W= X%/5\,(2ZT;,!MF-^65F<, 
@(#7]C(X<KUY"2&?W-)BE$(+]9D<(W>UN6 F$6O7@QQ8 
@1B63 B=KRE@5RQ65GJWH&3/X EO5=HD5*:!,D:_-<A\ 
@S0B:((N3/K[\I+KP_Q%(\XRWWT*^JO#FGW3[2@ -'M4 
@?Z2- /T)DUB$B> ^HMQL&V9_\<T4+GX.P2_\]3X'9"@ 
@R6EKO8*UQ>-30()F+TXSAUP^%>5ZF>4+BHYA0Q](!PD 
@IY+- J_>]) @X%!:<\F"*FU//XN'&..$FT+1KNEYXQX 
@MN"HD-F^G? +S"6VG=,X8QZ&$I_Q97[?;[2&J]?H+^< 
@^1YC-WDJ,E'Z"# +<3=B^YPXK&-NIU#GNLO^RKW[/$H 
@$QYK)5]Z1-[A.3+AMD2/Z5']A'"<)_>$*:*YX;4:FGP 
@J< @C0J[Z$WM]$06N[#IJ7Z890)T_G"-U2?&H;@+N9P 
@D>:Q)JKQ&*,3^?/$?*VO[)F[54\?62GAZ^U=>\$-Y^  
@"U">!EWY.R:YAUL##V=8!:#E?LW4^&4*S]#4&5;<B_P 
@@W9(.60]Y8\VI"4CR!=_7\2N"YK'!6Z'>L*Z=I%2 KT 
@;_?>W@%_9%M7H?<E ,N%?S5_9,ZY4!PHH7?.N*1SQ#( 
@GE FHT0@T5,=,V%,$;.B2P.;MD4G:A5W%*,HH 2%@ T 
@,8?YB,&B5^=%)R4OVVZ(BPS3$\ZJC\_4CI@BR70LR1H 
@H;(%G4B0LF(V^M9,+(X*OQX'95/#2RCB-8ZG7Q44;=T 
@[GG[95BMV_?>X5$,Q!-R"BV1IHW: $1<!7J(QA8'T"< 
@8F8=IRYR_G!V;@?&JR"2+^R<@SK]]Z%JN5^ -$;9SR< 
@V&\H[RF!@FW]5""N<4Y@%3'QX(1.R+=4]O8<$ ':$_T 
@3,0$-L3^5L\;F?3[X.3>T=?"Q G0"K: 1&4C3*S ''X 
@D#2P40.*-JD!H?!_&\>Q-Q4'J+[T.V"]7 ,9%%_%NRH 
@]C=PGD0 R8LP*MD5FJ "NQSF!8CO4F',3NXF1"LBB/< 
@S!*Z*]P/N';Y>/<$]D\%Y.2!?I0UAB&_YD%[KP0(WE\ 
@W[38E3BX,->L5>J;@._N8MM[O;IF,_/V(7$ !*AS?$( 
@@&A!G&4N,TDGC?S*0H*-X*;I3_'\0G7#O014@!J':SD 
@29!++&5JX(!YVRSNCRESNG./G90S](2>T:?2PF?89S  
@/$<Q6JZ7):L=>5'E-Y<1/] =Y_HZO'TE@(\0UE2W_"X 
@2N#K?#>TEWNVXE<B6/>-G<KIOSKDZL2B]A)1^_PDZ/P 
@^1R0T&3L[_]![M'QJ8M.)U\Q7_R]V).!\4'HTP5KS48 
@*/3\.1_K=8)4/2=F,[<$L4V?-9!12D#L<633@XR4\:@ 
@ :67KI?Q@&0Q[-N5*ADLONEVE0Q3K/P-<'1;T\N@$Z8 
@ )%8PMB5WL-NC9<#XB8Z..7:N@?;M)_^2I4#FT=S+HH 
@Y>RIHAPJ.37^7WZ%J/0J?N;PB&>N'%>-SAM:3:/F#U( 
@V2&/+UG$?DF<N, ZJV+RI"]Q]E3<*%&B?*/!V$MFJN@ 
@ADG]=RA[^/V[&QBPWQ_WQM\%<2DT=.,)C)WZ4;! ,=< 
@BC8T^F!*6YQW;[](M\&U)8%VR59N4A[/=?5/.(63\[P 
@/\S4 ")W- #P2W0F=+'&78>X7=DZ47@<1\4T2-8U[P4 
@-W!-23S7C,;N&Q@D4 WFT1'JN6C)>:GFI]GS(*LQL9D 
@+:F&CI 3\,8FS1&GGD\X$/+>N>4^/275*OYC6CNPW2L 
@JI@5:U($M$Q$>?Q@RTP-2OUG^[! 8:8H//ZTKF3]8%( 
@_%,Z^\P0E##R[N@PI6*]B?MUN;N4PA!F@F;U%@60N1T 
@"2Y?$UJ> X\PTF0KO\CD#0SILP5"*P<8,7)Q2BT5\"\ 
@BL4Y:-.^&=J+N6)$3FE2X[#BO=W;'R]*=[@"+9-)KZ( 
@&3V8Z"74JO!5'';TFEL-EY"92C_?+:SU<*JZGPY::C< 
@ENMJNX-.&;^=Y4!O7Z-[\_[$Y2&(69#.(\DU[:6&)ED 
@MCDP7Q61UHW@-F",< L"]/>W,':C!ZBB AG^C.@\!OT 
@;]G45UGP-*/')6:WE-Z9["_)$1S2")TC[O,1^;V$"KD 
@COW@"&382L_7>*Y&D;K="#(EHL.7W!STV )KD*[Q_8P 
@MY_?(>%9 ;UK&I+*3X//(/>&G*C/U>HZY<>192AXX!8 
@[10X2\@G?_");:Q03S?S1"[M@C=50J YZD\WJF%$F4  
@JY0->14W?0R-GT^]NGT+WP_N=B,M4B9$6% ]V7']Q-4 
@[+;<GB0"P \)M&Z8RRMD?9-5(RC3"\:!-FSKGU@F$HX 
@TJE#1DKPL8:IFTH&Z9&PZD=7=HX9)(SD\&2Q5:L/FK0 
@X/"<0 'J.%CVV"?+8F5*/BW2=W=43Y3:"4E3\2DSMS\ 
@K:Z<7_$I"+O6BTDB41;@I74"^3^[BZY#L_DR(TJR9YP 
@_9U8"!E_(=2U&NU*1*UF+IX :_$'/V1X2U$\V9[G.>  
@7'U68IG^7_UQ(0)P;#JE-&W4,.Y^P'"N/Y^2+/*_XHD 
@I\4[ORRLMV=&&W=>9=I:3,R#CX>/5MC]H%".IMX;-O$ 
@.CVC7A;.&)X1ZA.?;Z_A4Y_W;WNT3>%'SJV[[".32$P 
@J=8O50P7P^Y[EX@^*1TYQ/0[LZLTX:OLKRN;9S&T)(8 
@F)RZUI*@&'F]L*$OP]L<64O$IYH\!A!WY*+23"(AV8$ 
@6T%CD,Y7&#4)N9ID@.L]^L:^8I+!FJ8[C-RC=)!HT"D 
@ L#-*//V5O78JW"-:-);@T1#-:;=/ 9YN$!1#W7%C7\ 
@ENK_9%-HHU"P#N2#6>I( OFXB@7X88P27"3KRW_]>-0 
@'ME'A;^(V:M4]E;?'"S'6;5',K2(&BA=2^XW06V($#\ 
@5.0V3V*3@*HNN\E+5H5<+I2Z('YJXNVY_:HG(T( 928 
@8R:<I.7KF/%:R['@T((]P*[KHZ=2UHJC1MQ:+8.0=YX 
@:@?Z":0_!7[C%><[99^I@2:=*,!G$N3II%F @\<<?SH 
@:9X0H"[OC :%N'/4ZM=%5-73!#W?:FR'=JFFQOO1,/H 
@1B^L\@.V?^4"/\"U?:.&L61OQ1ACDPNR"/J5'7<5UH4 
@'CNS. "C;)A>3']?#4/*0LR8<].X5'+5[./2^83F1+8 
@[G*E#9@;$?3NVNN%N*OQNZ%GNT@?O99#)75[:^>E+]  
@6A=G/P+TO/>F\*+#$T>BHCE@?0S$JM!.S?;D*3(4F<$ 
@RNRG5@T]"B2E?'#_UOE47#^I_F4T\.F]VA?,]Y=0H(T 
@%KB[QWSV$5;O6P3,[W\!E%\6M*T/JHTU/L(%">MGMY\ 
@V,"0-Q5T:1(R,WG:Q[P\O@IF_PD"A^;0.H4$>YC/'M4 
@SQUCYJ5BK#!UMR^NJBXLT!ZF,KR 7YG1FEKFUO=K*OH 
@8JL;,Q]FMYH;5523QS9Y@C-.>4,92$%CR).!%WN3X[, 
@&G=#N34):M2#_A6#HEQX3:&50JR<I&[LUU95K"\]'$H 
@3-![=F)3YM16L]ALB8]V7+!1,@O<A42BPLFA^A0,$Q8 
@9=#8Q19 \8E&?&\E ,#N.%ZMH3?L<Y%;3.<HP[&!K2@ 
@\O@!\/DMQCUS3%&:C1]2LFFD6PT#"SO>D?^WSVZ/Q+, 
@$@W'2V.K\R7=1KX!'F%@9$X?461LMJZBHIY$Q%'>=$\ 
@)T5=H)4U.YQK&AP3'LDVC><;[E19^K^"4AL;&Z!1<2T 
@VSM159L\^X7AQ341OYW=,WIDNLM:W=7FB_UM7>L9&8H 
@8[F-)8B L'1.DA'XXW.K'15F;_Y+'$.EQ.3!!W^C1V8 
@.04LNBB;-"@XW57<I:;+GDV3R\B>-,KR6IO3:',+7N, 
@WI>LYCI('^G<H5;HS)Q5$Y!9GA- =*GD?5B9GLE3>V$ 
@O6M85%@IT()5F7.R2U4J/(=AIL'X+&R7R5-75'5*0L4 
@?$A"A6^8@)&"R+U,2%K@AO[P01R]C5NOJP>Y/>6]9>8 
@W?KET%.28%?@]O(PPX /:"'?%>3^3*#\R\XB2\I^:L  
@'*"3HMD[33"VW!^:G )Q685E_0^VN@,LU#19NWQ6X>( 
@3 JID!_B[Y3JD':1-C32'5IJ:%B@3W#0AE_2@3V"WB  
@H<CL5=CCW]KPK8\N8\0)'Q!DUV:07$,Q\QH0K!#A7Y$ 
@C,\:CDKA>"\5>>-5_;D(HSN2@Q-_+33 A<R<BZ=DM]< 
@)%.$^'5NT^@(H8OOH&4>@_ HE%;<@<*N40^)'0Q(A[D 
@1^/)%T%)6.Z?<=BG$G$AUA7 QP[R4YDVK7E[>SR\P>T 
@JQRIDOIC9S8-A1#TRF\IR1ALIA*942FSWY":$>J@UQP 
@3D]'#+L]Z1[?S"8$<'N >22',U CJJ4'S0P_\QHB #( 
@C5/58^MO:N]*\95WMW>0TLJTECURL(QVYOD'K-[[UWL 
@!Z ;8!@8NL?%UQ/C(LD.XY,,E4U'GZ><<(IVDB\"TCD 
@J&VDZZW>IN*1Q<_-DR^C/GXGQ.!*#,MSOPI@&:&I77$ 
@]R^=R2(-TS0%PK4[>8 B2*7HPKI>](]34UZ :;-7578 
@R=DCD+=?!/274/1_8 X;"I>7@,6$?:9&]A=QZ-A.B[< 
@B63 6R-DY !8C\LW:CGQZ![)T"0@?CC"[4=+Q><..4  
@1.Y;TBH<Z"R*MX'M0@7R>5],D9R!'^%XKK*5V)?%(X, 
@,$C=A'E<$O]-!$1)^^5FKL$[1D3Z;PRB<]$SP?) YS( 
@0V%CVK4;@3F0^J*1$P"$7A[<")?3,.X/,K7<J)3;9%@ 
@0PX3D:5S!EGI;WF[Q53QU&[=D[6&X R?L)CE9]N!MS, 
@3(W);\BNA0QGH.RR&DR#GU*J5K6]D0N6TS^%XBA8V_$ 
@[FJSR%*9GAK/ Q,8R[+1\+P83%\"D>H1I0V-$'ULXR4 
@I@YI@AH6QZ4B!F6+#Q&:T^'$PPXEKO(LN^9TQ8FU0O@ 
@C6"-J(OO5%;&5^VU[L8'G"_<R2*DCTY)'%@5F",%D/( 
@!Y?EQR0LL<\N="7S2(&&5,LR:B@(1IEHQQAT\PLJK#0 
@-KV?3!.X_NG^UL$BRO5W:0%1<^P,K^DH2M+A;0VH,X4 
@0U<K2@&!'\CV+,/$(+1__@4>!,5#=UT0+U4,_)_J\1  
@Q^Z%\KVL"!%^4=;\VX*->3X]1/HHAXOOIZBZ7L0S<V@ 
@2G\1-KU?S^S6YHBLW ,PM!/13X>6A,$NF_A7.+M2!@0 
@^W>0UAK\*>:41RKZ+F?47O*+WIIDCN9&;)TMC#[9RZ( 
@\^9L]"7,SFA! WN[JY?;AE04=,5[RX(\2UZ0;L<F1P@ 
@CG#P9,1>J::EY(9= +35+Y^:=IBH]'WWJ"V$65NQ\M8 
@;-90T3&[O@>\VM34[1]).#V<V6':91_8$H9O/3GJAL( 
@8<N6Z;^#*[#\P+^_:G4J]D*C'PY/XV/7L@U-.T'!\+4 
@/S?Y<VG>5./=N5;>\;5 PU/688<E^YU;9Z)^T.0/6>\ 
@NS81^"=+="LUK"-\6JOPJPHYUE'DYJ4G:7UK($A^#Z@ 
@]#][<!2(H%_D*BG;63=. &.>P(4R]I<QD\R@)"'46#4 
@C,"UV'ACN8(P^T$9)XCV,V&'W[+J*5C/N"P\DN</D$H 
@;OSGJ#N9_;];@PO"#NU23I&?.Z<I?I%>CY ZF>_*O6P 
@N+E[V+U?]8.N+*#FQ5D'I'7=ON/\,Y:\(TDXL+.#U]$ 
@!R;^EV0ZDQ$L?9-RRD]!,;P.8^6:FFKUMXS*PX,?34T 
@C! Y18ZE_+/DD55O#FLI%-I/00^59?XY]UKVDE5]UZ< 
@HG"@+X2_5N:FLN?CLH;=A@FO4O.Y04HEP_SP=8-_A$4 
@=0C78<#P>!U_-65;^LDD(I'K;9:^C=##G(Z_BWU7+A@ 
@]+[>_$5&*AS13]*>+@#F-9KI<I)AR&4'._3=A8P2H;H 
@ONX)(]GI>ZH&@ 0DXX,8XB]+H7\(Z.@^EP[6& J6&-8 
@)062B_B0E+W0U\=>%O]A0IQ@\\<7>N12ES"LF*ES.+L 
@9A=-.A!(S42(ZV.BE*)(#HI3N_$(M XC8=0)I%<GP < 
@/A0;9=L!2>P^T@94=M4!Z/\*8D/'=]F$$6U.Q).YD D 
@P&TD3./K)#!]2[6X /JUKDAC.JIX8^KSKZT 2:.)A]T 
@L_!J&8XA06^_W[FN>'99/\!+JFMZ-!8* 2E3+\46;U@ 
@ZH&_QS=A<P(M^,(\OZI(\@D*+8X5>76CW(\X&3V,U8@ 
@'?FO1*N2T;)<ODV2#1<_<C+^=-GH 37(3^EA.>]/\"@ 
@/?P%;##1;=SL"[^5::V]7W]923=KI^#CE6_9@98^-?P 
@+I0OO3C_2LIVT.,$&A$NF;SR #]#].?GY>I.@]Z/#*< 
@H%.>'@=KHM@],TC 7$VNY8=LB[MDMJ^9PEL25TTFB_$ 
@/;- ZZ2 =$@CJV#RYE/__R.UVH2S5Y5O0/BE?9>X,E@ 
@F:#\1,QHI%CI+%;^0'6(4DVL]%CLH!=GZY:<:2(F"$P 
@+@7X&=(. ^ZZ]+R8T^R!;GJX/;=K;+5&HI-6YJWL(@L 
@! ?X)B4R>+:T-%^AEU*KGZD3\UHLD[(7)*ZX!K=H(.$ 
@A&0LCCB$B8P@<J,T*TWQT/%O D7(#':-=\%&8OF@@40 
@*M!>N8:7;<68%8%_T5-;MAUFI91"4EO+D8+K\OG!&S4 
@!>H9MEK"/R(_0J'?S5?1, IG*NZM)YE'5?"3%,V0IYH 
@W^"'L><S3G!<I)JED7^T7 $T<+3$5.#,_,D.I5E]^0D 
@ 0$?<% AT*[UV^JD84:2 #\>:N#IB_M\7=G39%5_=L, 
@CGV JPUZ'E@$J/<\]. <WG.!E9YK45MVO3B#0PI-GH$ 
@&$N\?TL HNRJ.L@LLY5-/(C"]T:.E5'CTR&78%IDES$ 
@!:;E-M6L"Q$._G5%#F#O[EA;TK/1Z+.*(A:;LH9U^8P 
0];U^4*W34UWG\WE@K:^ ;0  
0&X17+/@*3B1>HOO*J,[3=   
`pragma protect end_protected
