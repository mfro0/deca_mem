// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 05:48:06 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gxb7yUVE44uOVJuLJ5JIHNFnwwOKOEeBfCWRLDmYB4f7BUD+z/weTQFe+wxECqfO
YgnPSGotWg6768dvOC/Uq5Fes39F7Fljxhfbvd1qC4k3LG3aRnZz0pikDjItRY6L
2eLhxWHCQNihVGAg00gYTTd+O2yEu2TRBBGHNuHDoh8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31440)
NoMkLwADcfIveHjMl4qHAqooWPXf/mC4LI+6WoK7+j4+boPuIl/M4TVKNx0H4Cte
wNx5aaeab4fMCnQrm3lW18CHFP1mfzEbhrv2qqWW4mt1b5s6iHLL/Scz+Talq2aR
j9EkixfHbbJmZ8OA5uC6ZHAULzV621xYhOWhghbo206TZ/N4CTZsRjzWOHUQ5V3Z
mRII/BjfGoETHfIkhVtpD0n0Sees7uGwLD165ixfaVSF6L9+SUut4kBySvrEMYFf
9EiT9otqhAx/1DyEB4ye6ID4rt+PY1w/0n1Aj7aXftytN43LrUw7uWNFRATdynXo
6yiLftUQeyPro4d0uh6m5q+3rBMWyQ3n7tTjK4KivujEN7QPN22CyCCLVjT/cVaf
vPIPuTDrgKqxpEIKHZjPjpmL1QvEoAdjK4P9pHO9ooLQ4t4nMkpHFNYBf5JJnY6W
tMVyERcFgOnU6RbcfjGHDUDSiWoh3jq0PUJaxc1y1VK9UrIIVPTwQl8A/t+mT7Nm
D62ZkyPlmB93BSiwwHT14wNPJe59wyVK4mQCGOcU8xokehJ539zpYWCih+Q/4dHh
4jqYUpiuYwpK5AOQQyRDzL8x2lhGz6md+dHZhtGtuDauYJC5ZbSDJvfC0LtCpu4J
jqtksKUAO5kRtUBGzVH7kWT1gGeeNMF7K+jbT4eXjxF8NiiQ1j1rRzTIQVPyoud1
iBdbrzMzDemt0HsamViWEdoDhNUfp8p9iCMigijzAiIZR/8fGRqRsDSmNSV8o9wY
Os09H9gO3z1dgYi1B8Qprz1WWO7EPPfarVX6wAM5qGNEpe/zT3oeXBW52d/reNTK
peNzq+nlrTC9fDcTtFXpB17H9EbWFzFFr27xDI8WNLt3d7XlluCJ35XITr7v5yxA
0coR+w6F/I9kgTN24xTWifPRFXmnELTUIWMTESvk3XKlmU+fniapD2v9p3UwP0Mf
czBDpKOussuBX4DDmnJMFUGTiU46rNsejxTPl3RJ7CG1HfDTHASDjnldZm8AVAX3
/OfdhaMVt0Rm5Af3lx2TLCgmybIdA9rXE1Q5KlVK9nIXYPRwlflJ5M+oxnHbay6b
0Ck5IO5lkPJEVxnPp73l0OMgq9KEC0zFDgfHmx3U+MwefzTGmGhc9nKfDzGf0pWE
touvRXGwJXRCuuqbnJ7Xe7kKKU8cX2HEza4Y6aoDugwSn3GQIoLCsRU+iM4pKNCu
FgaimuJykTdGApmV3oj0G6sAF8i1GmRXHyzWrjd4wYk3NgaoROrsnsrMimcP4Lp5
RQTBLpXKEFFErDo1yLj5Jr4BkrM1X8IL48R0G8o/BFThnQEMU4HEjmC6g8X+5ylI
vtmn0TfDbBrchztLp79C1DKCXpwGvSmQFcs2YgzKAg5brsbo+sQUZ8MQPSuHVsGh
dyKrLRvJv+Ct/0tV1uWF8YheeC33uHvW+MdClROqI6+OyREwPW99h+jW5ZBKpz3V
sDIPg2FF3TyiMNZAYCemHUHJcQSXU50yQ42LYmQrtws40fwzyEThRTh6uPVDztFb
tEt3msgofddEHNzhJiFDZerDoMxqsIaFfHh/e/rOFiYtBu8f4t0SNoob0XvC17sM
pwvSOzqhvqd6W6FzO6SMzAuJ6dOKPATriVmvR1wTGZACxUIqBu9QIe0c3CAv2YjI
dASsdpMLcKD0ElLlSzVBlgX7+ASzmmL/72kaR5qEDQkNf+6rjf0J99rmj91yYaVm
wZUzEYWFOoYa1Sk3/d5EiwxNtz2HYmmU5U2ndjBX8HS5HXdQrwTBJvN9aaMFUHrc
waLRVOZQsElFR9XbQd3IqtESrQEEYApkjtzyHhP2dfaxOeVhmOoedmBUB8LkgRfW
fWj8wZ0ycLG4jnAKiJfQj7n24NN+GeeW5bfRGbF5QHTPGmwTGxzNc7vmjud5MX/b
eYzfkpD3T95021AB5FMCbjDBTQ47g4yvQ5+0fQOjHIBUB5Km5pSP01KIfYh44fBm
4meFN94tVsv6vF8Vh5sk7AH1tN8fjKKofqreDfNVd1+Dp9UtQc+Z6OSEFyNVuUHc
n5mpXvPa45ZQ7z54pYH1LJWKopkft/G6Bz1REmfNvTiUmFsTg/YjFgbes9KKF98U
Kvx9zb1W6C6KEiWrnr1nsDejO146Vc9unxBsnv41wElSvkk/H8voNTmXaHpSGOpU
w1dxC4TePUffRAaAmSdFB4inxBDkkjfuKb4rFX1RzWtbihLWfG6N4nt4m0Eo9yGm
7MIjoDW3147HAxk59Qomw27mG1Cz/xX9qMPU2NATJ5XzAVHWYmdznqG4gAVs2lcG
HBC2LsyqK2wW2L9+K/AIxc77P4KEcKjUk0sc3WJuhVnc1rAPoqFVZi7Kbk18MlEK
CEYvQexuRhsiv5ipM2kCGBhEviNRzRME9L1ndgjMqGSmHW5Ra318tXpaQkCFGBlQ
XZWwhKZm5f65gRwYxydCTyV7/e7d5cS9AisCvwTMsAfcxQnOHSXVQw9zUKljaBtw
/qaml5q3LgzbzOQO3/OZHQhu5hPdnwYVOd95MsBkMwc2toLKQ6Crtz1/8jSUlWju
FyYC8zxRXZ5Qxur1JBHJ65kKxMkfaVZBkwqpko9UYsqBi1vENOaIrJYouDK5HA8n
YK8Nh9+4466lUpdJ1OSUWkqoNdoPu88hUmvNcyrFok1KWheF7zqGT+SSNwR3Vb0m
GcDh7pJLW2/oGSQOoKbL2jvJ1xlg2Onp5DHIoX3lBtiYBdeVggaToCZrB6hreUzv
fLs+b/jbW0+sFreIROK8qMWxyls8qGIW+CPU6alXVmIgKRHmSq6Ca+E5UBPH7IPS
tibTol9hVKN9XUJTfPjwmkGQvlVH8HizL4mJK61lue+hqfeUk2LTb986FkKTFRcO
ZUpFW+g9jTWEoMsSdqiMcGc/FhIEE7G8iqUBBddWhwmFWt8FRD/pT29pbVxJke5U
QTWaGdQPiNkks3rz45iBRq908OsXlb1BbCnb8FYwjKY7E4850e/xcVY/5OwoC/Zq
2e74FczZ07zpAdqDiQUedRP5O3xOR+nV3g8T9ZsVAdHKq55twkr1sZHwmS20cx+h
J6tlhL5VNZHKGByEea8CuIrlUWED8woNO2AZ3PgFic692XIvPUtNPQXD4UzezSL8
nRqzNfS2v1tBV6tmWIikFpEpI65GjAFrtx7iQNzei7aQ9UTd6psAGxpPVuEsTPAA
5z1RaP03UhK87JWoroHQT36LpjKzZVoIb6cZnQ6tYlPf6YsTow9xYJxbPq1xpLya
ZGuU1C2gof+5pHLUl+/rmDRkw7mLxmkZvrUlZ4XKZ+Ayo7oEi2xh1itRlENmtPgZ
/qYFesAqQEBpjYtwmcULxA1KEaqD///BwssOau+KX6n/GgU658GjVKQLwBl8Bfwo
DCTuNxQOy669UwRNcwmIfmtgm2Rkp3nxZOo9Y2EheipySZo+9qmSPdvBovzu2IUL
daSDXcMQz8U6WkeEeK9fNyYXDNHOOYtZrzhS2f+eiIZZRA6PLKHy/VMJQIHXsPhM
4/hZG9H971XfcOjnevUhRAK65gP9ZC1dy0AGX1ep1vjnJtf9oc51KSV1PlyPrFc0
gswhcUdc3ezYhVFYpzs7nQ1rTY0FSR79AwFLpCHz99pK8LKnVMGomTNaOrgpKdqu
SFjJhKV+/5uFeTuu6+QkCRyhAW3lPTkIIj3lrL3lX6bdNGz/N0V1pLYWyIXoOQd5
N4uzpndQc4DCwqf5I1qDHWTWeRCneNTJmp9q96BkPx3s3CkZyx0paNMy/IOyjZRX
34GqBlmxGTpwmzhGCZu+qk4B9Jorytr8Uwc3+ZJtM2AX2V+pblao0loUJlkq8R+V
i/yxn+lvEtV0Os+7hgZN4dUczxEGioVyK59fKamplJXsmSOvwo8xsU1dTQ0Ud1xp
v5NV9LeDaQdcr6WXC2i0jbteeJTfdH51EFQVcsYZCixTI42M3NjgfUGwHP+iikfx
U9UG+NR7fEltP86vee0Er0IuCJe6LXO855syc/RlCt9GDD7+Op+jPcdH2lkINdXj
lP/3ddrXHFmqyI3GKc4WHPNw/gUCtpG0ZnkMrE+tvlYAra2toeXQ/h4rJIWwtWHa
ukW9wzQvrrJvSR1NMAKZZ/YGA251hrB1xfmfMnOO1GNG8/Oc6QSq04ZYp24qPWg/
fDUqj41hZEbdJ48jXoSQAj+MPGxNf0+Ph0gGccdM5JUlwd3aY9I5iwttDe3rhFwb
2xeKKom7Q9XlcJ515yPKdBForj0K7kQLBss5MzLi9cfPFCbCLp6pv6OLrRYel+ew
ZHc3YR562FcjPyBBT3BVdZHnp4elH1WF26ayCmMg3j0q2E2iB8X+DkVn1BCEAxyx
Kv1e3DTa4kvLgtokim0G9BegPESVLl6Itimi9gw7dxh/HZqEWz0HAX/fy/1kkb/j
5XLKVH6F9vxGGE3h03rzZn0F2aJ9RSeEyl1BNJko4d08E2PLQbbddLdxG/NY+OWK
FXxf9N2a2nnZTCXIB//msyMEKpHYBtnALbi8J5na+aMQqi7/QwVQ/qsvzgDFdNJG
uTOfacWhe+Lh+VgJ7qvqyBETqYhIz5OobYiP2+jffq4fDannhTJvq9w9agYS2EDg
vxEU89CJoBU4vf40OJScy+Wh9HiFaHtZfmq4TD9BEYrfLDOcbVD4rcjRtYpxx7hK
IeWjaNtbm+AA9WXHlTWr+FF1wlvHZGW2XsbuL4r5+dRzYguFXiup+oX4dlqBPy+A
YNse8T6nOU/Dk80k/dfnioaXFYlTud9jXSQtpzQG0zcEcwP8bp+A0DynoqnG4Rvo
ypxGhAIkecVa1cNBFNiCdBRssdU98G6ePopF/CBerArG+JEPDsK9ZqFTYAhMbcNE
rPl6I5hrMBcnyhvp3dzXwBb7dKBeNEq7VdsKjm+u9JENnCnmFazzaaaRsUgfy+Gy
0fkgua0qZAm1IA+yRgprXA88qw6iLPPZy9Ga5QMJcBOFRfTibT4lBfHE9RJJCMUr
1L+/qME/SSOxlvOqxn5OdUBVz1dUOs+nrBAX3nv7OSsn8SNIUVCAna+7J2aZfaoP
Aaof2kZYip06lp48O8xNIaoTl/TFq1gHLU2bQzJSaAlgjlQfskfRncy5gwcuIihx
Vl8U2xdXOJ9rfqifp0TkcmPVp2cWajcJJrfzOYVYu+B67OA16HKs5yltfO+OJgVp
fbOz/F9qG39FJbEqMldz8c8QZRKhlZELRtosDyuralaFhLAhoFD9t2Ri2ffxUAID
KofV5MyE9YWcTkKaq1UQaPd7O+xPm8yykrO85oUVa+XyFNZ1IBRXiKer7sMH5Vzq
Txgp8QRnUXMbRjKPIg+wlam432rnqnYO0Xk8JCd5c2iUXCeZDDybph3F4oJitNIs
Sp/vk/ERR16958QsdqyJjtCNqWk3joU3CA3CIGY+BnJR5fCU+b1gF8gr8aiUOtE2
+z9c8YFQJoluZK4NLsgsW5/w/BYdcwu9HPJLjGxdcQR4/pncpBwDM16YMEEoj0Zm
eIZPvn3ir8yY6hPcAYJpq8+SLv73qzfykLPvpcpyqIEsCmfRIJ8M4dnrePKJiywZ
A5z1xvOYcHcotT/SNWQzRysi0vCmtdUiz4db3xR6mh2f9Mw3pdUz/gQd3w/SdwPB
OQp7h+DhWBCvW9Nhg0Jpk0Lcgx18h2HGDLVYi6VTzm/oItcZH9JYu3/84MxphkfS
eR0rbprire7CcbZpZ37d9y6HR8GrBRrn74evMBcY7mx2RCZ9s8OKCdKWZ54EmCMS
jIMpdmDjBBJf0QvRIiNgesYZ7gMF+nf/jlX004b8s8v2QS3X7JOV/TBfyVhOMTgi
3dtLUx5p0VSVpid1K/0D1a+DYZGKYE/CTSMxeQxHYSXPAHCbDLd0mDXJ3uv5sn8K
TXcPUAHOcUD/CRBv+gsH2GRfu1Bu7d6WOyRPiL3OpULnuKoivphUXvilhSRPaXM+
NdbtdWJKeVQq7axQBG1sZXNT4qyZ5+NyQpGN9rkUvaC8z/+/auxYnrhw4T9dkWFL
mUZ8gNcWufiExGKop+ZAWHd9XNqfAYhAhN9g0FX9K0zoVY816nQ3UVYTEEGlIG3N
okFad9Ytf2HGPyPXPM2Cj5JOqRZy3o+U6O1w2hqWWb3If9NALcR+2btMa3ZqIUVS
YAwSgM+eSrDAOG3/B7rnvxvUm9rlfpSNi0dvzEITIyExPlASHdlxBUSfbo+MZfwC
8nSjwwRkglNC9gw6T50WbbTuNWnM0Qw+FCLhe239Nr9OpPmro3stwM2yupJF/f2l
160sUffWGo9ptFegWj9IGlhlwdpQL7URPX/qLctMCRicr45iFAAXafZdBer6G3oT
8W4K0SqWm7cOXDVO0li1vLKpyyN0ZSbXS8pD1Z5Y1G00orNi0yoHPoC31ujczXW0
tMnisnZV7lBBjmvDTZdfiD4Oaj12kCK+zpBBa7b6W3bRxokRdTJco+iNbHXGurnd
GqYMRZ3fWEVyZk4BxGbYCjMUfU64YdsSOeklVpr/OZUFANm3nrz7OfNo0HbPtHrC
ur+sd+5zlnnPoGigpaECAGR6f5y4s7Q87EjuLKsRnNHSWQhy/PXd/XRs800sxBQC
YBJgOArga85V0r95Jdvce3SmLuUXp7LnWoT36Jlmj58hdm90Q1/bBmm9HeSjIywK
mR/Qo+o3QE4ICywrjvINIUlLW2VpVt69PaUO2r8grFto/90JgbIHrEPzw+Uw6k2u
XLROwyIMjJmo2VMKRC68CvMP3ACzKBO4mcbRkjwUSsesTy+HMxY4oKeL568O3Lbv
gP+clCS25ip/uZk6TJxWXo08JOrlLZr74NxbKvVjGd3Yv2CWFImg9/aLLbe5CBWj
2fgt+wxPSwh3k1LZJ6/typA8kGhtUCI6by4xEa1orQVjE1mj2/9Bn9SjVrIhjQfm
g/vmeWMlBekL0x+NVchMFMubcrQoa0XlkL2MsXS421nUklSJucu+Nz+kWP+JkmDG
fNpfumvWMrqMgXSO6ByxgZu6RiJa/oEWF+9975xAlv89b1LCY33XVVA9P9ebLsn+
qFz/c1Mf8/e4qmsxDtbqdsysWPssDueWkDbs2O8eOcmE6p3TNXHyGINWP/w6chVM
vl0EZes8/1eUId7t0S+118IB2URK1vOQYC4aWyE3oHdTBdb9R5rWa7N6aUIrjRB2
vefGLBedDucID2r1dQ9gY5sruQAK7Y84Ta404ZJSbHXZriRPBgfVQjjQMzf2LbV1
JdsLFwK3V76FtW5aQA5on3Q3HB8W7gNL3Uqi9ZdIted676Chsiv26GtZPBk+bH5N
zlegVpQy/Etx5IZEMSjZ9hp2YmvwDHJgMLtCyFkTEvgf5JlvjD701ZKvSRZXJrGA
pZALsGpKUuZGrKAPyLbLyp3Ox+WX4Pz01yvKd4RHia6QIin0TQqUXLBLYVSjToAd
UieHEb0buk3VT8KXfVl6mPfAF7PlO7/aZ7shgDyESjoOXElUOtsS7PwCq0yHhLdv
KNSzXdy9J+oZs/2SES/YYEAFgpFlBZgFjNyZakleMCJHPWn0BCp44rZUm/LeTiRW
Wt4W0DxJKYAHy8PD79oiHbRgQAFEdxfmEjF+5emO98vhLC0w0d/LqvgyQRedCcFC
y15C7fZvDoTJHSUZ9asLbDEQWSUEsCDdK1XYQ/t/uYHqZoJWGCHwSTiTyBzhKWge
MoNR8Z/5G6hZdLo7rE8IwJ/q0E80w7oNXJmqqIare74vsysx8zRoOcJX8PpfS3sI
LinqRbTtTaAOlSbtBhAVZdbdg42dWewUdlB2olR+lci0mFKa7tGHlSjnvPgG7nwm
hv3wr4MyHbt5ND4JgUbj9i32f14WaVflDjqCGNFi8tD2K3KR7A1qxd1qSRkqTlLg
dpnnWWNizosXHgrx5j2HB6D2GRMu4nkXPJjpYxj6zP+FtEMW9Uh831/LoEXH3slM
ueHcCd4CVoRx3regdjLSHQdP7b1yGGEvBg3k6O4/TUn3l9p69xP9ljiPZ+gTzZzt
ko8eKBs2x+lfu6BCTfVhBPCvLiipfFNN8lK+FA7Ixqany6gWFlisvXEHCYp1juCh
G/Eib2nPvBU8cOrEKK6Z0fkPQ5dT4o0WNLxXOH1GgzAYtZ3475e+csy9Mxz9T84E
txpwwNKpQKvpbKMhbjLLopG7j2DIvd0ViRPvX1pBmasGZuvS+A377CaD++tRO35N
x2GOB1TXr1Dk0/9LRRn8og7367gglrECbPMuyj5PZPvmiEqmJD0J9jGjPXs0uyBs
lFO395N1rcD7ax9zxKF1eykIaxHlHkKX0l7xOVvngqV8ygK6JbISS09RTUC++8Zm
616+XcNTMF/iZJJiN5Lvyzn5OpTrRruSvknotkRUil0Yao+vz7sfz4lgQ1zEKAto
WhJBjRWKUPW0s3MTksKQnItJzt3gn2zV8PpXO2tFfd3MqzwgmTDY0iGyla4CSB+d
+Z7TWEc4iUwIuC14r951AfIUj+9hncnLHYJ6Z8Hkbg8YkmKmPvqlU1LVUxWrsM5e
PL4+rn3h59wYcI3rf6sObf7wesYhRjL8MDDugUDZycLMfhWYgPb4OijQRwP7LbsW
Vm0irtseGrNkoFP82T8TqyGhzVbIznTMffAooQBE7zjsbzSb9XoShPTXTUgfThex
NGhKkwtqg1XYv9+TgyAIYimyhpcJvkf39utpJhe22fAu48xS9OcyA2RY0A3aMQeS
P9sMrQBzwMtCIO4NFxDCJzEvfcPnqBBbYZVmjFVYpMt/bc2nTXR/4qwfgLFrDUTQ
q9hnFgP1oLsa8iKjjbyzZ6Jbb2QbFEiRGBtoPfYOPXyk1DGOtVKO7PyhyuWOcFlZ
bPoPgtj+Yr2+v9K8KNpnvfQPGxSUBWTjQZQYPrxu3HNVOnpJPjRyU3AUhRNY5cNQ
YgA+RE1ZHvtFl9x0uDX6TLDSKKpFUKvgxHGXBtR5QgoChsElwqLJsCbuKrtNxnzC
rCbnof1JvDjoXXBSdBcTSU8rUF8SqP6e2fq2prfXv35lyHFJRMHWNJDTe8UCoK+9
+5/AreMv5eAqLtJN+YJ9CqfDzD1h5nRsp5/0FxcdEZn1NSMEF0SbfHonJOdv1kYb
0kKlm3/xibnmw9PoiqjdTT48z5FQ4ntMaqsH+vpF3Lfy8OicudExeYOGi8+vpLiF
JO3VRv6d07PBTYV2zRAwR+BKPfZolL9VkPb/fDham0J9r38W0wPInLIKT0MclRu/
7WWOM4Luz3VpQQBVXwtHOj9jf/lv1fGrWWqfyTbloGnWUQECAQDG6zhaobMbhLOJ
7vjtkrx4AZq3IhggvU4oxF4W+SQoqbw3PlA7QarOHGQ79M/b1HqTDAhenl+6WEp9
eUGYM3Nmx5ewhYRBdayouhQ4GvtUlKaJruZmsFwgfkcbfnC9EZsMUS+FPgd+Wz06
RWTXMh1NK7bAeo/QyH7M4Byi2Emg5KpOrNfRvhqFMI9jG4zU30TKG1r+2eESDMbx
wj0Yh2/ncMLxVurJqYhtYOvk9CvXEtk3uGUOmlslCEA+GDTR7SgVyu482vV83kFU
ImMoLhgpF6JrwXj/ZhH9rxRar2jJXS02ToYlMLdp8kfleVcfg7VX89hAq0BzKYrx
vn/yblJjXV3HBEQ7hY3ndDAA+nZbrN0led2iekprurzPz/WLYANiKHNj1lGdQNhJ
pf0KF7aMTpITcJnBSn9j/XuJe6i04DkACHbemvVC7xoyj+2Omf3D3TVTIDv31xfR
0RZ2lx1OAWsZLl1MZ7Y1+g2ttSGEtvqdDi3Okr0q0+nyKlMCgtO4wSb1Udw+vg8e
dm2eJGsyVX2jelP7Cms7QDAbrEDef5ShPJ9lAj1KoQrsvO5Okeh1QKNVEFS85zG4
fLT9vbQya2j99UcqaRoERaqLJVK5Ap3UtnSp2fDsKdsgjH7NwGR/5Lx5h+USJB9s
VQTfYz0PN23VzCePrDN/fjoPOY4D8HF6/fvuh6RGILYbTgc9cH+Y0WCotTQtxR8W
k7CgMxWEeZKz9xNPDe50ikkRjccjNfOJoq8yYJ4j9UI4u19A0KgfF6ZanQPYsy3D
CqonvOJUv0Jl+wzrX0nbnKE68NV/p1PXptJcw+0lfEvsax8aJ8AP3rLFaP1mHBtY
E7cO06ZmSBdMqs5MM3OLL7Qb2PWD2ktZtRkbgIHMU3w+lvk6bfodcWVNjYR4wq1S
RG5kYTAWz7RIA6Yt4s0729Cz/LNaQtGKhIYck+T33jpBkEUXQjS6gFaHCyrOfKYG
tejvZoPNkwwwPeAeJOxUqrrP9nI0QnHDIVk9IT6nmNNXCnmjlhZrR/ufr8U65FE+
9fHyL/iAHxOM+VRF7+ndKG2u3TENQsi2rtPTcdtpRTFIP3pbiLEc98TScy/cIY9C
JzTrLAdMPsgsOFL/pBoIl7Vt2cU6Hrd0Sc+YGcUM9Fe4JYhI5HqfxKNdMt0gDyHJ
qdsn+RgAryzybErUjIKM8/pAApT4HWbEY0ZuEitMIi95LLV6jlgPyqWoYaQSg8FY
vkS1jri3+3A9Rh4jtt3YwGRLk/Tq9pioa1HpWWj4wnlzNCWyKi798FnbjLvx4NBL
YkskoP1jELyDqm2RD+gbRWRSPM6DWBlNBykuogS6YLJ3t98lReuGyqeHH2O12IYB
cf0+TIO4TjWFKXIvSaSisx5IvZ0FeCf3XsB4tOWSRuxH2Kdu9S/I5wb0zncyv9Jj
S95djdHmdzz1hfDOM6kxR/dm1CtQ9v6rfoBcOcCesrr2j5oblPBFKXcOWjWp4Ead
DKH+lI15Y6ZRh86o85YGQuyk2tpe/74Waj1ct43Sfha4bJ5OpemOZJkUdvb4/rFq
OGpTP1UiKl2He6Tl0bXQyXyPzj/9v/yU5PgJrw+3fmfyVWEq6DAimEXFPDR0Rnha
5ZKlKzIB9HHb97ssaW2cljnLFmtRVI6SW6UgYZYqa0knypBmqNiDTJoFmA8I9WQr
UCu/bcuRDo9As7fzsSqNi1cGC0rYKOVyc3jPJD7tkohEgZQaI2tXLTSxPjYmbVju
4x3Y4eZ5Jx5s2npJIaHMxqeKRr7HPt2AErNwsC1wqOPK5MLshWwPXVcf5oZ3cwMU
iPGHlfI/rbrgeJvot/BQoYA3jiszW3fdkB2/hGjMNLGFBrf3OaV/V/iT1UUMUMMK
M54lo5jsBh73FdW6+95HmO7sdhLowjl+e6qjixA9r1+3jF6k/b1XIYPQzigpiolP
09eWPEH1l7AFnmyjvL+P0nPU7oRyVMxp7b2scbsRNT7gxv5ryOlZI5DfMR3d09KD
PAwDwDnVHwq4krwPwH8Nm5TZOIcmlVEUhpncYHGEV2qEzgF+P14czJnyYAulzpml
BxE6fjbHkpiZnkeqOJUwRfCpGRNZMfnC2bbV3xF0++lA9Wm3G8HsqhKWr8Z35euF
5JSAdk87LrY79kFhU0UUFXZv21ekJaRNxAkL068UcB4mjnnDD7G17BTtjRB4i794
7BplIuRS+3BCvFSSilcJuMBVajIJ1+2TC5UErY8N0d5jYFy8QKU52hUtEyHOLDn9
PhITkaqOxuwu0CRWy4twHZpeknl1xfotkpxE0F6Dhg8+syXIq3id5s1GyHph+jln
D/09kdfbzpouxuIySSG3g1rVL47GG88mMYi31d8dxdT5dQ0NXTj7+U52aJzzsDM7
jql0bbqxXqkkkBlz7s3JINZrsVY3L1x6pikIHb51mB9bGmIRfdf2rhuZVHEzV6hk
u/sxxGlQx8DkLX0ppo3L9ExtLTUh3e2ZuC95oFQn+CNa91jBFA+Gj3JgKNzJ3MGh
BsajUzklKaDKKNLbQr4eumR4XtKXcIP4uo0DHSeTUrtLVV5WBTZFmMEFZp1eR8Wu
8e5dfLoAL/0EzFHjBc+PTytxGrGjE6KIs/U2dFWw+Q3z24fS2e561l3nEAypaScb
IrTaF2QbeKmc0LV6YF9aOqVL1Sfa751zos/T1l4KlwB+JAD46sdQvmkcyifio1nk
sqt/m8KNP8FR5CgR8zVq2sUK1ckWxWJMVFKV/Zocz32olHy7YzHSfPZ8ON7pAPZx
axhVIhQ8xMg5dp3XFnU2EXrpJI0pTnO1t1uG6p7eHxKaxmDcySFOo7zsyjbduI9Q
2Kpp0JVseR7a1Yi7tQprZZWD5MNU8uAOXU91QddqhsgNqw/cKI5ru9DiXG9JkYvb
fgR0CLdaigzQO71QnzkrINrK4Ir5Dljy9dpYJZvhTrwIT6XhqnFsRgJ+1GXMJYrz
/MqnyKwH5m42lNBNJpEG+AmSJ8WIxJrhN1EuqJjDn9mW2GMZpaRaYPUrA63htmjJ
9WGcB/XUJRWAzL2yrZd3MCNRzpzVW5pguI4LYV/3Tzlq5/ZFlBPkMvFV0sbeCQFk
r2efrKH4EqK6db/q7vqZWUUbcoJlcbcNwr5F7k8JXdZM2n8hbKxPb/f9M1jAfnxR
SmDvz7Q5ff5J+s5ei2PsWO1A71s5/LECUy5ZFHdnR4dClHaeX0cKfiJsjCNYS1ME
XisJQcyd6FAXTBZgzOv19OuIc3Cewhxa0a2MfGy78abr95IPLRV8YWF7mFPHSm5+
lXte1Hf2sXcA9XtUiEewrY5romOfSapQmAkrhgzvyvyPMX28GfkzcvCvW/T5TOL0
nOx32j9zlqcZPA7JmoDZqgoi1vNrVMZGNtXlombJAZzYeN5/g0uI7JxIqDi3FlYu
LX3LrCzfBJ0A6BpzAlFuqAfd+a1yV63gf5mOju65omg/nKarTjJYlu2pnO305CTG
nfJscnkIhmQeJUk3KH7OF8PvTZkj08+AYXifDxWB4Akn0B4iPrw/gCVw57rdOp2I
955sm4vK8oX6M0+hJncDcuS3rsJb23wfjxSc44ZGKGSe67PyaakuFHBjlTmOLaov
0+rT41I9Lz85UOQUuAK53qjtFD9Z3fmEbCFgBGD3MCY5g2xZBPDRP1N+VIrqavlw
ITcS7m+DL6eVjsNK8MZfzDQUO36CruJYTJnYrnL5VbcInxOIdOZhhvrhAiZGm/Jk
eq5SgNu1UGMTOecCYGeECR5hDgSuT2N1SdaZl1wtIvttKM3MFYTjEC/1pzmRqMFx
L5T32FaIxg1t/8mfzYUDmgnR7ZL+LYWvn/5cRYZm2wbwEYG0WkSsVzr4ca27qD9R
jPyo4v+hxWLP0tsfdjIk+c//if2gfCiDLLoZjpzMmIcFBxO0vXESOYhUq5V01m1z
lgTmC7GVE86HzZat+gIzIcZE5yobKd5xSV0xyB52YDHuOT60mbq/gqJIdl2OZJMc
YpumJPIpwIXhULRXvApzU6OTRKzt/exCTtHYDT/C7rl2XosDnjX5B938OgtaQ9kq
a1RjmLT6LTFjksGN2wvReBi55giahaRMGvq7fSOw7rRwaS3Vrt6nCCfciGTLqD5m
vOflWJrEoytSWxvwjv9mHB4OCok7D119KR4wlT/siDD/ewhVcSm5CYtNAD9l4xhX
u59mEH5N0kw8RMraRf0pGR/wuWNM5IQBJubjE2xwBmG9Eufn9aWZ2rvpF0NFx1sj
1kRiZjYkpYieITYxmaiaULiCx5ieug2BALjx7W6tPP0VBb23VgA/nW/cFvkdJoSa
Uvsrxpup8rdvYtKpQkB1lW0lkcMTVCUAczT6cgnwwCqPRl1LqhNyq59R01dmNgBa
Q1/la8ojFQ0YINWy8wxcRjBmhZuRA8lFfx6g5nT/xT3yMzliVnkFpOTnjPREvuDB
yEb4xrtSvB/7kksFIE3Z6AeiM4LBpUR6mvt5N2w4fqk8BVJfqkRjfdQ79fjuZ023
xfVckh+siw7XwgnW3dTKs9kdSAn0k8FcWWUw5l5yrCKx5winVuDVvtlviY5dnDRL
Cw/xlSl291k56mnUQpFHu6LGiLdsZ7EAm35I1XSc++dA0uuihCu9p4Cq+OssCWMp
K9b6OgupBT1puGZhPyhqRGcoRcGF/QhgsS+/Tol9YyyYaIJjUt0uVkkKmo4Eay/d
Bsaq2elTxjQ6BOxdJsBrtQWoenDDD8u1N0grnd7asHbgPgWQFBH0H7kjPLO3Cme1
8oQLlwfpbXNSfDMDAdyV5EtS7szvpjtzKkgKyPHHSIzr/U2gFs62TbaaiYjx58bG
SG9C2rgjkbFT9JqI+Qbpoub/AdX3/tuaB1VUERZgnmJlOdNfAvQw9YN8uP5HtAFJ
4TGpEbpkHqgmbZ/RnPMIPKEFBLJkxzFCFAVIgeSlKcE7iF98c2PrkNlTeaxwp/S4
tS/ulOmDF/1SHO7Ai3UZPEGh8OMYkNg2P1WwFX6rHJiK29Jad9KIrItesQF5nXna
3Np9PVqCuMR76E4rREAuOe/IpFj0fetGUOf4UvrF7u0TF8zMoLA8xVdKocM5P+hM
8OLtGku7QRM8zzhHFyaNHI9os7Y25bt93wxaJjlkqC1OQpi+fNFNjob0dj467mnF
sAQJKF0h7hpsiEHqo5M2E3e3DTsszx5jHS4Sj+uAkCc2XJZlKO/HpojoLi8iGmlS
MikDBlPu0PfFQp87UqnXswbgAGJSATIrT2wFqL4aqPpUKEwDEN5g6ttWg58jOyBn
71LCQb0vzYBzHXIMI+/onqgJ2YN980dcLnxOc97V060vJsoNQGnm0Yzx/+L9J322
8/0itHkkv5fLWmOFD1gXPm5QT7xrgc9JcULIfPjWrxHqNr4AOsFBbCsg4llpWGke
CjvhDNyGCHvUThNHn/5FYXuFmbR4eNUYHlOaGOyx7+MEfhu8kuUeMHuvHP+DRtO5
UFYFwMXaMOoUL5+ofxfYf1y9o95v4eQoHsDAx5Dgf+Qj6L7qgQvK4bTwrcSbGJ8M
8ME3Gw0eT/PfWmaEVS/lAtnde4ZZasbhSqEarNmUNcpya5WiqlD09xovsfSVKJjM
Jbb+gATacLTj1QCIxerYbLBgAvVfxrx1BCJfxTnwpJlLDVC/Pnn/iaZx9dn36UX2
+tMJ9xBDkkZzaCg5GhR/NhJffFMY6riuvarRqu3XLr82tmoklXK1SvRzjYbxuyQJ
8wrnzUo8JP6safhV1086t9xw2/iybLXXMpZ0uW5emZoqPqxnddpHLhrPU9PNxNBw
ebGGjPn3xmipM/+MmALFrq78QtR3fneYw2MmNAKJixPcVEVcI3fjsaNblMT+4p9H
WJvTJdsBdnK4+QwjJ9ZA/so73TDU6XT57fAJvlltgjM4bNZzPhhnTFX9V1bu3nGS
zlxnMc6ymaw+nMwvW7kXdBAJdAtWKfejvp3fd82F72f+JHQ7uQZdZHzTu9cTGhOW
OMTWMON9z1oW7s1DLGjUC2l6awYFdPz6ZrT8d+b6THZObNkA+cyLcUB0+Wskg+xX
tSq5zTF3zMDWkgryzzVZG3ervu77X6mPLjcbeA/Ywpuit/eQkNh5+zdD9P6jmWUo
+TYruiarVw5PkDY0eJYAH+Sv1ti1Sq48R9CwYIvhOeELy8zNStsa0d4+v6dKN36P
9erXzX7/m1eUQZdi+M869hSe0Kt6r4cp3Rt2pDEimiSDZEootVwX34CzKclQASDZ
elXpw2Xw/EZJ0hiEmLBkDGSt57os07SYHtYiqLZ2MuEWxFgQN+9bNpjNNKqu6Im6
BW+71LxZvUwIALmkgXuDzE7IaeAJMRP1h8Z9k7bmr76xMXCxK1zBf3T+yy4AkCnd
uK98Pis4sTddgyBfSEvO0zGuLPOBd5hSIaEBVhYfHhfuxAqLKhCZmLlclsVR78Ok
JijhlNRCvVxCyaS6DH6Olb9qFxOLYzfPfVksRJ9jiMQqcRKfmz721NLCnA4194WF
qWAaAja1rOuwlWVZRxJkqFV4AdjjKI3ug99c3Uxp9587SAJcYuaU8MXNaJGnFXpE
QUO8hh1fHjskFkyIw81QewhIeatsLhEsQhtxD5sLf3V/x7CNRgA+y7cvr5OlhJOa
Unjf4VBc7Zuo0249t0fHaJdVg0UrZ0kVrhXRmD7eJd2pKLmIdlNMKllFUTRc6CJo
gh2jjnCZJg9cgi2EHb+ycpzRz6khHjyEeLyeHrttM1GaG7YiWdRy8G03Kxq8OpJX
rkM2ljujmwiuSxWb2GuzhhsxX8ZFUbJ9IawmfYK7SHMbODnwLBOCDaedmQNyGkWR
eMNCFGE+ONMbi79GMv9m3ukiej/6Q9huM86C/AXl5IDQ7QPtbG9u6pn5i7pYQk5M
qR2vFVKkI+17dos4q3Ji+xU/Ru7p0tetzu2kkQ3EMcJGc3u3ORkjrZhRlmdwA+aT
li3rPdCEJIMGTB3IQQFkEtZXCou/POf/kbsi4cldvgIOSgbnfJwiooIvAJhH+9JS
MBNHt7CO4CYs1dTISSrlP1zroh5vUf0wd3+9F8UBTaXbagcsRKPgYxHKnv0xkaMF
iwjo5FPK/hLg59gr0uVUmYRQeKmjCNrsGIGqIxJmtPESgQgyUBYCvB+FWzjc33GT
GoxYx7JfPjuNMQ83O8sH15+Mqb7RDRGGd5hzUHTv268CgvrskUfp1oemZX0F7ax5
4zTnblquOAEXVOkPVdKOlqSuyWtnXff9E26RJfHbx6SqwwSJ6f2VFNAikGUOaoFN
lSnEXwaKBJCBR3Us+i6f7eNQJBeR8/cN/FHVv5lIqpxNXf9scu1pjNp6eSqspG7/
fyB/73W9zm995MZqehApUH6HZEK/cZatmwj739ZCIFb9s+sTmjjgMKnwafrODsRX
wORsi+ULvpyybgBl/YbJ82KKb7EKYX0P8wKr8/Crznbut+8Yvl1vM95LMdztIW+U
2QOMwT4nhWwAMe1WBUMPYvRBzLWsxYjd8TvXACX3mJIK7e5gRX1Zx9ogjv4kNlJy
ff9b6droDviirmftTDMNl8Fyh18U8pVdIpXdpHDRJz7y7Jn1lW7xA8+4BHcdsMm/
wVGqxxc3FzpojTKTYJFAEJ0rbF+t76H8Xyco8aoWVC0cQOu1R/ueRvb4umf0X5zD
fgRGMXRaHbHMelQtRzNu+uCRg8iPHH+FTllriTd6qrZY/ibLUe4WQ9kCkUWb+5kn
5ntZMMNxpk1z5WWpyRtZnl1Rdr4+euN1hdelBWtUn62yAgOO7aywORL2ysND55Cw
R4U//E48SByysy6RpYSzlcVRfK2bQJW2/9CdQJBTZQPp52VvSeR1zIMvSUz6gkWo
ILykNyt3Ptdc+Dm6TpUDxciQ1psmUTCKzqS4AdIIJ07ujEiO78uNMqcHDqKm+xyq
VHXQtrR4MMivj8ATL288ZMQ1cjX6h+6+pG7uHgQ3LaTnOL4eRKmkSQybph1yKlST
3bnnc7cb2HvxnjQGoVV35Vc6tAgS8TSsZknVsctEoQDUMX/ESH1U4YuhaFJxg5wr
UHXkmhISS8uNU5w8+UWj2Yttk+qTgg6k4EDfASd64S6mp+Yn/PrLwCFU8MOtLtXt
3hAYIKoCoz4BSj6dtGz3FmAp200kOiDfq6wxIOH1Pz9B5I+c6grpKF3g0wcDYRCB
WW1CIJVRo2RhmhT0swRiY5DsKVctpuVxaA6GUSVf4bDHXk7GE7+urVdXleTd5ASr
rTU6ElVkrQbVx/FRfh01e6m7Am6TAL3i1hBR1aY3xEmw20u6T7y154SM1kCm/BuA
cVzG0uKWtxsVBZL8aF0v5Yr9ldcc1pk/KrLISPHPYJKq5SzSJL28kHqOF/eiq0Bv
LOpG6crOnwvOFYy+XVKJkkbmmJ4h+CP93anUGObDW/OPqxp/MZ/5JCN5/HcTdEa/
nzNVSkSeEhmKD+f2eFOg1Mw9UUOwhdW0/qIvpm56kyvYRdCs/ZU3Wlyu3m6esGe+
Ege6Fax32XzloR3YEDWC11Xb1qQjTPOZ247qApwGdYGU+bnUgeftiKQZ1cuxh+3J
eEn91AIE8bByjPS1iYsHhjTpl355cERKe/rc2jUhqyCk0uxpE3XLUF07UwBzQr36
x8CaRxmzeC08+hBNhod+2X2d6wuQQxsvPl3TgHs5Z4fKqmcjeswXZG9LIv/D7h3a
gaSCrFM/MpGq3MZ5nTkbAVCczUjpwG2lyvaKR+NknrQWx9TtBDVN/kNj8L0Q1X+J
6J5Gx/1nywY0D25XV6nGEtIHuxVEdWVZFQyJtq4HEJxpEfNC4RbCTu3B1+KkCT+Z
t8txxJ/k6blmGG3UVn2pDlabvFtMXKqQB4PY08JdGRX8n3Lm8Xn+ki68MnRf+t4k
eODyy+HU1+GyFdGjX554tluyn2pm3ZfmkhE+69qJp4lw1VHbKN2DWurPBSZhWb9u
wF7twn2N5kNxJZHkpZnJROFUpDHZlJ2Dnsx5BTQjFsIN1vUpGgOm3mzGZ3EUModS
3drMSEpSoKDPcCLSonOHpj37iE9BnHrCsNi1pYVmgXwOqpRospFSXq/PeGyPxsEM
iq6wwL4EdCNf3tZw7hNZfOgJS4D5ulIn2HnPnRYzVHOnZSmRRyqtlu3mwt+HbjJ2
uiVhR81pviwXt4J4SHp7g78MChwlZsJgkWqO3JOsrCb9HTZbrjJcro0dcIcIhV0m
eN/fIWxVvbg/LZaGz6WfiyFGtCG4FoMiawgXOV1nSw+oWwk1uZudOuHZDR86PYPS
+/4Sxt4zT7O149U//Eo1515grEmT562bpJwq65x1TyHdF5mT77mNmfoDe5TiZubg
2Qw14nX1Q+HH5Hi5hTt9oLUq1SjoWCz/k2wk7OCVMW9Ch3AS5LNlpt88QJnGIwV6
hnh+ZroD2uzcHIaCnJMuvGXHF4ERWqozQygFpeae9B2nbq4w7UXK3Hds7pNkn7Np
UQ4pu21Sxs9s0sIuOrE+qUhIzSMJYSJ9iQtmMe8CoZMdNCHDoRTZbBmyiKRtoKO3
u08T1W0hJ784BybkWEFZbxqUiyIHZV/hSt2iPmatZfXW9TUpuObJa8CvfV7omM6w
944HpZfJrioRGSU/duduM5ugkTySU56rbL0hLb4hpJnYfhzJTxt1FK5aTC5HcKC8
KPSvWjbMamvZpBAdJ3KAD9JpqJFV+T2cOsEEJEbsxp62HWR563+8gpjeJVmbodbQ
LYAvzxagw9vIp6LIz94i8g+yNUrkeXEwklHu7GPYSFN2Gzlz2fdEDCInLHx+fagO
f5yCU0gwn8l0RwXhnxnLqf3ndWWAkraRDe4GQA4/x+tSml/fKGw2D0XqfkJm//VM
ZD+CIby3athmkLO6lB/bu15NsPCxHy9MuWAK6urvr5jFGofPPdywBC5ijXcvb6S2
a6zyu9BZrzS8sjqpIlgiYV9wGaY59TZHXZejKeIoj97Z/WOtAPsEkjRv8B2rOKiv
jIqpocdH+rqbszqN1cslGqzQk2r+pL5Ldsdf6BtPepAs9BxetoR1b56TN01wcaHM
Us+19mkF8xxvCjgSnHbLI2SOCFQ+VW32KWCZZxKrUKSguOYFhTI4OiWVXuqIpVzg
jrHukZQirzocefsbfNUdXFgrxVl/fuHzRo8SdlZbrbOvAoFMSXvC5hQR756d6dqG
uZaB7YiagZkooZ32YZI+/WIwYjTyccp/jryUz0ZjUU96I1zu4HXks/hFWlUyrnTl
BsmdxjvikilUTB1XHnSJD5yXYQtd08zH3McQvhN7MFpBb+T26bfs80gFr98vfPWw
+9Om5Nx9/9iZytxLgu2F6w8Fd4W/6utWhiupU2e0ozV6NZc3EZAuRUdH7nDGtR0g
vS7qVp9ll4S+67/oHYik1OSTDrfCACUOBe/kpVA4YqzKvWkTv6q2R7cjih8nmiT+
c7DWX94F/Z7RfzV4Jtm0oeDZ2t746q02K+mcDPR/Gox6SqWupBFNv1q9GNA5ewlY
ymMaQHuld16vz2yCx/83x+LP6ouLKd+oPJvOGLbU8ZB6BYI48bInW/CjsVCtg2MS
YrDk7/CjyPlZ4rHRBZgnTvfONjtC4wu6pBjSOrcPjPYNjaPzJ9nc+F8t0Khle5Xe
F6EQxiEsNgHeSETI1aclbGo0i5yUd83MKjHyFofTLuswxb0fP2HObnPuBdm+Gb+h
qwiAvyP95QFzACV5U5XtwvB08q1GcQvaCTNxURj8vdR44oWyI4fL9SPD1CzBUI+M
y5VYuYfXOUrIrOTqRtAMZL9P1oZ4isbHjPO/fpUZcn975pAT7oub/pLUk1cQXbSR
pABL20G+mzvoGet5iLvicxEKRAsPymbEo517ztvbkF75i2TqDjHbpmC7cjVDh/YG
j4baYKHkM097lArH3uQrXnvIAeH85pLxKFSjMhc4dTCRr9scuA4CypH/Ga6z8g73
alA3x+wq9JclHiWnk4dFC0rP7gENFlSulEAE3xhFTOSEwSBjH4nqGaeibzmpybEE
zL2vbs+puN/tTRCpeMo5gvY5DlagEp2RRRExoFz6VzwpJBcKdV3fLE3KgieJqiCB
0AJjtaKPBVxizMxkIO48MG9NfIqRZt8c6XNbuWevmbrihbnHrY6cu7RfptAq0DjB
1NVeIjtsTi4BeXyRdUMYvzMom5EaHMEuNcAyPdATkx7JJcd1fgOnXPeo7DcUqZtN
j9qIHbNLXwHuO3hEbUDIkr3mOX9iWSFA/5ZDFT/vHf5tXRp+MLD8Sx+jO+X95uXZ
I02IEexqXWgMZj+z/m/mEla0kUgcPWvoTiijBRfSXFzjWWQPOWSO3p0GxOXGfRUx
CCbxykKihoIEAVbG4dRnPbTs/cg63gKGb5hnHNh9MODoovDIWb6VEgmrcditu/26
XnzX1NjJaF15lGgK7RqttIpza3ehIGMgjPKDMj7iI08Pa34lPnAk/2t3iw2dovKM
lk6OuA+EL8Iie2fT3Q4+CrHT42q/5xMhVZPkF3kgflO9NFkEtS07qqATZUNuW/u1
3Tme2erGqLDtAS4/EbzzXMKQXTIzFxCz2zTT9KbJdsnMR6EVlakQ01XEWvTKMk0t
0G9AlHS1ovjUt7d/tu2PakKqbv1sBQQawYqBVnBCCW4Ro7iRXQpqCchnujq7cUED
vK3bX1yy/TkjnSQOtaCfiHT7fgXxIItF/ymkZ6W121ieMmrp+UvEtRQ9x68yRWr1
8G5Mk9lZSYfdgaw6/5puO7FHrnxyKa/2o+X+OrDLKl6DlSu50pxFhe9kp0b0WHlS
h3/M58buDh783qDwVsUqkyy0C8WlRgDfR65eGUO0ryeYY+94cRl2JlvHCETtvatL
x5au01UYCoDY/chdPK9mipE5B2Mj8lXdZUXJ+vFHFbmTts5uJ32Y44zk/XvDkJix
LG5s4dPfRq5zY/+V1RQkTibmofTv6ZTZFI/mL4Pi9O39SFAkI40EgtUIQvi8YhaS
+t6EsYX1BnU1mUcwmo9zinhyLFH6XMOu4mB9/ichZKYbwbh9TiuZ65Bvardj33N9
N9i4LhgrHWpxaLgfSxzsa2tybEErQLJ+qgGzPsZghUfDOUZccoqRPR9EmuyOfPRK
3oMNCIMATJ3Fsz9Yp0XNaAO36x7Ycmk3/px2c+ob6CF6Jcct2LRNb5csAnu/IJes
nPYF/wPnwETdo75CaXFegi4GJT5qRORTxKSJxrYAWGXo6h4WVCPkLCWt9dg+KKCx
T+ZDleeXtvbXjsFLPJH3LnInVN29rhrMVc9WR4TCqbsRJDYqfWLeahn+wKWPGhpc
wg6PbsKqtPfWSoLZIc9JRcOpWxfG5SrcV3Q20O+V1/nLzhznIhUwLtkKB+/TDzA/
cExRxLpQlPWq7fVjBv7b5gkZ37qehpzvSZQZky63aQxybIMBApqcs2KX69ezWySK
IT6Hcl/Ckrsotey/uAmaPkn5XTVfloqwAAhZbMBZShlcI8oTtKwpMgW6etoC+b8p
3zCfmAvg28uTUvxSvZoHGTJLh3TVFSNpzaIV99Z6XzXWdl2qN4axzyLQuwuY6tVx
kGsCLo2pTgJwKeejwzBEoMJkeJn6F57PJlUbRDEh4+wLp46G54RZuzEjr9mLBqlX
u1dcq9WOvAd8xEIJCtxC7+8g8JhH8Yd2VxuvhfJbk6mdG1rCm0eSES1pfHtUkm/f
aKrk+9ihLMZkgNaAav1vhRUnXkMKuyiYL8UREbDbexFOZ3fUVUpqR2S5FjraUmn7
HSYMc9XtHibNUUVjV2CCY47C9vSpc90etJ1Nz+OR/a6lvZ57e+eW5jgSe4Dem0bj
+AOkXYuBnr1fin4XhGyv25kBY0nvRvGj+J982eSRJbcpLYQ6E7WalEZ2RONs0r/Y
DmXVPO5aXohn0oSRjyY1RnPizL2K3SXbmUS0IGMUIDgKaf+SHqbaBVDzHYeSqqf5
ODZ0MoP1bIfgQEezmfzjLLvjfCv5nyQdwUY84oIZ1zZeoVdcfdf9Cvkqfc19+Mkd
EFZyreQQ0CB/3TW+Pwx1qoGKEOHNKwPAOwrg2aPhHk92rRTYnGn3LZb69gQ1C5NC
JLK+fKUB2hDT7x5eiRT8PkLoNDqUq0wZvktdX+MHArv8qLC8+b40UIihPePX7OCp
Dw+SBxh/+/NgRo6TDHIoLsWr6/y93GuLQPQ4UjSaAH6UB2yuCZIih28KhvrbduPn
h6iyp4GcCZQhHKxsLqTr0tax330yyBHZJXTIEjRIMVCsUIHaAqSCwv1CbISUTE+P
7oASIH/Ahr1i5uknDkb0hxbAOoSm6oVCvHYW0vKQQrHSOv4faJi7DkZdtuLyXJ1W
B3e4xUA2DU3gYc6pbB55B8Bld++IfSi4Z9j+5/1zinqCniSV6WwMga5bT0Jt0daw
cf28dGGY45oIN+wRFgfdBirtgrmHXqiw8JeD96LPQ/9ML3cAA9l6SCuaFA//0Cv0
1XWzt3zki3LQzQEpIECaacFqvbzEhzoXG8KC5dsWV2Z1n2kwI+CMN3Hl0dIlfquh
tjNy7PMi3uSN3AF/J0TSrugGYFSK8CoDV7V5Yv9SbVjqiSUZBXp6AHaGH2X2f+or
hjB0s50e0H4xdThcr3SvEZL7+G41PUvzcAfsq1Twiu1k3H3F4C42irsPSkdDSFYX
xDv4l3xi0wjTW9wvwB4tU4UpITrMKUBTk+0z6tdcYIul7+MWbNw9QgqSeQROI4Dz
Wmh+AS5ztHBdxRZfkUyralJsylWrOs3ohkraApb1vdanjEoBLZm9ATFjj/YQ6NJM
EF2FEm4To+0Ipe2CBf1TtrlEC5nus6KtyfUNXi0s4327ev7RR7JrJO+AtqlNbDs9
4BiM+a+LLAHhADnDRZy88m0MHcIZFscYx1549aE9Mi0IQWb0Yqd1ytzYJpV+rZI1
u/gKhaRlUbcswzK5qWtX72sL+U9D1d4MO11XcJo3sgpNwZOYFZyYyjn+NWmLVFZR
/GKaNLTFlGn7Pr2wy6lF0JRlDgyzaiJ9Ogo4gwEFewS0n0pM6V3lbFnlwnKaVfI/
dFHmh+8jPPloEsTYNDgrQw1fHLPLbMrLXBUfGYycTIKnwKL96kmMywydHFF/+uM9
JR0u/ImKrzeRqjDai5XR3zPn+9mWvMwNSsSxLmnf6i+mnjkHydhxRltpo3o6WsgU
5UsNrwD7wamNbevfTHs0ewf9fSLvf9QnPlxjdg1XzLvcgNrp2ANqciTkKfpquI+l
aI2oRDBYZYirc8rL5XF1oSI7sN/Gmb+ZtclNKoWo6pvImEBqKYWwtJSbZBkZM20W
5zRBnq14Aqx8v+hvJxFeHbVkUX2vwpZeKBnfN2Y2+RJ8+6oi0cqqQYe+XeFRiAN/
w43ovHnT3AB0nfEo6kWlzMMPKUEqvnqTyPmapY5WfZTtkqHWYaLeItOk1aUeiPMk
BhH3UQ/03hWAfCiYwzOxU/fDJAchTPZqdUShjrN14zG35xNWzp97BC3iEdC/Spdb
e605ETqDm75szO7GopMlfij9/D8bxttA5B0nJ4solVc1iSQYR1FAC9pJzdid728e
6vyM9zTj6W7/b18dN4O6og81F706LwadWbXR1Kfu0hnoTDxOjOMBx//E9ZtA1Rkj
o2EOWsadZMutnKg7rvxDTKOSavEgg9x4l2H0LjVny+KabIXh1BxulSsQmZppEN28
EaK520Ar2HzumP4QTrr9T7rRQD3ri8/yNseRh7O8Kn4eNTDuTZCwfz0C989YkLwU
KL5V2w/WMuYPMFwEskJaGtLpE8PFVk/4HGVnXelqmnMQA85uxjahsQU/n1DTtBcc
yZmNUwfVOP2RRtmg4llLTrBNl8l4qRU/BD5WKFXlGkmpiXmm58WjH1KFtVSu0PFq
DDZfI0nrI5nBpXvRz6byxemgC8oBkEnhqDf4zHkyHi1cBCoZS2GTvHSSJRL8Otek
5P2kmpGCQA1CguDXt1LpIR0RebyWjETcw+4YzGIGVYKbwYjIm2NIAeszWK1yPBZ8
VyMr1B93yGfx+XzD0DkhkKjLoDjxJtHdB4vf4KqvhE/PAyj64ObegmG/UZDBkR1W
OxdBEhnQel6tI0rjjwFIjZ0heUCXSIQeIxmUmpG3ABrh9OHcc5KQxizVOrC8B1s6
djJ2aMeDeJ1XaWKe+aIYbxylkYp1tGE/PBT9agP42t0bOulO2PwL4WJOyyDoKiYp
N9quei8miCQiGeO+KYH/IwqlILkvF4F4roTMd4nmdtbadXiQCQjMnXnkAJWXlK2h
OLJVkr1vNhk0uBJU/kU9fTXuyQf+gs4TVb+EQpOxmdx8RPvlI70vnbfSRPPosgtM
2pHPWrY2i7TyYnSr8tQdq7g6PIwJ4UmvZcrRpW1iSSVwLt7HGAoJU34F+m1gdkXz
UjhcS93n12uTAmrvCgDqcVYj8nI1TXP0PfPzuKczxURJ2lkviRe97/004B6fXZVq
Ru/k0YWclJ+6Q+5ewuZJ33ayeE1ZfwSFbOr2+XR7Cgb/myXR4qjnZ2hen2irAqY2
IGs57XXb4r4m65bJqblMniwqmZZL3iZGyYsXGDBi4gjXKkBI6RMjEDvlLxE+cHoY
jKHZi6qUStoeoZcnE6ntBeRR3b1MV+tTnIUWvbBbO/UJa7pLMUx0UwOHA607KCC9
pbmlB67Ob1MVGQn7ghNthyVgF+9Fj6rr4quP8vOCnxTv5U/zhlT7RDT+ufQkGT6K
pOcTLeTLtEy55+s1gBqLSy3GxNmskAK9KNYMahUnqkMjvl6K+pXlYLS4836wr1xM
uePEBMiU4DAp00+ncsxWHX3Mm8r3kfJkEr9EvWgzRXnJ8fAlqwUdknxIPq1+zlJZ
vFk9FXiXoV5SuDSOdJYcy3tsFXekFz1cn9BhGt2SuCNesQ2bIm13AU1yWl7BJgN1
fLuqfTP0ZLkMZv1vA2HbP9WNjkLC23nSIr1tykL//zlc4edOHMWqQQNdJCrG3VcF
bIafROH0vnk+w4fwOuCspRBvoP/FWXMcD2wr9mv+hofY6xVfksO1pYPxVVV79Xv2
Sc+6GSi/9p+l0eAkmbf4BR/0o4qhURxB+PcbIoKjZGXGysBV5Eft5lFD/idg6sDG
vM2NStPu87Ee0UbciTBfopgxD0UzuEHboA+YOlkNEcWEwBGVrMPJGVEdwBB1OOMm
X5jtSrVovkeKJe7yzByktpKaq+Npcm/hFwuXLI01dJ2781uIZSjtIcJcEyyzEzeR
d2QqluHb41BiQA8106Oz99e+yqMqENvnb5/Jm9EfCLZueoYd1R5RA0mIo90VR73l
f8jW84a3yCti+1W/MSoQr6jX0laFUc+ODac7vn/wNm0F2C0Eeyi0rTQZVUEz7haX
rEqv65BLZQNX4r3XyCS8xeNfuybjs/MMkG472OxkML2+4YcgLDrQDi25fUp8R8K9
hCboXc37BdZ+CPWaPT72jWKTCWSdOxpZSofBedLPezBPXswSrr3cVeu3mwhovdIy
Xx4Sj374/PgqMQ+M1wK5G+XW4MLNdPDMiJb+x8Pji0TvlkUthOEcawacBDfILNW9
ws80eJCdNs3P+N/uvl3IuryaoNQKSmtIbYZ8gPQRcQvlBq63OtM0hQTwwAt2Mu6l
IReFBSWwx3f2QXtJBTO4pwdjusHDNARgbzTyO7ImjZWDRfOjTv4jw2LydfTYTUJt
fxCbXS1ET2rnw32lP4TgP72SqzM7kckGB8XOCmHv8gE1D4iD11WV5TtzKL67Uld2
U4WqpfefRXx+eF21yeGJbUrrtPan247M+n5AEJIa4T/r2DL7QUkhQZGqVMt3qBO6
JqPvpiU7PkU0Qp0Mk/CsMvDjbOqsi41XZsZFDvSrMgheefj+hXN7Y8XC4xKhCyIr
2Y1P5Cc4yToeCicOxsrqP8rdfa9tvtFeksaHCVbtsU9ZT2qwaIEDPcQ+qgpDbAF7
37Vm7AybAISqn32jdsvGZw2dC9S+fv5QCJgNRjZHx6qYicucbFIVh3mf/m25v4pJ
LSXsfN/nho4cgPbNE+LHkrjtL/AFj3+2uDy0H8ZbKK00fA2R3upIQEhR2Z0t5E2s
TrPfzLyxkA2gWVrTQDhEiSlqTQErvNGLA/Lrw/hAchBawo70YquogdRg8ya9954f
r9UGbdMfUbP/1+iDJ4y2aSFHaZNiRsB1IAQHugf21f7hTQPb/e6eZFFvDOzYoaN8
qBdb/FhM4eBBPXIlMpUhTDbXU7U3KAsxRe/j/noGE1AaFi8S4S9crjV3rjwCMHdt
5oGGy1XrpVGN4ptOIPXIAP2/9c5BnhuPIif286Kj8vXDhD+28omMEcK02KxENCfN
oiY5QkIZZBix8GEIogwZcMyJNfFe9WtTZgSfT+mfuz6qJV8ikS30yuCsaykFPnxH
cGZaN12d8E2AhN0c0nJqG2GIw0kziqE1RBNpsk4Ns/dx8kxIbtzs6EFABjbmkCj2
9EtOVqX9rfthgshGnn0AYL0w+1X/x0O/PIQRpBgiCFcVAPHQDJpV2iO1EU7GNEWW
ZkpagsVhLzJ2rO/ZjqnQ3eGvX1QfltmPxYZgcAQjiSRS0l+hpqE/pOmr3GFgquAK
MXSpyrbpt1PvCtDhAkkrvDM///FnoJyBRnNU6lzdOSOIaiRTAilN6Yy4OpHRm4w3
iYP4ne2+1vlRKuzjRe5sRolEvSjZD2hLMx/DyQTNQ8lNEXMpJ+ZMa9y2RpbpxWMz
J/s4cu/r/DUhZXaAV6+rphY/CVj4EIx+yOlVdOojlWiCaZhMX6zwN95JRnWoU7jK
rKjcKKGTWGPEmFJQ8Z1yIeAYQR06rRXzNmjbgAPpW37VxAOj0dZd00rfG6PzApBm
jna2Pl19v38z6UGfFiuIdy3QIGvDptZqz74ANLBW5FQi+Y7sAC9taAE2qIHHx9RM
BBz+CI58dBo40RvNoxyzPiSHK00Z6NtiZkdd6jLBXwUDfNhr3zeMJPWMx2IMBdFs
OfxE8e+j0WgUjsLRBw2J2xxDCrAhkN9LKRbIwsKot23bF6kMWrKgltcTycI5dQ3p
y2DvkMvVWD/+fCxDUI9awnsVfr9G3LNdyx+Squx9gU/BrUI0czUnlDzf8wj2P5jP
bL2GSO64MyLarxDQ6QhE4d25d8Qn3v7OFyF7uh+S/V5JpKHsDjtGekGxuJtfrVtH
nu+dVNj2zJRt/jQ/yUpHo4iksJMaLlQtg0HnRy7vH/+Sra8+0uOV88m7uvI1c7S+
W5Ct4K7bXP57v0JzgBy6KNolOFtKlR3eR38OM90mvEV6MOYR4HPzw4LFLgnf7YXi
YPeF75rJuFjgdo9FkCnZqTXwcW4y7gMwLDkj5mkgGY8tvA+C/2krbYB8KqQ+ztEW
23kKchW/CDI5hKIssNuE0PINBc0i+OG5wT63PobmUyuhS4tRfn2Y2n/LSuwo2qJs
qvU81mbtM+Rj7T/CYqtCBZ8+7unMu6FTfaM0HLV8g3Ziy1Rw57z1zyqZfF3ZbQQI
i6WVlGdLrM1NmQbz6JGftFAWKy26aTVNPV9F/Sn26m7mpfRQnQqOKBuw3AYwC2X3
gVFetRqDdk2LaP/4O893D6XphJp79D/FPDLVRQahHkmT2/24Xa9k8r4lp+BmTRGe
7KXBtnwi7x26lR+y7fDHOOduEPpvNEDoIYYA9iDw7PIvpbLs+fp0BYlgS4sXZIz+
L0Bsn6wh+JcKrebD6NdpCXToh2QKLa+HDP4p2YB2IAv0WrH/Az2BCk+g9pfepH+e
F6uzg9mtAkQZajHRomManjsbp73eVaVu814kGv3+lmgLtMpvoQu+fNJHUQTWZw35
ZtacO937lFcPVb4NNFJEJ+3DGwcosW/oASLF/B2BKbV98r4rv4ZMUtH6QLjcZ0ve
frfDj9Kgb4X2xzA9NWUvOCTfYwqGCiQ2Hm3jORSJ6b83X92+o8DzGE8P+pbpTFaE
I6TiKY1JBeYLpM7rFlkVKrFsLclvmhFeid/gkOdOVBEABBONW52esRY0qqmcMpiZ
4WmvwanFInP7shBPKm0MnMjG3HSEmuaAW/onPR+8I1QfFp6cTgN8oP9ET7Ko9ET8
vzS0xWa0OFfNZWlwE6jzWyxdfKNKYhaueWWota5eGWhtpHXZEmkhiglwR2MZttZJ
5yYOtR3TOkpKgTNF9hE+8f/v1GhX+zuUE/nqVq2EtXTSZd9sqF/f6WiLTbb8xnzd
VMY68lY86jq1ksHv9Se+HM5xyCGRr/sJVos52lRcvhtS6T/VA8B2xZYDSRNCUf9Z
Swj18S+C/KoRCyengBjLRS1DsnJYdi8SY3IT2Zzp+e2Ltgxf/f6z+NoXO/CCPSZt
sTERyyfTDr4r7X6cCxSzXdTVkGCq074u+66iYbnTcWGFkOePoOCbdFrJMA2/h9+w
Z8luCZ7Y5H1CEm1mNtbiFoJjnRYj7detLyBnGxd/vp+iFwI/Ja7on5mXaCOpd+Go
whRb/ViSFIqgUuFAkGcGbkcZll0xgIkZf883Kb7RTcFiZWAm5g3SAQq2S9QRcfkl
MEyuwjGuI6kYCgJyePTn3298Aar/BJpSdEFXw7qfwx3RsQXoFwYKgBHsqgCa/q9V
VkceJu+ofAGKEaCnL4BsSZjiGxILjdNTzhg7gU94QEzNl0CkuPawxus66vCl5O/b
SwQY/IvtvNQR0zTft9NiVYeiPMsNl6pkHuJZV/Bnn4RYRTz1Ty81aaEoC5fflg0E
IKwU6TCwf6UlldkfGkihV2etuYqDLSa/+gl2A0JbvpQm+yIkQ1Zs2a/ePKMqeELU
Auxc/P5Tnuge5WvOlXzSoHATlpu8dpd8PnMsFEDy85YZ/bwvf6ldGeRiXhnI3COi
VHyJzSGR+awTZUIzILbXZ7tiooQEaOVUpUPqcx2H2hkj+Hf8gJXt3RKvl9NOyIEl
dVGZJHPu4U9cP9RSnV41E/v2imOv8Id7UYz2M0WkmrPPvqVc1Mb0hFP8kE8OZG+D
Qm2Xhy/46/LV/TF3BIIDJdXF9lShnVDSm7oZb4sZJ3YfShOdlDTIQjY7kMNbQdXN
uGlWtOMq6JdYXgzlmtWZK6CiEnsZVzTe4IfNtl37g9tbjsrTs2QII30pTVGhsOzW
1wgKlkEzjlzykV3rRda+Ds0ZVPPKJX77UUxRUK3w/mIGXresAV/tx/OGGB7NRRQI
KDY0Qz1iiLt9QnqxwMSSkz9CI2Ak8ODp1MrWdGWSFM1Pf1Tpid5Vpng9hfOK3IfN
LGFPWz7UnvenDh4Rpuivb2SHQTRNCmeP5HBYugc/OntjvAqqb62igOzN81vvLGFj
2p/GCnOeScL4BZxLOMj9x7A6G9/HmUT8bFPbY9rnA5u1+RkAVY1FpbOLh2DLAa5R
+zqZ0S0ZzrMK7Bfs2UlJ6x3oJyVqesZ1g7HA4AtIvslJiURu5RyQGAvfrau4zKnR
d/Nlx5g9HNoDcOCMDZtBovF419mknGMUi24MPPb7wOjMRZb9hJIxOYYkPSd7H0KW
L4u2rqTp0yYSAS/yETGxgnHyhyGHeCwamhsSWMw4EYjrEz5avKk+JrqV3HTmOObC
042nmfdLf47/LYsdHhZPBvgRp/E0mxZbsehmaHMkk5x05w+/GOKLqiCPQQUF7EiJ
+VzjrJvmYNXyaiaB9ZtLbc+3TO9WWPjqD/ZUAG99/3ZvbZlZ08I+9OkjlVP/d43b
FCtj/EleYeXiHjztd9X3MEg3i1Aqr/uD04zAqJasakec+y0S3gQ8x3IkFgrO8Hu2
unLIAm06ohy1bNFNdPmmC8mr2DmA+FAOPSRUJgPARTUBoq2SvGNcA9Mq1jTLHsHs
0wRe7KEkHE7Dy2NstGlyS86qnbPln5+hgYdzfMufQ3ktuNYz2L0j6TaJJBsWvVJ/
2e693/Uy7T56yqob8t6WSTn+3NYmX8FV6vLmzyQyvpSf3LNX5ol9I+zRix3nDoQI
umtQ4QmYg4LtGH+E98VE4H2QlUsRWN9iWDW1PxnxTMB0Vm0aaKLy2ahisebza74Y
Re0mHnv6UCA2QquXDUKT39njof0ykbGpXmiJwUdhNOw2BDLeVUTdvDdftjN9Bk0R
elNdBWDxmNPkZ8NzjM+JGMqFd8ARYdRofPp4ynutDFHn64aKh+IXLcb8z2XCCEjA
S86QmCBBIGT8d0z+QqXqqN6rJTzqn1LIgJpbnUfOfCef0BM6RRzLR57hK4sKuZuM
OmSH0rPReh3PIBJrRBxzc6hBx42NBI21n1IcvSy9PlxCwdD2rLyuFaoNJ+QI+G0V
otT8wm86K3NPeqQjJhX/50jg58blPIr6qQdfOROmJvSDgQfdpgCKi83aKz6gEdGP
Yj18bLEd9nVtJnXhop0na8GGxkbrHDXHzl77cJ1mpW0eI91Td0oFEKi/TtkG8gWV
RR90Qhp692oSsmddQnp/mBo66rkkHJGT+ak3hXI8ISElf8G9AR4cvm6IR4MuOrkA
bVrcqt4Sa73Z8nM2xBGeLb/eHz0L/XmgDTSseIP0+/jE9tDVqNpvEXKKGf8rDnyp
Q073Da9lY7add9NqJZPD884cbo5TWwB/bpgKx8SVHPmh7Dy49kCkUfz539nCa7xP
qvK3X2uLwAhtBuItAqPM0iLrh9hUPPL7CXZUJRV9ZziVVdXAcSJENWP0e2jA8hJI
7dxPwAhvo0KWb8aP7MC8wrf7xt1WwYNc3IOoEKYh5y2Y6NeNaqvLvYxYoXEtekYs
JOAA3hNBeHR4M/BU7FiELvMux0O1wfeyig1uK7t6pAN786ghsyKF5qZbSyK8n1T+
FvltyvnlSfjwK+pwyiYw8GJbs/XtfH5BJ0UThPWc8HSUcOjeau3OekoCr/oq721O
kYV0WCaQQOoBYg756uOf7twz9DiA+ru/OVWeA7cMXIHc6c38GwlRgsboir+uL7m3
xqXC7eaAdAbPALXKCy1dWPcoJKg8xug8b12Jczp5Mw/92gbfrR+4C3Z6yGIzIJmX
kWnjgvSHbFnxe50ZyRYUE2WYZNj71+ZxAQAuPnXHk8TX7BMI/LHQyQbAc3K7BZpF
UlGmpUqIGjfQIXFJ432ogeXJ2jbodKxd4LnzmYcT7RxXAJvvcYfZ3j0w7UEv/YvD
+/Z3gRu0RqgCZIDKVGtqOeVU3U9ulEk+nrKSsbxcamfL74aX4R0b461tS0Vxikhv
uWkkzlcJLeA5aFqGXEW/2mOJ6Wwic3NnL1j1BdXJuYTip7iaWqTH9vqjL0km4u2/
630O4eQLcjtU2y/em9r50HZMi4Rb8RYLoRzIj7nn5/GOz8ig3NXm30yOszi/UEdo
MTvP5b4Y85wZiidFahz84sqkrANyGGwp+7fqTrrFuf/FOUYkpUEYCh39eX0O6KwX
2KE3+D9yKPQNawqXPJCQzR6a8IvC/h4HzsHDEKGwbtWOqfegUFSjVGvvIJLS94rE
u9W4X+zJxCT12uYyyM65zm0961zKtGNzKs7iy9PVlk2JP5IGlCI480SPIERtBopt
6dnZKpAEbgBupGQymR+7Lz1BWNDO8mpZxoN0lfbq2ssVaeVWUzUwb4XuCwJRMygV
Dr0M9T5A7yaUeg0dpunrEbJYWEAkeugmnk1cWBfgmbegxxg5W9uckrx6E/Im2RHD
Y+2B8BrB1jkxZo7oOBwif2aIIHza9womZI+5eo3+oaK6BB9DjbC5OcuiUSL5Clch
b8qI5w5PRr5eiI9cr+2l7BrjU55LGH+MiTzE2Des+dCc8nPKZqu8k1/qSMdBYDS2
T1HXNjmj5/DrWEvU6Q0XkrPw8VqYV9BjWqj/3Fk0H90CIMzQcFLymEPQSuTHegoR
HYhPK2AexyCbEpjDw8bCVGc/Y+iptljJlhW2XNbddAZZYCNpxZJNk1yIneWdH2Eb
lqejk8MIM5/32ZXXg7D9MCMx4hJ/8V7hPfEDC+NJs6RkjMFJDq4RrhlfolyUfTwB
NmxAl0gxLpbvVeDRmAPNfXGfquw0KQwmBMqobrGXDeojms9QD9MIu7mfjxoFJk1w
Tc+VHaV9OzPXUgy4Y6FZkf4Qh01AnyYKM7dGNiSXOelHVkS1dylfOTQgmeWq4sar
TReKPHnvheLXsHCvbOOvr5MvbiYF+W2ZAC25cIC0MvmCgd1qMwhY/pd6H7XHQ3xD
La9dR9i/w6zt0pJi2vcJfhWuBDRtsQPbiQMq5+ChXGiUwMkwogGeuKEVXdjIZI5F
IBAp60qRc2ICmswuc1XVlY1tFbtkCNpPbYaL+zMG/fV+NC4iSF6nE+pr9q+A4ZyZ
cnVHGyQV96bDLigsTYY2H1xUY4eWwsjzIs/AS+Hmoi4p97r5BqlCjaH5PvhJOtUP
4Of6ut0dJ9OcLSWiFoYYK+mx+ZjpvQEVU32EYXyu35E+HnwOLdj+ylaLzHeS9m5t
+8pXNERrrK5NHwPzYRfAdEAW+xt//jH6Knst92FeCWtpSEOIW4sDnsnB5nCpjRFa
pDy1umRcWZFwXzAz9X5Lr2MNkF0j/Sig5zz8D9uHMhJANTr+HORI3NUjOjwgeqWM
dlFLBLa0m1p+mJxLm6kBmALDmQJBJsuQmBlR+aAcUFq7NpjB2uy+6IeRt4+MKdya
Q4w+gtE9GK6C9rfeiY5UmxG1jh2zFjrbI2spTWNis2iTz/1SZVfVocQPx83cPTfi
E198850g8wehKFm1gFyQxWmh1cl1CoEZY9SPXR5sQpPc4hdO/slR0JWu/te9ydVC
o0yMOvS7KqhE+MGikP5QMNzaqi2JJ+B30LYkyJR1fSJvd/tF0tGgExjdz2+lGjhj
k44OYDkPl5FJw6tiNw9zNBxu6HWKIW+Go+tkciREzwNJPKLfUsAOHyhjvGejFU0o
q3+RNpw7Z9kHwzsXZrbmNLV74lzzjDhGF5XPWOd8YwvuORYRocwAf5kvmR0dds/J
I23xsAly+CVX/3PHX/JMCSd4X5Y2iDVh461O8XqCvX9f471JtWEwtrDn7Lho5YLF
dkiYycZDih4tmL/ripQa1dw6WOC2NZ+6iTXYuXXr68wqc6ozK0l4rlwrUgBy9NBU
rP+R1mQKERiQv6ySHHhnXENdE1PuFCBXwvFj7xWrTXsxtWmhqbolLb+jUB3nmcFb
RqCRDgNtiGZe84D1s0mc4KGx6i1h2yChgzS8s50VqdJKBZdGLa4jmCh04eZpchke
dZMTi/v3fc36OYosz7Ot8byNIhw75Dm+bbuxr+JQo7T5D3xGKbE7Umfs46/+WoPt
yK2MqHMo+YY8SUuz/5+i6Mg5qDDX97F36mSoM7Wc7XTtc0K3sLi/3AYrp+pcRSl7
8s22gGt9D/nKQLystCqBFaqAPTumC2wlQFFwAiX9Yb1Ol4v+Wfdu1C06JSBZ9RA4
+90q9uxfQTUtz2AUxegICBqhvqW7Mj4JNXLZsbzvwhM7HkOY49ygtOPjY1Caxx/f
GVStmFiz08Ti8NwVmIY2w6av7RdetvIK0WA2chhtGrBmO8CZ8CN8ALrqHKHBMbrQ
+ufvuM8CuS7JZ0pds43kFlYoX8s6jnCQJtqcF4yDmVJy1aoAYWnHwBAykrVqqH0P
vCi9eg1yKkiAuD59q/UFME4EowJk2KLrd55Gw+yhdMA7DipkH0SQYcJDuXs4woOq
90kAH14N87IYYY/iqaLv1bW+GeO6Nb0iwlzZCqmXHnQBjJ5GQHcTxvbzIWjipB/K
tPkKpnDn06JoVn9wgEJYSNod17n0XdZzuwT+RTV/UlMHT6oqNowbcAsLzhnBtBHg
I6LqUsvEimlVKtt1r1a88Z/6aasWIw+DaCaNpHgsdT1xHj2obiwTIK1D2PAX/MZy
Qvi1L9jNlyaxJtvtjcbR+dBDs/rnCvTNf8qA2Eb6c/QwUkQqrpFVSwaJgSDLzlId
T6o+5fTHFOju4upzNvc2P/Wys5IEl1VmyZkjdTRKF03dZvrulM8+GP1VL721N2k5
yJDH3Llh0zsIOYxGsxQgD4sOxlBaG+3r5rVA7dFMafbO+ERIIsLbqL9HmLwQCIt/
DqEvALJA71ZV7QHUXb2Ph6QpKGmBWEr/IjoiW4wQYOKAcfBFlN82qNoqeRQkkYIH
JOulk2oS1Jg5gfPSo4/VGyhmMfPdH6zyiDPEX3B8csuKluOcdlSu9u3tsb7Bg6bW
8mtDPwhChKdCaKxYPKFM4ywW1g4t0Q5+pw96RzdvDkNi7GsrE9Din5wwH85ybYyn
t7G0SpaSh6jUESMEaSjfdpvPFYA3I3OWqIqMK3aCv/TRFQMPGCUcCaknfhF+tB+2
ZrT1tIRMQjL6eLE40EgapzT+Lof5DbRZZxJNrCRh92Iwwpelp139FY6KiEuJoOGa
pBdrTLgONHGz64HTfEhHLyYZZI3IktKoXxIwf7Bi6qx1MEuKgbif8pWURN0zN4h1
q99OUACYNxlpr0cgQAg7NZJeEMfoQohoODkOBO+4i3xOsE9BbyhrQNQK5Szlxm1f
l+aZdFeEvsjR3WM4OiMpdRqZpoLepDb3NXH+ugj+GMG0UDLUmFZxqwL79hxme0VI
USGAuLcAFPqZP8wEWPTrWWHora4Le9toi15BSYQ1Eikt8C6Lrz2NlYdWtxYeIQQS
q+V7S2mYrmhumH9ak0jggfNfiZV7fcQpcj1YIp2ZnLY/JQ5jeA7cEPsCStK0sggu
WYiDplmglbrLZ5OjM/YuZF+eRoS1pXgINBkyVH+4wdsDmthcPVvjtMqRvHm3saBs
t9K1hJl2hBBGkxckaVp1RW0fvOlWrXF5Vsqi81sGmz9rGgPd1PIF8laxmPkYDbdS
Q1FhYP9u/EFXvPhXe7XVfSNvAjB/6/xJN2+8bHNCXSAcXjLa0M0AScXxkEuH5x8W
fjmqrKjUz0mLRWpPxm1NokOFMB1fdOAoznS0/vuawY4T9iMcntAJ5m+cB53iYIKe
H6gUed66h7QhZRMkFl6OWSO4yMSf59avbYJdfVZ+yRGWuMcGbv42brGw2QuhA5eR
i7iockMvwudmMm9nHXhQsl97ADb07abOLSpJx5GNkJ2X5RMh3VReHSJ2HLT/COkz
Vv/k2qQoef7XO9oJ8SVWB2QMEELNntQOOj+9U6aAAAyXNZ3E4ouUINqVR4Xit06J
4fDDsAZ9mgCozjZhzJ3j73WJKbdtZ58NURhahC/TOaQwtp37sr26qxKqE4y4oPLK
koGZzWT6RMAkLRbS/3toONiAaKDhKHqLgtdOJWjQn93sFwPSuMxbMapJLMTBq600
oGlHHbB7MJw1U/3LCp89C4HiLXoo2EPEwGItuEqJ/FQq/Q00xSwtegZIrOWrfJhY
BlEKuF9V3luzoyePldwBUywklPhx9ge6cGkc+4F6ncjTlreTzkKRs+SDDfo0YlqM
ROPefMJl4WokwUSlQl6cI3HznQUy+2Rmk836NcQIkQLFVLKe5Iz9w8fnTn8eIunm
zd1E4KTkRvYo0+hnv3Sf1kyxhjVQqmkJaDAohUnjMiAJp5pa2Bfocox+OrONZkpz
7Ugr3XuqqH+tjocH+J4MelmNV6HSLSaX5We/OTCwpjWgv8vd/6sg6YAkbLRJ2kvE
IeDJKLsFFq4nIEHiqFqGkUtDIJq0gY810QPhoYGWYmNTS4D72FAXZ6HgYIidMin/
T7HcZwhBQzn+seI4FMVpnDfKn77WTpRVVA/jTtTlFMVJYipJaoM4n7BQEx3T5YTq
3DKaTSos6Hs5EgFixfGztMRttFrXDokxwKTL+/RAZGQ9sxjTzjEOn/idylvEe/7n
Y24ykxJrhXAySM6mku/GuFDu7henK1iPWCwHAL3WKW9QkrM2Q8ud6PH/r3Hvd5LC
luFGqlzTfMN8X/ILk6weYWba8VFjGcIcE8qr4h7zKRfd3P36WUc4w61ws5Buo+jQ
8BV04vgSciBt9xNwEhPyqGdjDk8bHrAsejgMYoDZ1eNDQVRigUNFqYrla2BvGX4T
aclc9yiGYBhvJCq1HYVv7M7V7LoP/23TAcXuxZXDcKxAU+AdaTaLmEwppd/gDwnS
fc4n90L7hIJ0s9DeX4ncxX1lnXrYrpqNgDQkrret+eQw/UQmwTrLSYxZ3EC336GJ
xUneVBMrkLXDFHkpw/djYvkYhy/07MBnoJJJ+sJRdzzEs5VINsMbsjdNuQL54Q3H
kI5RiRkHwMSVDP45c5ZbqWAcbAA0ITOpAEPYoUInWYN7BRxgtDOpClRCzFJ43JMy
MLTsvKd4yR78v59Tjm2qEjpXQF9KgWDjDYzK+IucdzDsOS7in+i3oCu6H5kZe5XT
UEIH9kLjjVkp9WpR2pONIxG0DZ7SRNhwNBAm/rDSGpiDQaIPC7SVzk7WZAK21bU8
IJAVf0eusfWw8Ylaxnnpe8IkLcK+vYxH4B0Lwn+QjkoG45f2L6//GFJkP6qzOWk5
s6FL/bt4eUWj+bzsNGBoCCsYzrH8nkjXaCgd/woXkY06NPz9iu4xVWE4mT4UIpXb
XXw3aNwVPd7hF9BeK/yqObQvWcqJ7O6CH7AVb03fw1vFqKJkPRp2i5xO1qhSUEfo
JRG8E0l7CfzD6bYuTTT0SdS7fxmZqTXiQq5OvjbcxQHNoulFlRIxA3esGDKzeP2z
F69rQbyN0wNslpM9BWSfJMI4tUtxXD4gi+11hnaWNcgAJVcajdJUputbhrJZuy/U
3H9btRjKYel3w1K83KmTaRsSYlOe76rMIx5K8dV/wmshxYXnbs5/RnlsnQTiQGqf
HEs9/SOVvDgM8U5Q38eP3OJr932JSrxfyyupKnI58IEh+OizxcXQB3dyiXHaLAw1
hXh9MB1IP5rxLlh/cVxsBrGulXR9YZ5RUFMnBb7JJ+cHA4w/CAKOllGhKv9VNDem
gwDd7hyUO6pKUrq1LfS7tnR23Byy7AO9u9SWgsEsM3jNuU8oXJVAq5oMgp2ZoSKw
xcYhoUel3K5oDLwDBHAReSZrIloPSrBIDQzZI0EZqBkgvGJ6d8GF2pnl1b44sE/U
C3I39h8gIBcRezcrhVj40xM2l6R1SpagR5LvSLndGxC6mSrKF16maJdD/rZdnKG5
BpdaVTz8UHj91RTbhgUXh7Fz3Vi1jJnJbVxPBSpe4n7nHcVrDcNGwzFXskTUS4JE
auknfmkmETeKSZVeksX4ncodlYNZ2YxXROlF0sZsrDUoubbIb6OXtj4Nc5Z/K5Gf
GwCeqkfJ3yR0Bn0Ee1vV/iJ1N5kRaF+tauZxOj8oToa7ixzxpNz8Y9mfs+qKL41J
kzDAEFkPoWNq0q0HddF/9yDrZ9d+kK9f5zt7GlsA8XbpGbJdPe5GVEbyGWpdkq+X
bFV/vALt7FJ8gCfQuSNXub41XBpIpD2iqxNziKu2Ulo4mJk1ulNezMbPW/VD0FgC
qq6kKsNexbngTuzjushq2N6U9yUlRAeOIpqZvu5jRiRaJUXBj81L/wBUzZSEuXeU
I+Uypvk/E1BzBArsy7lkKw/mheMupXuxEQqpCcEvEmH9cuaId5GbCLwkMT9gn7QU
Y6z8K2j92KkHUXCBvXi/K+WkW0p821uflb8HPfCCCCnnHmaLmqB05SONlB7/qmGB
k2SONsCf2HxzIfc1+X3klC5BVV0GnBEwy8/dzl9KEMZnVXWyjJG9qe6YFLSxDFs+
rl1bM0WtjzY0JJgwVwgZJC3iZKHTrYmjOed0sp8VZO6PKzQpQ27EIA/dFRkGnSuI
xb2LZn8KOySqPuyGTORZzitW600osSdevmCLVahtaVTdWYSWRYn3exlEPMi9etgJ
PxpfCCs4iZ2S0XmyBlnJBZ8rIWkVE4e2K5FQKxd7kXaSJ8aYvVqa7hswY1wMW58x
iVGUFpFnQR7qTzvWfTJLCZnrmiXj7RgcM7q72xCXUUyicJ30UQhJ0meuiATIhg08
EFyDwq8MrPoiNx3GQnn/d08fRWWZTQ4iRcwNwCTdgy7T3/Zfl3mKFcNlFmgs05ar
IG99PUMw4f3hDLQe+HBF5ZGVZYmo9PD6q39YRTyC70yhiz/lDCEUtHS0y1QZ/u6E
sSmiCUv0gZCOI9AF90N07z4Ef3nW1aPD3Zoc1lEQ6DPusjCwBZsOe3JH+XFxgZnY
iROyOqv9UUie50wiSleriM5hSGyF6JJDKP7DsnNcsY3OtsRyB3lZb6KWuectGLZT
uIk6uml/HfhO0MmCsVwrdb0IS42QQFWlvKkijwJms9XWXUW8VPNFrZUxwoh3x1mV
2+3bzfnQB0+b9HhQEiQkzh4y6J6d3kWiB+r+tmH1+E4oRO5R62hHMIl9Ey0X06/s
nXqPELJ3g4WOMtrKuQofGVnSi76G3/wnJiGQT3Z0wX2xTbfJKPtCGPOBF/FGJI6e
XOpt66AKFfvIKNvKM1R7GgKGk7NN4BVnEJuIAVN/YHdFHjppnI0aC4uT7TNS0VgJ
SMfgjDw2lvHAaW57MMULu0hnRflX+sC31D3IHhEYePZT0vOBnefVJkvmsKN7MBNO
ONy5XfEMKHvl34DMu0yJzAdqiRJr36KnqZPVGwYcph0pz3djcdEjUim7ckVE/N/P
1HbaaX+B9ztemXEo0Wn6pvGzX01BCF2BrReeR3G652e54j4uFoLGGx9kmZKnui5a
gUIQh4dnUspPcq+PeBvSLXqJvBNS22p3L4zkTtiN+cfNJAIanbipaQulnW2V2lYT
WqEsvz7tm8QfM/GKLEP1YCM7ZBHi303BRhxC/RELhiQrQJqkQt5o5onQe1mz4LPA
GLV126gT7nzJfwIFfiBj1te9l72HyyHMJsFcKQ19kNMk+LoSERE2Mb6c4Zi4XYkW
MLxLkXYfJhkOuAurgUHPjAbLFqUFaw+AUA6i7cUM8Gnd1HuXNI20VI50/Q0ELzX9
vpFdeyQ0fdDr2SOSSgI7yGvS8SFc8cXVDtb456iKy5uXFR5LQijDWgv50MS53XEi
QNoI0t32ngwGcPYXymZQJBoFx1S4W+z9VOuqLNgwa2UV285WJfIt8gqSoLYwZqgp
zVjluGVRemt4toRsZf5Zn81DbCnytEI96qfrHUCulU+hIUhbD9wyVUcIYO9C59Hk
KkSWSnQbBXNnpCMeeqVMOvY9CKPx7QSnvT3VNzVBdBRJvZ0rrC6Z1vxJMk4WhoQY
xAzCoUY5KB2ymEFZ2Zt6uz3rbtDmQzeMxUlBc1f+NuqCRZHC7HlAaSNCr9IHaGzl
KGaeCyOk9lz4ZvFB/zyHP5M3FY8aQENAq5HbS7AEsltjW3GZtQHxRbg+x7/Zl71c
3ceJT2W33SOSuq4eLmUgWT74BEIsvBW7x9ZdxpejmIn2WmXQ5KwJ6/RRCASxsEk5
8H2yvl3BBO7J17FnJukmoOz9qE9BLIa7VnNDqLLW4IURSwM+XaHIJLLJy7zWYV+R
PaMrq0Uve7XEMfoIwB5xYAeXFwxvQr/vNsiawG4RoPyVdWiUByONBnWFtGR7JcTN
NQG6+x2+vv9YU9KrmclahTkaJ2oOH3r0IwfBiUEYtAuHm432CSHWQ89xaW3RaZCI
dsmeDKbe60VAofbLjOKyfCYAzDR/FzFf3uOb2kZJivL5k3BYKN2czRI0NG/+4Olf
n2IvizS6TmHgRh++5n7NgR3U2Z6+/4CBR+q6BDMRKl0MmdHgJwRMlG3gia7f2n/b
6ht52Z7Oa8s44mt9BlzOcoUOd/bXhgraMdkgBvKD4AmqloBojI+Ozr2oA3AOuLo7
gZq2e2cWj9CprXr1156uyT1QHZThucIihI2Akr2PnVcapjHiCfLfe73+oEOR0kg+
SHFANUk9i6sZuALFB8XcOh96C1I7FLF65WVfsTwZ9a78yKtLIdJIED7L8dC3hbyX
TqM7JpsXy4ylTt6NgaiYMW9uKYj6WNNeDWpbIonBGlYmNCessNAXIqXFuozQQdBE
JAunfwp7m1qWTbcTJGHgaZu3GNee3kNtGujPbyfulcMVKWbSPhOXBdKlCBcRoS2/
OJkzbaB/ysN1cesBROZy5aewoH8w5XpHQr89qecczmX386gN3vMYohaPvPewT2HJ
aUdSj1DcK23WjMKlee5MgIZyKduLPNcB8DAOz5FSEJGv+jpJZAV+vECFpfyPSb7U
HE2eEYBd+tpDNZz6XOkm4j5Tfvx4lfkjyxoEfT3gxk0dLW8VsGmwB00aWQKRYoeG
96hz45m0U5ekJWTH7nJSTQEWG4zfWbjnsB7nZmcU62O4czGPaCW3SwQeWw8k0Ghe
0qNAIFy1VqT7mbeC60mboFieuaq0tp4EhYvaop48wzL7PTVQqBG64EXI9h3hRTHB
cHMlO0p/RpcPMS5Q6P2LLtnfxfRJ2tLoYNxyQST44NRToOndCLsbEpMOh8kQ+q03
H4jkQ+L7yLpvvts9lrM+9S1TjYvyM5rpDuKgM7qqvNo7+/fyvQG0/QY/WnybLRb9
ftkaial5ZKSOEvNI66Sj8z6FirZ+9QkilyFtORbyisSX6uAvjnSDSb944CjjRV6E
YYORCbckoeA2HI8SDf4cHUT6Q7Ba5extHGyWPNwYjlth4n9m+v9VPJlvd5kRvlGu
bwOIJ91iRjSbBOqzCoi7tyCEImtkwX3UN4NFLjeg/Kv/wBBQN0J0FyQIjJ8gsCnX
XIzYY/odM3LuhcpuzIb/KNUQP/9GRQIB2BGxpkFLvsVayUD+6X/2ESKJbIi5Aq08
W8Eoipj0zY7e/RVig3Tjm5wefelkO1YFqR0ZSZJDEdtShJAWe3JoU2yf9eE4xAIs
/54GJ33J9Uw4fE61Bw0qVAXUq+8IEUiSyv2a02amPh//sejBj45k0RZU8Arlb0aM
xKt6Ln+S0ygOVh+p3/521y4iWf6gjQ3YqAkMucRqKcShJ+yONoK7PDSw7d6VvYfy
XfcYo44ICFd5UsXkBj3lPkwktI5qwJyNVhZkzj3yMeq04ju5QoIvTk1Gk/YCd9F9
fTW9azTYFUHaQlX7nds3YXwbTk6ajetJ2kcrxj8JOW8pXeBKUGYUX7LisZ3iAOi8
Wwk2JU7Ccvoby0kKwarVroPmkk3qc2kMDcdHa8kX9AbgBHh9k6mWPy/HiBt9gX4E
MTyAND7NQnImHyWLusDWmEk4mAMcz6c1hUMPz5YRixpSDu28OLPrSD2Tzw9RDr1z
pBCQ06vchFdCfAhn+541ddHolYY7E5mA2YfuegxDPEKgPR6WSx6TtyNW8bQ1zJZN
RzGs1WSWZrc9bxEWbXlw7D/UaJuZ1FWzkHIVaVDvOt/vvSGHyYOo4piHVawwrxxG
xs3QsF6V5p7i45ovFJmzKQKNrF5ppmNnJxI4TKloYvuATs4zIVSnZMM//Os1/pYB
QvZuXMwb83Pz+tAHhXrnZ3U+Y7ZYijXNoewDLkkvYcRt/oJISNVb2jOj+T6pbVym
+TuUTwFdnkrzOM6RoMEO8ioK9gBo7/3aCweWi8sEPsY5kRHI2QoA8RlcLUCi1D6f
2bPDahRiuGbS8yyhW63GJSpfQcMPSXiMWNcQsr64Mk9HZSlNRSjLE45kx7bIRHy/
rMf/yARnZxx5ql4FAPfxhFqGOw1u6sLQHgRgkrM+KeXaHlftW6R9Gk+FQukRv2ab
cTq1fVrESc0M3R+Eq0rr8CNcy7I7cM7eZXv6AcIBJ5qTcIJBD5lXUFkEMBF8DIyC
QVp1ORIz8VTUKE7j8HvImv+9H4Wp92xoGjgs+TuOakk+AfmiJ06ompe3DLohg++u
hh5wXwYd7uvjmYBtHuZwrGPDC+oCYJD+g57EGGAC00SYnmyEzA2/DAJmsz78NfNI
8+UXxZF8iUhuNoR3xyPqzUG53Of1BRj/bgKMl7OwRdAq2ty+9AB7e84V6SC6jma7
RALNgrW8pzfALMTKRoaMWxi7GQlLo6Tt4xS2fBbhzFHrLSohGhKbGjIGh24xkkeY
`pragma protect end_protected
