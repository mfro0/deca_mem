// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:00 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tIZlTrkEC+20i57Y0j0g/wmKn+0NUTL5/4POBMv6KrltIV3otv9eolIyOVT+0GjT
k9qrNIW9yw/9WD1d8ZKAOYcd4K2TTBX3JK4xoqeGuRTG1BPqOGOuZvv1hL9etDGK
KmHhq6KdfV6Eb9WLxf8eV96F/AahMMMl/GOquMWsr18=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18864)
SZatMrsBAcRN4pP02MrEQs5x1/clq5lDYnlfcOdbECTorCFTZ66kr2Qj3iSvjMMA
5dlOoe5hmw9st2pW4avNQPGMf93Qys+wCvxSHTQjDuWlvLiU6+K2Yw0ZECDgC0Md
E7kryaaWI7UN+k1LdheBFCCPpRHKKSYqFgfS1fVw1b9oiOnnoGvuFTuzq4TbWpcB
j7PcExTGCuFyJHxiBDQMBav10H6uL0rWOLkO2NHChyss1U7WjCi33spVBfgm/nFF
4p7OkPXz9e9ybaUO6s4+uNl/GunAD3aqR2XsGWYkz0ogx1oB6M3rGa7/NylP9Kzu
MD8ejDET+vyJxAfIydfqN87awM24DblCPp6y4t28mo97spEbDvG9cgcZAkQKFZ2C
uR29RqKyqjdSmo6TjT8t69Oj1TEwY7DI6nWnF0FMynJtDcNuO7O6fJvcyhSZ7GWA
IQFL8jvEFQLB8qVqALt0k5uGZw2sYOsMzfLbF2H2+PdtfbZ1zEdKSO+IzRcMlUp3
og8/KfnpZCNE2wSD1T91YO+QO1LvJI7D416ZKty1kYuPiTtz15rdrO9ge2UQzsXg
hM9c49yWGH7/PZwDuAsVy5S1ioDw4cmPTIK9Ze3LI3WT7Nl571tuvCzX05HVOUHj
yIk+wQrnrV5jq0vlgwJK1BOre0irgDAG2DEIv8TEctjQ9PwRCrm8TMQa/T828F8F
waFDvmIfhcr/CDp4d0B4crxIv+gn2DQMq9ho6JvVCuleoT6IWV3ip6HTPV0z7ItZ
i5c2VoAf0OcsJ3j+AlEiD5jWJhgYwE01Cu61PBY12mcsnPLG57xoLe3961m1vlI6
RWFGX/Pzb+QseKefU8PrmthZbQXpggqPGpUPPrY4qo5hNZEdrM0tn6DAgmX42GlX
EguuRsa1tiu9gGw5zvNeReC20omQ2UVwTGMw7sy2D9VqHtE7csAlDCJEZlZBDIqg
0N05Jbvz42BlTUBGhfNLzrB6UgxkMmZO1jYqoQs7U9UVZA00BV/I10zCCqrDI/BT
5nSCC9oK8rWcnUFG4aEHDEa9N93qN4A1+51tMvE60cUSikmEwYViEmBPKp9v7fZa
LLDGoFzRuXfXk+kYzVj9MF9ivb0rXyJFbt+JzoYNcrDfI/2DpXOzaMGwPZIUFGEx
S3sfveOKV9GBNSvs9LKb3XbaBaVufHcKrRKO+AFOZa4SaCutMoUfaBu+vUu9bUWN
/xTIPPP/VHWwOQ5qHfyC2UcLXV7LUlVNCPYyqyqMfWYzJR4vBpG+fkweY5fzXdJX
iYenDF/d/ReRi4E/x8wuKQtffp8miLKD+S85QZKDJMonrWME2N+F/WBZ3eSEmbJy
/95alCRJhRspGKO9hxUfekWW/V6QxMvuyoMD4Yo2pPEB18rmjacGhNCwt30kMYe0
jacP3ZMa1uooLu1qjNocJWEyN07pTJOeoiqo+344BtSBMdHU0BUyJz0CFHY6MacJ
Hl7ZeKHal5sVql3okMRhNHV91tQRJmH79ZeuPQVl26XlLN/WDsETHTKEyAixw+A6
6dk9msw56YJJ0Q80E9EBdbLbSfFWZGx4xoBViQzFO8UmvzETqubvnn6NRbyV6suQ
4e2yYUgqn3v4W8PUY8/m7fbn6w8U0VpT/ARWPrO31aoaZUqVQYoakNiiAtWY2Omk
FRdVqbElDV3V2jr/mOWYccUJMK5DIWYw+TPNrDpV3rwX3eRSplfSpvzWwQPvHcd0
E6Qp8w/AtolTAK/sznQHhsHFfinrADPUqpwbJb487JLcg+qGy4EjMVQ5qOmh4w8Y
J/aRpuoYKZixondSojroGXS8G8CKLROeeDWmBmV4t/h3uSRqbpMTMvbIIdGQ/Z8+
8twVJYYLHgmmjf/NSKSU8Yhc6aBndBy6cGSevBX1iKaGPMqV1/6n9xIIRfwdV/On
1Czql22jjs9P3y9a6PsF3pnrNCN74UmBnvIcKXs4LOGsNIi9iusa9Diz4vz8jndu
9DQ7Wh9KK4GDbLyjBCb/Nlo5BXlRtQWAnidOqkdRrHKTZVVme00LCyIeAdY570z+
eMHw3h5KK792JRUmoC/CGNd3Ox3FijUm7aVmBeOyqbt/vhYxXWsEdnUywMweL8+W
7BkUN+b3PBPeMAbHhZ72MgDerCbYzUKP+RqA4LsQ6vcU1vNvOWHpkU8N0aoIM9OI
lzTrDXiWLZK+7qyT09hte0+REFumB1X5vUuqxr+Y6boiwfHcY6EDeXRrDiemyn94
gxuj3T07rumF2m5Q6vFHBrjv5NX9oV3N2v4izd5sapQLiXhRo9qO1rhbz4im3Ep5
LyX3m2wVxrXXKlNYIi08MRhQVErO7TwbTCD787FKZV11ig/BwPKHJOtAE5SN92WC
QccUDDkCafgdKsRAmz7a6m6MK6AR93onAbhVN9qbvQXyWCvYf0GDO6FFy5E64L/E
Q6ks1/eOf9rGQ6Q6+bhVGcMYRjjxZUp269cwY05UZ3X51hoeBXiixS57OBRZGDnC
re4P6nSeRYSC1kVz/fBvHS+22BpsXc79npUjzbOG564UJy/cmY4PEVoJV1LC4hg9
AJDwnF0A3T8YCzM0bKSSyL9F/TKTOa/Y+gBaTHr89N9lNNDUAoN0SzYj0wiiZs8M
xW/cvB4zcHRTXSqDlqfbSGmJz1hErfRbjOEP6AzWtAHS7TFWf3ZcKYgWl31Kv7OY
kIalhllGjzcG+DRwG6FwIBTTB9TsDYMCd+yyBaUefOy+HJ0D9qxDoATSscxBBw9N
hqdO97XsnRR//84Ud/uGKva/KLIJkjZwzOvr/yus2Qa4amty3RItm4GevbLEc6RN
L78he7p4jW4RunQ0MH6IQdtpNH3D1r2DulO0IcouMEkh/G6QQCVJshYnOMH+T/sz
Z1cfD2t2eTpGPiq+MAEuvEtbQup7Zg7B0FPwKRu6LMkpn2cGWuTfGuUW3VZRL2YH
LZvA1ViVW38YMuUViRV9CtcnURo8gXilrEv/NT4c96P73tsoux2W5ufu41+mXcGW
xYdt0JhCbx9NxsEri4i4qPFV47P2itinqVl2S73etW5FtieKJIsPSeuk5fNw4uEE
zVx4oQlxHgeO4g+lo8mm2O1q2O8GfsuW4Zt88YIFugQ8cCBu29/FkoDkZontum/e
mfg/0EpEAWq1xA4P7YgFG5NklcpTdFURt/EvmTn8fYbBIAbcuh7w8BiK3Ck9Bb/+
CdHX+7KHWPV8cgpIUFyMBRKDVowQoHplUzhkMJ1WJneuu/qjafF17Yew0nmrDU9n
sD7eb2YFEW6r3ES/Oq+Ry5rveOqqFKvS0YNWe0mg9bAylTnA6iWcg3McUbOwYG8d
vjCRoSdSi0qSDWq5m02aD8/RxzEm7WQilMeij8jcngZidIppxNBQHIYTOcILh7N2
FtSrrF/gNrRskLZoQLHXZxHXKmaohLRYo9Q5Qztza5XxqvJklu+cBOSi5yzjg0Hn
hCJtnfEyQP/pncwiDx0ilBldWqDithTlJqgKz445gEkzC6P0ivMjx/G7odEDstr0
QJW9kqHt/oESg81rH6OUMa4iRhF0wBGSVUsxED/TXZ00meF3e0RSINlm+q9r8Poo
G2HgFAeO6gcayhoytMHzz6fXJTqHGJ3ZqW4aUG9MFMiqPRfy0n1K41QkClRVZ/St
TO1tLalHjm8BKu8fW/pANllUL28J4M683HYfXAlFYE+Wc/lOGlFNKwwtXXXyTe2J
PdL9dy1Eyle0nvZxHyJUXofK5iRsGtvtk2fGQCvxFgrntF2JgffUn96Vrvj749qv
INA2JRPF1gtUEtSUo4tlElnzUUo9QkfZvEY74QP1xroqNt4DIFW0tZG28a4VBjde
OObBZAEH3lZQ6vNuwhZJu8U+WT4XYV6K26Dtk/+lyr3OEdb7f7t5JxI5YYa63Sj1
MW1pJ4x5H1RYg4bDG5Z8My6jCLiNVQRTrTxn4WqQNf87SdCjsGCwI/WGRawxcz8Z
lp5y6eFbHDwibQLjhUrwiiRYxzeFVv1mjXPyPUgG3aNSjUd+pJifOCNtZRR1vmXB
lBnop8p7bJWcM6VzR67I4/hvxO+Fwz6EVeG4RPn2iIugZdcwXZfLTr3mJUk0Pf36
HM3gBi1fLl/boUO5ewLw1oV0Lbztm2VNAeVVM5hOXeUlNzb7HQONQfceeT8ho1O9
DqUkO8bOWKlVJzPpPo9sqP7Kt16Qi+O2f2HigSWB2GA3g1R0sCkN4pVHhufFfqqC
GsQX8JhOuv18kAsFPTfbh2DafU4v/rv7vsKrC3SSRhDwa8Ry4mgqsx5+W3MheIAW
xbda4YMphujFWXdplk7qP5mSZB186vWOybNpm8pQ0irmyd01Y61RjUxnERo3Exbs
/eY7VLRC/Nqr9y5pvy5i+/BkX7So1GIGpGYkDaXTwEqv4b5yZkBBe0MLAKpK5Jzm
hS2q6qmcpryWAOrTG3Ta/E/ibsWExgdE54kU5sfGJ3tRpaBcQaMVlOe5tFSMGbOx
aA70sj5IzGNQvNvz5DI9Wj2ngPc8EYEObChcToeBMhioyPfFPWlHyYAOm8mdiLCL
eSiDC5FP0RY+RybfGMUYkQeW9cUcWkk7Ka/iugtwbVhL/m8qu9AmE26iD+Qw8PS6
eiwMS9TJGzG6y6K8jtthvFLQgFib2BmOLhStT3/wLMnUvx1RQf0utok7vAMaXViT
RDeWgCOm6Ft/Eu4leENAJUUIKsVWA0zfzYP7CFKqEF0/nOimX2pskd212or4zvTT
afQPRndnkl1Mfvurk6psUF9aOrd3O3VcufI+StcHXnDQa+jJf/Eq4XRAFaDVGbxf
HRi45yEfG3/rO/W0+KNZg6f6tsyQmhInDeg7KGV0KRTZj09jzqYWSVK57CF2f2Mx
NveTB3uRmmvSjcHFmfqvICyaVhX97ntWB4PkXiTG7RPYfOt+t7D7aA/H4yS+RWa1
qr8SpaGyO5d5fe5F5pPCM0Jt++4DzfpiIYwH3bVFHvZEPPP24l8FXarp+Icwd16r
o5qGH7tjr/VKiXKNW10dHX6FKPrzyvbsoumvV2e4rmbQu8Xu7vyvN1Sft8zfBQPN
t5SnFrw1NUwfxotpmWHs9YWJl4P0eU3yMHTW0CnDSd5cBn14JdASgK4G19fCcZHk
0BcDA4C+eZyBxbw19ccj6UJgrK7Njzp8mSdSREdxieMbjGqCeTh3dj/lcPYDq5+Z
qXORyO8z53rfsinFfSdFSbZR1zPDFDIGS0DEO0Oc1BsLTTx76I9XAVdNsYOeD+l5
lbuRp0I9r+quVPWT1/4EhDOG7acicn4QJPJUfve9pD54yr9v6kR3HaPs+0jCM0eQ
Kmyx8v21kzu0FYW1d64y8hgHqUIAQ3HlymDKoi9ltq1T3dmjsUpNatL6IPFYV43z
HPFx7mNylnYpDZUd1cirU9aIBc+FydZaXdQhz0KTunmbAny5+59J21/J3AeaJmPs
q7hpx2fc4wusDHLM02aFBBi49mgef7ClgJiJhXyQjH80aRCHUHSFdi5k6PlY5rO9
2bM4v6SiM5oyYiOjzaWH/qRD4X+BPPw4Hl8LUGrwDnlJDB4J/FzDuAETp/2xVL6s
l+EpD4JetS/RGtfm+nZlN+/FEi4gP8+HK0Ei/BK7VIwFj1gggWbWVyEb83fKgxsE
ZI224r0AGY99cjZFTIAcbtM9ZYVe6KGmEQYcfgwzHjY/G8FVmFF04qMn1w9RDKLs
wfSYuErJuQSzTvBnlZZqNYYP5fzon4zdGbpcfbVZ/NRnlrql/zOPCX21HPzdJhu6
b8WDiUrUmbOo7rUHDJPd8aKjxDwkLAwKfuZBkAbvUdzEHijYuVHRPrQSJ2GwC8xm
VseGAlNgK/PdiwfstcOEpjjL8CtV34pbNMw34mWh5RsP9KScew/QLXWpwS1jekMy
LcuGcMQ+y9XYXBVsacRWQHVlDODZ1INazgth/Ukxl7ahOXSoA4rucD4706vR30gM
sDxTkiTnYr78xp3+iSw9/9yPsLlko8bwSXJjctLdYl2C9orX8OTqgF817Tj9jAUW
RhySzvbHvxfxXUMzu5tJfSEEB3To/lYEXXJGNtLRvOfKeJhLlWbtAhUVGUJVtzhU
uxEe0nHt9l4h5aPzcnBFqZKrrSEiGltNq+eqyLXa6jWWfx/wXC+f3KSgOd+pwWwe
+CDcEkenci7WVCS1Ox+CfbovzJJqKIAIfDJlrtljyz4YYQRv3CX4zSl76DOD0kV2
9z6U9nA/WVTsJDyoyhO44ExgW+4nwDi788oLE9yxwLsVh3q701WApf5/Evu0DJJI
aFvmRmw/3bjXuSm9hHpBEqYoVXLFt+WLyVxgE253CLp2SvQ5tszpbfBKLBdHje7d
ZmU8wVhkXkUdNC4NbpQSiUeHTHpChV0RB4/Mz/LdB9SFKLgaJLKIWtFR/KSSDML+
SusAIVVZ2gGmacjS094SllZD+zydJ/7TD169LWfu7kzvYIJkRIVvJgzp0pVrGUgO
51B90j9oIRCfwwkanM28MY+A8bvYEFlVT1moQ9OTUfD7wPPmpb9fZZEQDcuScP8H
kKcfhgrm9BbHTMRCkkBDvIQ1tKJZr/w4Yy81icET8nGr4UxD3dDfCjEc6VTr8dh+
7YaDBqeXB9wpQuzqYynpqI0apkFzZgcqOl6lQR4L4pn6gmareHU3Udfp8t4OsUOd
TPePRIvTMorvlOrYS9b9DB9aNjeb3nTnuJ3hQi9OBSAZ6bnS9EkycGCMxjOb/XQ/
Jl8EMndUuhxaMsuiW58O1/dtkQoqoACoWQIAncn+ZIrH3E+qy5ubOe1EX24AQALd
kM1PjAhTa9LFeCinQF7kgVghQjEdKh1TOwk4ahNfA2KB7XFNZYuyVgRKRpng+SbZ
e3RL56zIrJeM3/7ZmgsEOogN379lK0gqFQHzp9O6D3Pb+GEZRfHZy+ZP1SOluQTj
2E+0d6ghxvRa4aRv/iJ+aHd+SkTYYrtm5b+zMp2fnn33dtOfJMC6HcaUy1/uXvHB
xi9uYPabDG97zL97wWqXQ2RkDVEHxldeixPUd9zXLtQJNLrZvjklNzaY2zaW6Ijf
1cKSnDj6eaZn5uSQ3cACxUA8ICBxErMBsp5IDSMYhXWLogmlkEMmtrUTp0h3nJWn
PB7UbMIOwHuxB2oJ83Ed0eH/wANPhzgQywpCeLt8ZOeLz8ec6RVpfp2DGwF3q9Om
arzfvt6pley/flWTVx9RKdW7mCDyy2oLIfoyE4ulFAmq//vLVWFXreMemovX1eNG
oc2X6vBa+GLJug6OnIgDK9LO/c55NpYskTi+Pt1jVorACBPWlgq764uqcHjDcPUE
kiHHxeLq1xNNggP69rezNeCqQ+I7issXni+FS8ZisVvppoqJKWPZ+ucOAr9C+1IL
q7mzus4ChLakunXR10rCRBgMQx5oD3T8QNfFfL8LszvtC2U9zjCm/IWanp9GXL5E
VsxAtEtQjRCtFBKWZxphsEzqTvhZfyMHNvH6n2gID572KSfalcx/4gh4PcM5P8/i
7qO69Fl9rOW6JmFacxCuM+CrBDcU4aWHKquU9bS0EkqYH8XYde6Pt1KHU63KYRZp
SnZTS5D3VQ9R1NbLDGwpjMsvyTuIteWebkbaVfYHpwF+488DV3RN9fgEVwxd2Yq1
E1E/EL1UWfIvkkwShKtIZCOSeUAC9Z89xSSLFPl4+cZeOsw9SDcwLBTbYDDjx9mg
+9axywclKiIhkqs//nwCKRqMNzo92wSQV7dha0i3tBa0kvZyUYWy0l4DUd5Cc8mF
gPrqo4MkdIt+AQ5/2v8Ihm/FxhyeOSW/ude9GOoALH1K/5HDsUw4F8YHnqTWJfZP
Uq98TU/G8nI274Ns2H/CuwqBKnbbWXyuTguHhhBUSA5z9twnKBHB4pkhPzUldijb
/PXynXGSg9CK0sLYLcHYCnf4rLiE8XLesy+CPfzN/gda4qAXoMysC0DewrnGhtnc
snRjoHC7f3V+p3/D5A4WYJB1dCKlPJv7VaxKfnOdfKjGEGfEozVnEyCQmADFNCKz
WNomknRsii2vlhjVzET1FHx85QM4HD5jtn3UbctAIl2uTgp+okJAqKBIl2zcdWgC
3Q1BuM/EFDGV+imVEmxAae/44h5gVbFSsirLpsgxCjGW48Vwfqg7dy0zo4cnZkO2
DThoFY68lzsUiiWd8Tca39uGQWpMIivHTnyndimNeamqASAwp2H5jlnwlqt4mQs0
dYAt9La7J5NIsxQJi6+PC327f3lCBSI/GAJfdruOUXqfjM7f9MzGsDFwhyynQb9E
dot0wd8sBApB+uPTMtjb/tcSF3EN07lk3t7KMjtRfzEdg2FR0S8dRoITQmgdvRcI
PL0lvi8ytNkHPedLz10tbsRdO7czLoq5Kh9CnDBBRfrmX+GKmxaPyHb1d2nQfC27
dZsZjE2D6V+nXfJS3ChlogPril959PKUvvzqwv7NX0i72MTaysT2XLCrqjJ1z8Eg
vO5OA2Kc52v1ueIzJOaLIk+XB8N1lJ+P5XWwnIsoxGsOGWtqbmlfqetXD3jAPQIB
zORDxzADxBXfyeCZzf39293Cmu3Yzq1g/WiYHrOvht6t/cNKL0MT0uKTmKIslP5y
fJO+DcbqVQ9PVgtX1P9kT8Ih/2bXln+Ei5u+we5B2se6G2oD+otbWYYjrNKurVGR
PtwKuypMyluVqm05VADCHHf36v7trOhoX6oj1ZhDj8ng8TTv9RXiqFrPl76RK/Fv
KaWzYiS4Qc/aDCAc7rWlKhuPPMl5I3HK7sbeSG9bY8pCZBpCUbxCaNbbdFAh0Jpr
znsnBcyaFWOsYVbPJY5t4SycSwY/QeJo0Dn7ee1+FpwNgaZdUOGcCQH+pBaesA8I
/ebKSQmNrFTrHzRmtrBqPdSsYLOGN2F9UkqDcFv1/8EoKTh/Ecs2pcmAZz+34Guw
Rj/afRhzY69GBEdLUWWhxGz2QDy5rkt4QgvQxXLpnLEDs+bcVUtpI3PDjwDBr0c2
jmT+TITui7OlC6dMcoyWVl0DPb29eDndRmVv08b8fYDu6VxeLFTZNvo0zgSQ2gQH
SoJp8q2hVXWty6l7//B7Zr479DeIkwSPEdOguLjx9jtudXUXTbCm1qnN2XxawxoL
GgfDl1hDnL/5al8URuPrUKwWeW9/0CPWZkIS8HPcM7SsALtDkTujQfitu4AHvn1L
zNQ0yDTb4oCz5W35xvzJiZUh1eEJhEWH8qAReEUweyodv7FxZK7qKN+1/c6FKfzc
jcTTdBD7E1HRVIBq0BHh3wvm2pgsWLwfEcZDViaqgbG9ILevSpRFFEoP7nLmoZ8c
PfI+8I3ik+v8dI7uGsIMDS4Oh+iqXTEFHMyx2Hcrx3PJFQakYAEFDgBpsPWtEiSZ
tXaWM5hCQtGrzWpEoge81qpFa2VwF9vPWwCEet3ML2XlLjpZek0a9wTyebBgLKoT
PaaucRwFYWodxggbWGODG4yaV+csAxn/7dgtRPiuCvfEIJFckFRnagZ9QIafeVG3
IVrLzZFHw1v3baNMsZDSnolMilmpvrfnbtp5uRudzWXRi2wD6Jakp+qruR4d4GVl
x3WB+dIgn52nb/xDvpK34ZHG/Ct8HdJy0kvIhnaFF2x0YX/8glMzqvIB+YD28aP0
MphsiOpGoL0yWDyw4Xup1at+Yo8WHdB2wlpinSlKNThR3UAwKLmNqGWMYto0p18U
e5rtiOapFqKdK413DPHRLntUIx3VI4Zdnr33xzD9HBG/KBbZsZf4TQAQxvd+lkaN
+ib5H59DrLDo9i/fXyqemF7g4Cyagi+35vQmBL8MEgENJaPptyVLTg4jIyz19R8p
EruJUPRD2Mtcxi7FVW5+2ElnQWdY2I1gNpTu7/vKqyk1+CDawDMS+MzmSHmUJLGV
QMDVs/fzT+Ze+Mw9GK6glk40mIoxCBSsz4iMZveEj/JHxWxmI2JSfNX6WXwSV60b
CUCwnfKuHcbJkbLKMM0LQpEmGQCutlWag0d6iF27gQz5zbGgG9HfUTmGj87S++zF
QT/lm+MueNYKsif5fEXZi9De3QIEFrXrxW6rP0v3Y0JOY6BFq9PBhjbLXGyc2X1l
e47uxsHIpCkz7CrkUhdoKxnrohN4nvkXwRX+5ONZ0n6p1JcEpCSql+bBBEykH9wR
gL9rV+SiDwFnX9yHZFcaRSSf/BYIpTvIkMm2yy54JV4SaHuGK6JP3dv5KN9I1u0s
j/1apdmQHvDCBOHRsyxnQU6qDsRU4LqkMJLGQOGFokJF6yh5Hi6dqBgiWt0WPIoP
WAmfuqj2R5NxeR9FUBXu+vw3m2M0YVk99SvWxakk5yPsLS8HY+0M8TiZOeMIF3e4
qCcVykDIAw74qq+GDfQYUHsEZu/7Ds63ef8U7KUooK20R64/jM/FKtA0H/qBvqbZ
1YWIvokCZtlIKN/8nXjnuPz+32mrqFrZzcl/kHJT1RgxRZ3N9dxNcjen9AD7dHZ3
baTXop3sUk5OmYNMVUl7689ptrXXi9fKkyYUfvtsG0WRegFRyAO+lA+OEw685gSu
sbjh/UQdro0zt7rN9VkdVeo8ggDt7LwvmGGSwyIkG5U5TPJOuuqfrKftgDmetnY6
+ya7nzHs7HsU5zLpxpLZti4WLVWdTnSlA9oVBS3Dc/stbJWkx+pzn0qX7ZTCjniO
ZUhj7CJjYAlFCQGySddg0wOyYsthHLo4sWFjh9JIS6Aps7hFNW9tH5wE/rrsl/9+
2srKDf+hGjFY8IRciVtvv1cwKRqIH9HoZsHJgm4fldLYOlIHtiAChU39yA+pTYwr
rXi+V8e3/ZXw0JkNhlvtARXbWfYU7K9+V25vHXhgUZg3HN/+o75hk4Pglj8BTFOZ
7LUwX2esxqu+xYYpa3jGOnFKWVEH5XilN+v53IqYBU2HY/pfUkv1rJk30hdxs421
f9ynEgr7Ln7xaFt9itBbeN3pOtG8jvGgh0aT9ZJQJe1vIAcTAxnULPb4tvHS+Tou
aNRyz9ZUP3SenxEtZhRXlSvu/GkCcNrDLrlaa8Z7TrSZEUhu9z/XeSQmH/B6ZiYC
kn3aSdQ4+gqi/sGr9/Cqwm9z4p+aTn9jwUcrxsNN1WDyg6csPkuludbrSuR9QdTw
l1ZlbVyKry/QVMWBGjwRNWh/Bz9ttJVNzbZNN53ZC/PZ4SX69BZNWXRp7nsjGJSL
tZbABZYzfTbcOg0ICBWpZjNo7mHwpJaVDaFtB2ZYJyAIGYhqLi+KeOFQR9aJM9ot
ztedkM3e3/MWbsCgtC6N0q33PIVtrh5imGT/mLTflJ88dDpD2FBfnkhxS96ZR/CY
MUxQaTCNeTBpaPNgB5Q3U1K/m7yo9K3iLuuBT/Mpns7tx4YZ6F3sImCE98hu6MJq
E97jhVH63CrXcla2qMJ+vyiMOFeXX3euJpAWq5J8mXVdq7h5S6z6b1S7kOYv7hMU
rMGBS+47pn6S5WhVb48n+akfS8ztrYd4B1Z5yuwHUJ4ff24VE0eD6M9yz/IGHsm+
/miW6f2aRKLz9IdEZ32Ud577IaHPCpSnax5yzG0NfahLNtqxMqLj7mL7KE75mdVr
sHXXRkJ2nkhI05OY4SAhxcHmSGp1FSPponzdUgOoDzXwuhgtJ7FY9xZNTuvxtI0j
5vvd0YEkqivQwYdr7xLmGMr7bQ1GDHtdjSneLrouaTgHgKp47d0YIrjn6anm1zX8
C7onaeD++eeKh3YkhXT0Ow2mzix2vnqB61BsucBnme5AfLxgX8aDQUoLr4jnSHl/
BmuzGyT1RvB9jWCyEWtuhRHnhYqayg6ts08xHwtAofymvbnb8U7W0cUOPUVHY99o
GVkaIE9QW1suGXyOgW3qngjr6amZA235TK6RZrukxBWKODQ2sW69H167xnZe5w9H
LdYBcV43ZA/V3rMwsA5win5cL83vebJDN5y3BsPI9U4p+TvK2h0yhc16IT4tPveH
9XYs6ohmQsYWfFu1qJnhAkopk00nEHcilejLqASnJQdKYjZ3DCOlvvtHs5t8k7Fh
OE/vF7NG2uVvRNfJnCPiIu4dVcVqKxafLgXwUBrSRnYPvYyWdhNMJ1F7hxpQqctB
+JIzqRnBSKC3wCwL73asXtMEsVqjl76aRGG7eoP+jwEfTjA0k+KqKccoc7YgJ6iR
gcurDuXFKxkcHzQHcp/vTT/xMmSEMcFKSfeEf3oFC+taEBr9hXMKXPgBDEw6ZQ5E
yJh+1XlbXq6FvIrStLzmB6EUrPvfpF0JeDGbaRNzQLWBzpGGkpqBML6zsxRrFYMR
RUR07Py/8+h/6kf6HFNY4ofq9XeItvTn25ZBX8NUY0tMzaAzApuCl24oEhOeZuY4
0xCC+tA2WMo7faplhDilxQ7HBTu4o/37nnJd4+e55rlGvJLWy3nzRRHtvU5zS75W
xMzTf2/dEiVAN8X98uHlBdJAR1EKSkQedkwz0mRCqNw9o0L0zNMO6UzedvK3cyx5
y8HrhBr2vUwaIjpXcf19XFUZdEaqIHOfomg2fSWMa6UNxQCWV2Pd4AlhzNLCa0p2
yy4AqqvY0a8bQe/+79ITf/BX43VqN23y7pCt/q3haeOF3fQ/z9wKPIx4epLTnxHO
1GgSkvMu2wtek5R/1PJBhZSwJLu3M+8x78mZ7gFoyvgVcESVqW4N9Vq0JhG8HrdN
V/OXc7Es8nbI96BpVXU3aVsXUyGMKU+HSaMKpe7qqLJzngY10n+54Gx312u+TjDH
gm1TqGyAew3po4gFfVj6XEd4zqoomCj1iKcOQCFfK7TR9UqKNQPdEIgAAuTxmPCO
o9bguMR+K3+ws1iSDkDA55WYRVM54Wt501FeN/DWtDSLjodxDUGXoQuiD4XPH8Ss
TduzRm2t+tm4E7IWlXYx2knmRhqGf5y2Wk/01zbQRHU1k9uU1xl3xw5Mgi+jYka2
MtONXqLM/O2ViUTQatHKdTng8qXHUrLESgdyN6+3AHO7tT/VClHOkcfo1VNS+epE
R7APvgYEbTfCWtI+Njtu24L8Kz85Jd/PLP9Qq4faFFgGLhq0TSfL79MD4PMX6HPL
JlMqCl4Kz1YWILKlEfyfaiJKly0im2jen7ZGiYr8KB0Ehesc/PaQw+E4JgqXM2vR
xtE0gOp9XZ8GKMG61y9iUYZU/eoLx4e/2iBbLwcBYmcsOmy5rUgwp4rpgrnLXdIJ
qlXoZs7eaGnJ6K/8sHzs5qkRS+yORTiO77SjOODRm+xL2Wwj6u2Ru3jxywDApojR
3FlcekbMueuZC5Bqzf/YpGb7f61Z0n+y3XiLq1ShcaCx7sBfJLKgOGa9KZ68Zq6e
tNm9LJ3xaAJb0fkcCObD8c7IzzabVFrY0nQKmDEA0+a5iNXvzlABAKW8YsAAlQfr
5LmA3F23G9mWfAkEMnEZw/GTbGmhLw0gYn5gjApIBjdqjUPiqFnA0N/f0f2Oko0i
FStU+ShMYUYREQU5VZuo7h66wQHgWYmcW9yEHUdV15fF24DNk33ebpcSyT48UCc/
xK9M0ddxhP6Q/gjE+jOrMA9Uw0Iv2wi/CJ/x5FCk9RB8G8kmmf46sa+kYWjRKKHd
pvCvB84DzWVW59FzBkwxCeB3qbdLDm2NV5ZBKymKfQP0jTNnKTzJYyIEmU1wlf2e
zFz/EyByBqoWxttlSd9Bw1iYB5iUKRa/cMib5bbztRxNIUJ95Lga8LIOy9JiCsS9
iKr44oXDNtQ4/TpvZ1MRvpbxKlq4Beplne2SSkeoTQ+fv8ly5guuWGg0fa+PyNzD
TtP40aqAtWDPUu6IANLXTNZEViEDkyykiMgKwuN0C/S4hmimFO2d4XDkab7/5UKs
S8TOwRv0F7rJ2Ecs8M6aMcPooDBsdLMmTAwjek/Ddy1pERlUU7mQnbvqdaGKXnO0
DDGWkxFDib5Y7dt7o6tyxAPwj0Xn08KlPOX/UQIZxRsD1wFE2ldEoJHfsanGRnsv
1woxMMiAXSjXeOC4R1l+y81ffzD2pg9bIdIrcQLwIyOf8D1I02kcN/Yf2ZQ/uQKQ
nkDOkZRQmEGebhB5Yz/kAP9Gr2XOVnoLq0zJCqCdssZZp8FNWTW9Z+qeFKKa2W4p
EWg90jyQNGqUvhy4nJrDONdvV9ISBz9JykN9tZtHzsBBVFmEsFAbmTkV3zmgnSWk
H9n5bX4MAeVw3wPj3wMHLleEuTyh2oTj0g+rKz7uXIRMWdNkbsMXQpORlTY31LBR
rievIwP2vX10+A3VspytAOp9QlUpk4PWE+943h0rwhMF7GI/i2ZDsHVEaxZMxzf2
ZJSkIQXwUBK9BtkBbvcfh9PqTcMMkjYKFbcsxxA88bx5ekPLiYJHKQYbCnbDwH3s
S0W+z2FErqTGJyn2zFbH1IGjSaPT2QY3DMMswg9GMISNzhNTGT6yA9Nx/IDxx3kT
TlPIliSx+/4IivcoG+KTAPwn5z8QfI7XpMWTSFSVgiSQYiDOGj/GA/w3v5T5Suvu
JCupPSUPvIeubtYDDtvR8FMOApZvEjBhluuLApw6dkzOMOjYyGmkiVY3CafK9QBb
6dAKwm5qPcH5YDZkHNAoZWyNbPsU34I7oCS4+M6FEztZvn6H+XpgOMb8NpBJvFGp
iLlYyOfAJmm4JtuHeCMisf34UOUWHzyc2dyQ9QIwnQefL+DvEnb/7NXQS1BJsj2i
H+yX/ZvHtHxcos1TGYAMZCFAZDHGbOVx9QocHf+yBzE8cVMNtqbBi6zVjdH8XPp4
SRaQ8GAnCxZgO/WgVSjx2vsSb9TfK4PjUTyyXBp+4jSBVjb+PV63pFlInMf9wNV7
k9OQVYoH9LNH6K/rgm7GF9zvSFz9Fke/U0thUcDJp0BWTt2tM6xRpv24bHy5Vuf8
OPMGEsWOu2YjKJizbErJAtneG+tLeyzTfW9vc+ObrKNDKD1xJeab1RC1JO9IxtQv
b+n9Mq9MzCee7uuczEUjq+qzebcD4ny/kTZJxS34YyaW1GaLq4NSOvXPurj6snaF
6Iutxgc8A+SoGsiUW1KwN/AWjXXhoJ/xnpqwg1PFWSf2T0cJd44W5mS843sfAT9I
Rdfj72HxobhazQfPixXDftM1FrajTsjMPgUyUm3yMaFMVVjA7sXgDtWwE7v3fEG1
pa6DMtzY7IslwCB8csuj/LnNrnl3Xjrd7nUbVRXvBsm477ycqBLsDOFgoEvcfC2H
2ltTqYrozfJuaI51bfV1HUIgLZdmtdwkWtYzhfjXYrfCgKkaeQCS2JWQX5qgBfbi
bSJyt9VyLDOapIDM98L8r976xP4M9hzFHYRJEgG/SSfLnXvbmc6pmeIYVFPf1+nc
tDIeY85Z6Xn6xSrALYC7jOGQsZwcZTyoB1B20jtXbdwex7GfBSgI0KsRkU3yemPG
rphsutY21oZrNUDEm75Dz4EhpKvR+NcB+bu47p49FCm6cgP4czPGF+W1lmg0NmrY
q0tIjnXyq3AlWwqoYw4vpJ7D3Bhbaurr8JHlfyoPbMrkcHIM9S31mUCClTTQJJxk
bR8puoAp1OH0FHpHCP7KcN2AFiAnBdBzGouuTO2l2WiWGVUgBvONbkCRpJ/YaTgz
oZGmp/qg29APf+F6+TrLrBom7drsxr2AXFAxa2DsI8N+MWkdIix9dplwFhN0+HJ9
7cGH44ER6XAHiGTn0xyKjjjxdLlsEZszb0DOPJzlysoyOhBHXFH/hPwGKMEmiVvK
W2Greiw52Uwb5c/eWKPuRPbhOmr2KcTlxpPWSK7PuUdb6p1UEawzHcAEolV0D3n6
XrrEve85XHoYTPXovQB9xbmTnumTUA8dTWY+ihDCiVIrJVVt4XKQn3J8F8tVUmkd
Id3PtBycjtw52UldSTpz/So9FJDOcvhZj/A7eVn4jDtjd6D262a2r+OIWBrJrRpp
yd2sxpaNLwoCs8M0XQSJS1cqBuHEb10KCVfBJuynjBEWJxZe2E6ugTPuRQZOEdE/
9afiOGBEeFxY0cBCW7ZEL6LVkIlwdJBn6hPnKUUrBoYNv+cl8rgEwXXdLo2+fqnJ
IYnUzY4VJMHs8/XV1rFh9JXSgcZfkyHB1ScUYGSRNe3rdjg+HuB0rtPUGoq33UE6
elYghG2yEE/AEPKYYTJf9/JqQ+8J1FvE+fafdT7g3N7Rf6YQIzRkQrKZ24/j+qWY
nh/l7I4aU57Zzme5BdLSslbaLARJu5OKMBPnuUWRzVpic8o6hNkXaXGLddG6eELw
QYU35t/RnnQaNHB77C1kXBXWKUy7+aNCA4OZGo/LI8R4IBl1fhe3oADkaHapk5uU
M4ijS8bD6go/oY9gnelqdxYvaBI5Gqayftv9MZjfx0kZcP6qnyuGkPPLpUPFmMhb
pWKSQKDfHeCgswrVNdP91LDPHpg4ToA2eJAhTpzZg4puzGf6IuxwDwmzZk6EbKyS
BZHjse4AQGoTKVrgh6utp5CRgQ6DY4uGsaGuhbg79BOSTngVJaWyyWUGbpYH/pzK
R1MVhy3QIP78S1GrMOi0CAcQhjoaI6oLiJBSSZUt/QSL9BgoS/nJHdKlKf1/vYgQ
iVMKMKnZi/VaSVRIZ/R22gDV/kkhqgQbD+T1gaUL1sTXRy3dJ6cMuOpaiLjIkriS
I+T9UQoTbJQLr2dnw1sg17WuBZeqBMd3C0NvvNsNCP6byk3/yhk6BdrD232IaOXY
3r0ZP0Qn/KhIbLLtXvfEMG+7i1D4iIJCKuLhFEX+h/ZW2LiYBvAQID5LZAAyYeTp
740yNtU3bsEsg+Fj/+ep3Juult0V1ptkIzeu7QKehubBxURqupCWjD0nV5BTx+pY
t3HmBMqb+NiotbpYiQ0tTAbJQEaUiu1UttXNlkotB4fB27yvOCANSX4qfSyeXXy1
BiHeo8XEfse607MW6yjBxX8uv8oNKmKSvCW2igAnIumH+ZfaH2rfkNcSc7erEuGl
+PPJQlFvBa4ZaVsDoet+c41Gu8nz2ZGljuxoy7zTUhk/1N+wRafODn6kVeC33f08
N/XxyXpvIEic2mh8HOIyclGKGixDoS+NdsK9+YVQANfe2cL0KBOoTZVWD2Ma/w+4
mNB9Mf11LE3qhxzaL1UIRepDRF+kslHsGI9uhb0xBN3yp3AqbmdrW7C1NN6fLdVg
cVhbZuwI1q2dS9KZUASPi3yyrHpUTQuhwydSg9bU+IPcu1DFWKVEayTOR/yOsIaS
Xfa0WPkm7gyRvJaKe1SPmsR9Nl12ogrv8cAjCbxuDEOlNNYaMM8bYxPTGBELxlt+
tddXodNwMMhBzPcMC2+CO/MiLd51lCQEDdRXY+D72Vffga4yd1FekD2ohg2Eg2rC
hQZ7XXjxhkJL69JzM4lD+hToem7nkbo18lGGHpvsEKcWtT9aU2eLqicq8niSIdhq
I8WRnwWlejznrNKkQDOtSqad/QKKB6+mhab1NGiowGKc+AWa7XvPDwqPfhuRQMZ0
yKWjBJksdYF1Ps+B0HK1Z8etqIBuu0h6e73/xVPfwLf8Vij/YTRF9aQDcXWA4AoE
Lh/hAbz+n6NPZ6vUVlbQXlgJzPuV1nTxwYSaHP0GY8FjDVX/+tzWBToENr1Rg9kH
FAEpNBPwW/w2UzUSdb0g+4v9g0BNwRmp3bYVr47MhAGFDbrTbQPQXUXlebarNK++
0d2d4yp3qsYFZbilZ4O/ppamU7DGYgoQsACDPH2hGZpaQm81l0eR2N5z7NEpf0Zx
DZ0/X6EQKvJVFrN47QCk2OQN8nslDCouKtOWiGYknU/bdhoE4lx9jCrZm6UFvlui
+8T8MT5+ORlyxtPSW4ziO2XQRX7uE3bvLoSu9rUm6f+4VETDYuglxZ6Yd6uRnrfI
D/41SCqYdDoGycoIf5Q4XeFtYqEzn7QIWIfBDg2V0dqwdnsCfARryftKaNIT88Ds
MtXtrD0E5pP+Hnl9lPrckQG+Tb2CzLt0Wj8oc3peVgfT3YGDKRHUBv7wFURRZS5i
HS+3pFXa5up2QJMG8h6i8UAVXh01oZZpDPX2fxPGhmws/khBY8dZhfAKjfINDNNk
CHuSlwbLiHJYjlrXlnPA4EZhkfVQzVhJJ15ACB6V7ub55oMJ0ey6lOUj/dN89t93
WyERIIfGf0bNlC1XtZ1+2QIQlPOrQCgb9ltgc4us28ll/hEKsKQbXki1aMxMvcfk
qMCCaJFw6saL3olZEKAiIjEExR5K5bfkX6n/qaHIXDju82/P6K0ehY4Co9RUG5r1
qHL41t/grJxEKPRTiRjH57aFcvwzzpoOgRVDaVrKsM8XG20ShdO/Y/tVnr89LWnS
BGtuIX42M3gyNDHhnKL/3Nye2ExRgztPjInUHpPrlXbqMtX/9YNsW4/reqU5w+Q9
u3KxZ4FysBpj3UFF26hrb1YOjORNG6ns8/0mhA5MVs4gDpmQgyqbGzm3XiVev2bV
MM+GPVAvX7XI2ZNo/e7fMM6iNkVolF+2cNYAz+U4mzFwzq7NHIvKDnJ6Ga1vmn25
jHmnortj56FJIO9IUbezXa2uTb6K4Mo/wWimHbSUzRXlt8Jv6KRGut4/Cev6NR3k
u/i5HI9AlcYKccz28g9A3km4gyVD9Oage4SfPMCmA0VgRLXF8gqbdUNoxUbytUu4
OG+s6v8F2N6F/7xAPkmnbdPqVc/OZSlUIG37WFyXciI6vO4/oLyYFVD96Zlnkh9u
YbeS+yTlw1MUArn54obCsRD2ioOGIiG1oZnu6qRt3XWhQj03IaLHkipUckPAq2gp
NT1vYIzP858EF+twTM0Sd6ucalZF+jjrAgwPPH5hVAoFWEDSCQtq401FAFcExS8n
BDY7V5xIHck9hw2RQDi4no0u3jCCZYnl1mfCvmi4DBs6Vl/kqFB1P8bFCyIfNsD/
WsHckVGNyGmijia2GfvPQzde2XEvNHzna9RUKs3pX0iJ1yaCCIx/wDFPNzpCSlYW
zLgwIG55I0MThqoiPBqizVYFbDDKh0DgVLbaTAVGYD1IgENZeHHovwv7GPXDF85B
4DvnA2Bvu1XqfWg1J0PnpMKqzH6mfbj0isJnP2lURLwxNVoZU9YiISBhRyDmqFQJ
PtOk7YawJFhaEsrkdI6j27Kfgn093/gnD6LUWER0miJhjC099ypU6QnmISOjgRHe
X2YgG1aVJ4kWnrMS54yarUo7Dh3gF9XXjvYapiNlgZCHCxikqi4HrPeHrGE1uT50
94pqgOvkN9xGxIcDPAneDtM/orOeD21o18mtZPnVzk0hrJZPZ2zn9pGPUPB9kcRz
FA0mBBg1/nbKDOGAkumNUqu77V5FXCSX8i8axt9ZeyT4bRq5Di9MJbxnljK7yHM6
G0atmmzyG5HNneZMdKVlLYQN7qRIBDS9BTKWMMJOWYEg0EkyIQclz6vb/PjPwq+M
l2c41MMTtRUhKTQM2Ie2GJa9GFFb+lDR4d1mogk82AoFS9D/+Lz8eJ//92eXmw2d
m0tWZpfTSmquMfvPkc7KtNFR+awt29WEFXZBmjBKEygs/8Eu4dAD9NeWb+Coyi9S
FVKUr42PP0GZj6BYnSeuwrchEVl1XnryobYb2oUCYJ0tCvJxoAk8Ixp8scw2JBb9
Vb1jM3cB0MTuQhCZJd+W5q5dF2ewtNbxC23Z7mD2yAlR+nl1TXoFkNXreMKmId6H
gUVOtgMwcqMXLlCWoFCxzQjG+VBfFo3AqeJpUP2x6sGRngqsi/9DjDragiva/xHN
eoQx7WNzAT9r2w3dxlu74+der/0/u9Jr7l8X6XmBykEmEKuEEZrUyv2zJU/A0xBj
cVj0azAiX42EDbGD2zaNEB/XHIfT2TEjkd4yZiE6Qj/ggckmvxplLNx8Y9V6zrZo
3V56y2Tf9QQjUPmMgspEElIPV7hF1l/yYsMkTtrskRRwXGOuNL2qh6l0UCg7yy0y
Danr2gpYpdiApwXWXel7A25F503e9IRO+4vH6PxyzM0AAES26NCzSq+ybp2UPc4T
mcMLkHfWchwkqoNPdsQWsh+t3NJ7/0SUwOiq6n2w3dWp8cmMwpZp9gWePmLp0Mes
SyiRVMVjSSVpx+YEO12GIh18on1EM3tPMLh7BZE9HRy30eY96ZOUR+LY4ETXAR/R
rm34/JEOFashahl0QbJOpFIO9uf3CKBPKs2pOdGtLZl87QUl0K9GJ567DHMQrNHQ
yjKIBLwjOM/xxMII1YgwTGJWqKwDtb9p+Y/IB7ggzSuzgzGs7Ft1zp7KMy+l6mYU
L0PvAxSBKkgnPt8bvqmabQvQ44q3ssVKk7tnsA0r3XgTryYRQHgZ2/vKLas3oQp3
3WiasmYBpjQYc2gNnOBlXUF6EFrIMUr6SfZJN0UNQHEhIZt+AwuW7wQDalZL0fs4
05VMcJ33KdrnUkzc2LHap0IhvZOb+Rwf6R7ymABTcATl8sXap01iniNMT+Ixym0x
wC4nrMA4nCSbBrd/rnCdLK47w/R8q6I+93LIvZg1XKQxZn+0JMJa8KcNfSMRe0Q3
WDEy2QEmICeukXKrfdHYiBogmIpVCx6BpUFO9pqgHvSACmLO8CEDTr5yNklLgBlh
mZ+/BuDbqeo4/x8HreO9rbmW4mS45sVYEd16u/W8+wnuz5GeFEByLLGDLrvMmFGr
muPR5RClXespmWW+lUY0KleyACI6jU38XKHmnb0YN2CDFQyrxHa5dCMrcHNzMKka
DZJdq8cx5Xv/wcWIjxRRtzBNtBPn9waZdmeM1h5hzRNHAybn8JWmFbUcYRQzEIp4
cDwgyO9KqCOkgLYirn8zSF3c+0SbqKbEQHM2blBAwLGXvuLa7IxTICmt1Wbf5Nf7
jsXm/1f0Y8K1di2jZ3Gp8RitCsQiEKVtEAESWK1PIZkvP/nWgA7I82aOALAieMav
Mg7DxKO4pB/Q9aY8K4ahinfkmZeHKEJtfRcFeJCUdyEvv706rwybareM0eU7zBh5
METwrMoRKwUaDm5Qw2WDrVlm//YAurYMe+BL968mOhDCIO+o1gJlyb8Y9+k5d66W
3Bm847wmGYeK214a1DXB+BzAe47mISSyVCqMg5tik6JQGUjg/zWSOSMCMsuEv2sG
1aDVLyIKDMq1VwtzT5088KW0sUgZHek3x8PlCNgX4CnvMeTsZxXZz4WVDHjnaFyJ
3JpnqFZQgHgR7Ao0ftk/zwj4bX7RFtg4M8ba8lZSuAAzWJOWW1QFU0agbRJUQh4Z
zcSXGHU5LEMVFGfUiwRCy9yt0QVyfEtL8nrrnO7YkumeyptFzdCbIsvfE6VV5Yt2
zSkwS2zDc5X0N7HGcUfS15+lODCFuODpmGYLXCYzxEBKKIeoaEvWSh/FalsbmalG
65wiPqs+9UPrR0hy5wOFqd5773o2aPG7R3jF7jKRqf8R4qCejqHWV9ViYI1fuYD+
dTK6PIgR7csREYBwIEQjD4MRZFsq0XQE/wwxnaMhd1QUy8F87YIgboxhGcb00iNk
WglOcTg1nAkN4YXVJVFJY/Ofhov7db2LgXwDnPY9eS6XJp3vziQJ1xWMI8sMJgTp
+RekSkAr5WRgtZdZbcAGxDDQKq4YUYQ1o46h4q6sT0pnbAL+Bbhhkr7jqLLWRlQL
3L3IxMt1zRvg/ASc3vtLe9KEtV7RGFp0qfkYjqBNKC54amOOcZItbPCKwY2XrLC9
HqUgxg1ytQcMxBg1eQ8MM6Y04RsVMHDXS2F1O7jEOTtb/ISUXFcS0cwkh3UznWDd
vljkwYgegmfsSKTZa/z1l7jkZ2laQSpmJ3dlxhm1FiIQjDKnjQaZe/Ys+AeawCEP
/w4U3/HMhmSvZ5V4gwk0/OZhRfUkcs0/JL5gDaHQINWU/I2UFiKFzluF2wsfH1O3
Yqom3GckXZkd/lvBA/WvIVbO6jck8H9RPyqPnmj9r+loP9sc/B2iqt94pUhR3py+
u5P6OzGHNkKQ03nWOc126MoUVLqjVlFGak3NsXrl5FI1ka0FVxjRkJSyWXOn6HtZ
Gl45hYZfEdke/As+FOsmHOjrmmb3qsePC9R4B0+XbHbTtGrwdI0W6oG/BDMkuebW
KOoTxovdA/X5od9/v0TfJuCfqygUJecgYtbAR16TKoaZ1t8nAaQAgOkl4OMJOJdB
cO9d+OcANoLCu8OKqZPfMG5WR4kcTj9C0GDRIm0qgVLXBkWaPUwO842Do1GqZ2u7
UTuhPd30MBGmrkdVhzEM5+PPH4BXJ6sM43v2odCWgrqn0UDvN8kYk5bZIUpXtnJK
lA7ol4WW9nUSbw4ii/5WZji+aLHuVcBqz0jaKIfV9dN65rOQg796ConXB1VwMe7u
SZfl1HZd+7fJspvxEVCebZS/ToGa/VSKrdS7Vq/h1LeK0/nc5pwKsT5ZsLdq/Y5s
Kl64SkR0Nr09nFCQgSAKg5i+Ksw6rngM3fZE8iR1kWAuKjabsp9Yy5Md36nwoK1u
PJKo6rZL0pm70eDrg9iA3b7IQaUBvtvzk7QQqaXmWbwv0UPlLITDVAf2WB9UWLXO
NS+C7+KRxpIXeF+TpjfamGcPUQ1vHV9BX3WxSNM69Nxw0g9o/g6fKz6xLwkG3m7q
QNDsPdTX2HlGuWCEmmgE9LVqFe2pXUFJeSd0Cm3T2x8N2BOJUrvroEYnBac2GyEo
FM6iwzR0+1HhT//kbf2hKfs13eBgYjhvPo99DIylrPurUuXsYjQunbY7ZJiyY7Ke
UUKgFDX+6WqbuOAUwbYGEJH+Tkoz+9kX5xqGb9/agMVYdqv21gnfb+UINsnzZbcn
eQ580ojqgOQC7Ecrw9HQq8Db1wR2mLeZJ/R4Qs6VDUkn3EYW3K5GNi4b31ShB8vj
654q6B071E9/C0fLXE2nb+TvEjw+5JGRtTbZ3stXDA6pBha+f25oRNjO8vmjYigV
KWaI37nZuo8A+09h9I6jr5lPsiJmkf6McJVdzp6UiKMxicWRwRjHF4Kq9aT0p0t/
2AEI0pLOnF2c2FWM4q8Ang6GRGsALiSRFg07MvxK4tteR+2HVvzewLv1Qn2ltW1F
zNc0L8cKKsKVkxxWCsUghHFvPakP8/8aIBzswvIM0n7epRuUqjEJqSttpNmIHuGf
7rf9LxjXwlxBUHB74VydrWcYME3R80AtYWYYBdMAp562/xTqcGBOztXxucy/uzCi
pdN8r3jgql2utEhdYY7Wj0zpwtnBQWsHE4s/a39CU3YOFEfrMg8EAsO2ebXp+ZyY
8JCqqp8YFP9J1T8V1m+JbKJflPt6j38xOyVoHLkcaefWvMubcPg8IWeyv8a5vtuR
lL78jeWEr+WlgQ+eynXlW5Tfl4p5ILZGaJW0m3VP+WusYzj9FxHWrklZIAdt+qx+
KoANQwPn8CeKXdMLmghuUw/lkJg6M0BiqLYJ4Mub3DoD/3lZjoj0foff/PHeDqP+
GfiC8CUF8YUt85q9Uj/Phn2JHGyUTXls1xr92r8zId3dKSHZUe5tLRK86/ERpHqD
6kwWRYEAW/pz4Fairr5aMxa4n5WsJZ8mcpu3DH0VdLJ1te/kqK32368IPZN9JTJO
+n1PQRZPV63GlhaH4Ep9Mm8qfPXvkSC3zRourF3HbJ3bo0z4u2py/sycsiSEsbb9
vWP4/Sho4YEGzw6qhJ1nmgQbOApoa5EOf9POZIMOZiRP7FfY6elLR3wTk4c0lK2i
XWz16e+vrEkqEvmlV0KEYdAQSwXYWNi3/dp9L3FyV4Vo5on2McNZKJrHdFmBxpWG
SkQ+YX/HfK9PKW7jrihgRBFsSw4lT6KB65jKz+RJx/ZykJ+PhAooxjlMPrmqd2iK
lr5eGGSY0VcScIQYelQp9aILa0ajcfNC638o1Lh3iGrNj2HGGyvi0uljRNQcnUyq
zzennA47l5//YQIJX6x1NikGt3Kx/lA0le/ACKBnT1HIzUrbLgDyDPPs5pjq9Syn
Xhii3TXkvzyI0SlpZpwDGojxhCJ0vLiTPin7SI0HVnd19huxB8RqqDEiXoAp27mi
leuL9/YDZSU/bltAshhMW39WXtNEHDewQ6kI3F67bPO75lAaK8Tip+VRdFCwD/iG
Ynri/jC0tuSh9IN+wijO+M/oqRywPF4zLSSpC9DxtfJeQxGwjEnOJYb8sKnrVfkX
GCfj5AsshsX1Pna9CmKKg2Ks9vqdrBLxPePTAnwaxtTQJF3WvdHDuK5UaMaQeWCX
qv75Szz7ppwNMt+m/hDZL9j3Dwuy9rZ+7Ho75QhxAd3RWoOxOX2euXQI+hS710T2
qvp2e/4O23lIcJ1BpBINKxyB62UHEEpFqg0pVkX/MsE84fHVALTvm+IAClhLvGF6
bXlP5FTYo/rB+Fys6EZCHT6gvlfdcLMRzGtPr2eoiRJXGk/smcKDwQfZgVT1IQDo
KCTmXYPtN2wnP3JqdbLXNZICLaHWaEiOsPr7Bkf+TxuD5815o8wOgQ2FkcYMpIrb
9+AFKc0aUWCg1E0996UvpViqwgGLlBWE711RLFz0mOCe6UKlKSGSAynSy7Zm5YJJ
RWrwDXS3SDPRKFAkTWQ9NwSqDUcoWzadf16mwC3AkPz/gar0Mi1653DG+V9XoZ3k
ruElgrY3xU0+9qysykN7vDBdbNhHCNlml/Pbd07nyM/ZUjoAzf7uYyt6vpYSeP/2
m+7va43GwHTMAJZYERi6K/pu3gud8l4GVzIlwR5mvt5LqTKm6b5Lb8g+JJ7K4IV/
8ihkpeAg1OMsYdGOfhtQ5X/apN7/yGyK4rkXJHcZJzCRhCsgvjOTZw+at23AvNy/
5jOS99PwwbH682V/D+MLoGT6V9MRa1nrzNxmXJPdu1s8stzzI/7D//z9cFNKmdFI
JuT30O3pfSNwGmPEAa00Q4fZA22AXZiV8qTSGYQGrdSf70nU0bixOJpmG8lamkrt
GnL3+8d0xYT0ApuTuIMZDJNJVxitWI3GoHe3fvwRUNINIAs6cSkF8XK7K9RQ8I1B
kuJPyq6UW/PCexHRbn8hq6aguQRJkoQoOg9Z/yhpdkNjHFj3W9ltq2d3yD5Iut80
fvTVh/OgawSRXwX+v0dalE8g+P1NseN8lNNtmP6y0yJbelacA3LQNVno71lggHTA
CaVaR+qJ4uysYrrZsqFwISj1uxosoG3vJhS8rUfowR48KlFZM7wLpHyqozTAM0iC
u1RM0zrBgyGujqFKMOKQFQngw2IBS57PTBfUFIgdg+u9vtp5sS7I2oJ2OLVbrhWP
Zm/5No4ncTgrpWihv0rmB6vP46x2FnN7U+/HSBacMSW1v7dvkA2WyaxOb755QbYd
fQtkyuGCuqT+IDusUMTuRWDV9G0RqD7qCRykK0iFPfzZXS4x984qc4UOj4lJxopJ
`pragma protect end_protected
