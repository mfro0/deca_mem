// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FQuldX1BSgpK08RiMHdYDkbwI5wAc8sb0ADkBNn4SKvN1ToP0w9NFx0nwR/cbJtr
iHJEzT4kATRiAtdest4aOxzp4Bf5ZhReI5AE0P8pM6LJ8XejsS+saxpVmpg04i2m
iUD9oXSWULVXeYtc3RX1Uheo94JcDEyoqkCQuMoDYF/0VKq5z2MhnA==
//pragma protect end_key_block
//pragma protect digest_block
1Ovlg21PBfbqGumq04Yfvzdsa+8=
//pragma protect end_digest_block
//pragma protect data_block
/e5ftqiqlKwB2h5HcVSF56RLTIr9EQbNzMx1z1XWggCgh3WsdaG77fZj2aXhQNa3
6q56ZNcZ4pJ/0CrauoM7MloStNQ5DmnivL75pkhm2Dj25WZaWykPbmsh26zUJvSD
v6ADH3KU/l3CZtpWDirwSRXsVXWt0z2SoUivbeC11x2bbB4UCVXDEe33MZEkvkEh
sqKuUflYjmc1CpW9QIIU6yUd9WYjsvGE7TF2krBmEi8VAch3hfghlNAVdDkos1SG
QkhFX0aRBVag7wrYNByGws/f6ECqq+uu6MVpVIvEDpL0VKFCpuZSUJYO4kTyDd+Q
VMh/ZrrHRZrTqyzcReDf0BbgK+93R4Z8KxKvsa0qzppXxokQyzFBuXuubYp7c0TC
i/v8wxHccl6qHtzM9JuVGy06Ac+ZowOC4WycLZu3SDW5DboVWyFbj8uF8INomcpw
gYpqYVfnJiY+DQLAoxlVDwsQvrWG1eIcOUetEdnqdnn55FmhlxmWYR+qTXaBiiW/
vjRMkLZ7YNNgc5LKKhU7mRrZFyQxuQlL2dFnT7tj2JtEm2PSFJwInBNjyAElYRn6
usmEg8CAI85oinfziRqyPw6r32n12tJcWZEhSGBzJn0MvRSqrSEFA+0Twa+zYqTU
mz9wk0gdJ+AavgdwQtlYqAdb5AfsKo8BN8TBaWVyMz2FgdLmwfslLC6QMGXnXggD
LgPVmWsmyvhAw23ewY/RURhDonmcHSoqGuLsZZAo8yg6Gc14F6KHSkwXKhFKG5Pv
t58zTyUQstsU7NeVKMLELt10LAv+Tx4SXccBvAK33OQ62GouCzQr9tABT5tpxllH
4ty4xPmhzJH0VpF6sNWrXNIr8jyzFnowrGXGhquUTF+Q5pXIT3DNPMiOYaDeJbTs
6le5I3KdKWTQ63xDSwzGCUjjN+MZG90W8sRjlhHz/mgIqYrWcn0mUDPhs571SeiU
MU78n9818RdQOcjNSLWa9RokV7XmEUsPSELtZA8cCHbEwPwGGmYK0mS+A0cDxZLT
ociUtkmgi1OjLReN2pf24GbIFWWFfbG7xLFHrDOWui5QeavThaYLpiOWrQ6V8bEa
Dp9/EJj5U3gbRIjow0VHLfiN31FtbYsmU3C/i8cO1PelH+8kjJhLyFkpDzJDI+88
2k5KInX663i5q/U5o4YGq0JSkzqhJV9UPHumjt1MonlZ7NtdT8yuuP0BCmc+Dzu5
AcmdEEplfzamPEvyLRwN313ZWxFqx9IMLwnaVOSlVmVTOLq2f5E6mrif28hGMBup
311kR6tD/SSa5nwJzb2Kjh6JNkYxIMq0FiIzHLMFJVMfBlYdudLLsBiiKELnlAAc
cUuzbdKHTlZMaWFZ43FqMlxkdTeTYEHrihvFAhG5r8Uqam7fLljfPNFlSr8P5zM8
mLo2StF2a+h9pvgUths98k3ZjFIZ/6cfSY6JwK0KCxhuftygXuSX1d95/Kjzy/5t
lJ6liMV/8vI5unj/it7uyaJJ46WXttF0dTfuJ7zF1xGfEJRVthBh67Sm4AIbFtbb
NURacs67kTmaUa6fwba59IXZF/zzA7tAIErugi8KGHnZ6q5m3etw10JKkoCNxAyO
X3YvUN0EnEXtWiOmcxGymxrrFmpR4oVUKew9L54ES1lRSXZiBVmTIJAhYctyf2ou
18v6kwANVKwuD88JNHkdx+7zsHme6UV48KQDHb3NtxRx5LW5F9U8VYj7O0yRVX+2
ea4d3W7bl84WxxWhp1Zqs7+V9iSwh3vfEFVkgfFlHZkoiGk+gthQWf2nSTdONeNe
iq138d8ivTBKEeSx/Q1nxCdynu/OzYE3OPnzcDmaZI0gRevvpwX6sE4vDPIkc7si
EL9p8+o9jQj9z11Lg2EvXKVImxtuWrHLGvkUptLcVVrW81fpJEZjny7yMMtbqb6L
l+nkbNQ7atlZk6ZxgESuP1b/jPg6ztddku9ADeh7oA+HWY+VAyvxeEr15l43AQNb
DcQu9JP2Ax1Yun+l76QthOzAApoNTDToLc5GXJvAf/Y7XaUuaO7+n7tg8b04pcEx
Nte+GoIbnuGBb/K26O91WnMgoKZ+kHoRXbRoghwTtdkPF9l8+okzi4J68WkC1oh3
x9gl/qc0/nCL08FZrU/qcFIthhKPoiOh5GX6iqKztaBBlymUx+vI8U7SU04wuTO3
yPvi3hfdihwt5ccVDTgWCeQNlWwx+p4FgZPGYKIjZphPcYTyFGYXK515od1PPCxI
ywPy+whMRP7xmD1/d0CDJWKgxKp8NQA9vJMIpgyA6mdayIqrzyZ5i+9m0WKgz/Cm
SnQqN5YRKTofF8TS6cFBE7nBteNISKmumt+/ny+Ff4kxKFSDIcWp7Ih7WpNlcF/C
6KlSZk4d6Qr1Yv+ialNISTbdnEvHU3bLrVKd658AAImN85u5hDAJb2UhuhLq5POE
p8r7kCpf324RhiVei6pc7I2wDnZgaUaPYzEoVn5oT0PEfXkU5dbaWuBZKFQxl1de
WRR+AsKDQErN3Rt7p/Pk0gp5C2nVJ84Jjh04IvIysIDV/leGNdMtXRqmcbVu0cD+
IXIZpjVu7beVuVYImSbo3jNXhFCwleOl8DGRzooGZjhz+vlyW+aOpJEo0sv3wiPy
j4mE/w1ui+6/6RtXhUEjv9GaahyFjvVICDbj6Py0AYLvgyTfBWFH/coWF10fvCVS
4NEyEpkjbcit5J5gg2ia33X4bxaTjTn/2gA8CGniN3tCpBDfMK+QtmOd5QkNHQsq
drKJNEZrbCnNezTMGlp8Rarf4yTu6DnN9UCwksaw0LCO/olvhb6FlSgZyVEG6LLJ
WpTkDMF14RjXHgYjqv8cOCX0HumIY1aWsQuC+hhI11kCy0gLGk/1uhaFLrrVvA+4
MQ2cbyU2OUFsr3ecJ/8AIyJ2Sw8V2vNxoHCksMFcoshM+h81rF+N+3hCeKTcUDEu
M3s7m1keaCQTiX9Q9O093DNaXUlLX9HaKAri0UR2QBdhfkYtAxlIGidzEWpNS8Bo
9LIQQQ+zzsiLzC4CxCWX1u4ZJhbxPceFI3Y57Y13YyjTHlf776JFM9DkU8IWqG/W
A2kkD66MWEyLKRJPYvaYJYbSe0jS8SO0zIN1blKps5+o1quPYe9r+GN6oSURPoMW
uI+NrF2nw88ebxItTwUGYOEd5u30LJnRyVjR1d7BdI/Yg06URzuCC8oBwm5Dr/81
J8HIsnosXsm7pwT+ExRDJ66UsKr/nwAuBmOupNuTVPfed/0ZujiXt8Ljk3pdxnKH
Y1fswTlDkPpbGrebgTVlw9HyiymS52OL9LSBIlXGt2Iyg6C5WB19QBdkflgUSwDt
DbGI1J+EGr5qcBc4T0ueRaJMqmK19K/0iVIgx3iPBGuQmnRcZ6pkCXeIK30UvCJP
xcifRkZz6GtbCK0eUN3ed/hZusQrbINihP+Bi7WwEzqCby2GevKJIPeiuiVX9Lid
jbmDIeGXYMMhz/iW2AZTh6bxsWdVGviwmv5PJ6seA1KB1kCsEYjRSSA7EJe3tDnb
pyUrknZ5fc2FClPzgqrQyF2mXXOfDqZS9q3gVBHgMHuBBr27vM9xHVTcljlJGiOP
JsSpiu944WYBCRQiBV+h+OiPKDYyx/WrGN81Hlj2vtxsBhbcL2RcXZ+6WU9AFm/2
S7TwO25D+i9S6lIfhWUEWjVLIpMA8deaInk6kQLbhEQYy81e2mLNRq7MSjyo6Pfq
xGv2gh93O17ur7z1knlxfgJUE7a7a+CdG6Ja5Digj90QOKA/bmAk7Pc1Jz5zZ6hd
OTY+dHR+MBKQVcvWoXuwBk0R3SexujRIz7on7XGstuvh7LpjZdOkz6d9uY7JWPM/
eiTGAgyb8DrAInTPKlg8WVNIztAS4lnaq0azvUaB66lualvVieE4TU+xbMviPF6l
drlaYx/Vo/36QP6U38Uf7Wn1L5boZne+ow1p2T4xdcyzPBVJv1kLNCDHV4vbZiUX
kMcHpnkRmTmknKgcjvTDzKLpv+w931ZloemL09a6ONVwA7FHk3noPFrJX4bPKOyV
ABgp1Qjnr8AwgCvLBXV+3IW4Pl80a62iS0dEMlbLBipsH00I0/4SpMRHhhgRPZIr
V0HirG5sBBFbp87cmMlZex5Ia0FPzKL0yEkMij5WPDc2qqJMfl6Z87Y7a5t3GxDO
Jfxdt9hr3LS8xdP/kd6CtZwWKoxdH2KzesPHf5D4u5z0eKRqbAs5oIWdx0t7aXpK
VI/bPN96n1mh1R6/HZow9qglevJAAYsTFWiaZJ4tzNAoK21EeS0py/CdyHuCi8X8
ER6wfQnr5t+/eBlrF8BXBtfqgZYcvgqOVq23YsjcrfDp8B9kb+x1euPaCOZLm3zU
GzLW6eUrpr2KzSJY7MI3++bospfARpDUiuJlQ51dlLPv8AUuda2jJBaWiu0OIr7s
oHT3vMKpDeR1VEY3RcKNM68X7Yb9RWC0jtHSgZeHchW2d8Px6lSQF1XluSrbweNg
3g5jeTVO8v6UbUVWkmElDJuiDiIEs9/7RBuHl8OXqk+vFbVKnHKhRdNpg1/N/aVT
AC9Ql/33KBaHWWCPviXTMLgFQZTkTYsEwT5LTVsblbSFqQOXyxvwdxteQYxCQVWM
sf7ZQuK6ert3SMVgbqAYRU9avRBTHAIP+oeNjmTK8Bp2OIPnQBtPtHJ5qrIP2XBg
Rjgo+KcYNj8qTwm4qPycmHAOq787H0JOge8MmMQsZ7jgHAlMP7r24wpa+OsD1PKB
vWNX6JWwrVSz6/wZlTfSqdCmLC34R28dRJVJO6zVcK4Q880eNkqH7H5Q7yYDlkSp
UdfEECAV/F/Dsirid/qhvXCoqc2jBhAkcjJKYQ2lFEzmCA7QljSg08zTakUy+bGf
Y6gkgJ0YKjdVUic8RnVTyXBCbEn7UT/qhFp71XIumbUn53uFakRCQcUozNkSMyNh
S8UdggnfsSTHqpIlzWl7yURM0NtYKHj0+H/fb4N07yZeC6QsJ3c8mCJXiz60CA5C
i7oYJEmC8KiqZQiZzewqeCcj8XDVdjnSCoUnPv6vyhCTBSaQvjIbEcBNPZTuUe7b
D1bxBww2YvYdBrv/obGqCu8EuS259Z7MJSD0Dj1pvVO5COcqdAATN07vPPRge78U
yiTrcLeOm+oWuigdI0nyN7gipegAo7Z4C5DFQKScw6M/xFlae0+OxEOAm0K27hPT
1b/GluWPFHzrv0lWFOJythFrViS+w9SYFjcWcJRSnNSwtWBWRb85JcyuYKb6ITEP
fF0nfRpANtcYs3VqYacSrHQcnF2W+wUu1uoxuInk/p2V9ATe+BkIaoiqFWPth9tk
N46eX2Nl7BAC81ZUHKd2OWrz/UZqzzHzPaoaieJXtX/6PpWePdLRrIlNGKCjxQYM
pS5YH/nwpwCFVDcAhuG2A2itBkGFMLF6/TE46Z6saizo9CKDoDlL8OFnyxVxAieZ
2pqtCpzKOBic4uoBsGjvapTuseMuKsZaGJ5fECsGOutUmlOfab5VObY5/T4h28HK
L301nSddKN2oOw1UyJF15iLDnik4ZuouNQy/WwKsmlWnnFH/wDornVAHmybg6DJP
EtBYlYF50R6kAbUsEF0MuA3XK965MvHaUNwHNDJu3Ck9Ir0FycjwWEToWBiX+Pya
KodhZGPLYPqbo/l74/uHy8BoDN1bJ7DvSxJxU6g+rEqUgh3+qGBHg7kGsPBRPYnq
yN/8PXGEXhY1nqxIbYUhuG8DPS9FcuoNmvAASaTvwkqIJtFKOdM1jz87M1d7/XjO
pv1+hjNzcqgyKVc56Kf4bCFfl67485EFaNGRPYESOT/mWODP+/IwPk8kDhdJhkqH
tyoX/h3XvHgYv6pOF8t3CxIwCptM7bgBbngZC/ffQ6BJkt7GguZW9GPEMgUjTApB
JEHkkSVyllXsfpXMu4Jim9qWKNm+QzZHcOsPTw7EwK1TbQym1B6re5Z4f9HdpL07
CYHF9BcVyRDk0aNSRReRkhlSKwFchqMNv1m6vPZoHLGfCt9vK7FxSDlspwatnH4y
YCEqaEzaDTIQ3i8/RHpCPUxvDTuHVklIcZYeKOP0XbVlAdBpGHZ0GeENT3knc4Jx
WwYEAh/kF5MSzFnWVtLHJLzMY212KVqGD1Z+OYCSprlyBp80uyRIdWW3RDcbGTZ3
2CxLtNX3lOzkl28TUkp9+pOdate+FUrW3Npf3j3DEoI3jwtni5n/c6n38SJl1gbQ
2fQ8saOASPXO3sEltf9ue/WCpjPS4X8FAcDDPMpYvju5BZAyeQ5ECpwBEC57MQk/
11Ne54Gc+GMow5PbMqcqMNX4CMlvlaVC8gVr8tKjho378S8eHS/Py28YaCsQszeP
Q3p8sfuxcF4pSZFfNBuRcDaO7Oy40EGVzrpyuZwy7KMqLbqWYQocQ8Q0+QJ447zM
3eNJCySOiikJmlftH+sukxifxAEKldUyPNltYvRv0TnhWxfgYH7J2injFW0AZKna
KQ2Nr3lFnzC2ENHSQUdwZeOT3nkEUSQ0qWMMtmusafmBCFgYGhlo0aW+n0PCKvL3
nT179tJKcrwSGpLXx61YVlUq2pCkn/ZZ319O21KeCsPsy/4WjfYO2FjgrP4ol/0e
aTepL9lyFDoY7p0pI5o6dBBU/lbjIziMm7q2SYz4hlIWdANlwJ+IXJdzTwyF83OI
Hhk+xVxpO0nbldacvZKYCwY32A4897/0o857V8zUKGvgmxQZWAimLXJWnzMThGKs
FxVv6QjbJ8ga4E0eyGPHpSLhm0SebrZTZH2HUXq/yjBZHeOjc009iYw93joDpw2c
h2jPizihDEqWoaJuYBWzCHbf/XoAR5bFUYcYVvghTPp8DlIK5HoOPqk0El4Ow4wv
09Nm+TJSI1E4DH4bs+Scdh2okWIGAvz3GeiM+2H36YoltXitPygV6Zzr2rcyK4VM
0Zj+R/BlUtIrD334lnMm+Cna5ihOB2/RGKiMZD++EPA1zGGXgvgZUmU91RrtpDn5
Vh47/dfPiywHbh10qBmrdkApQs4DkO2IwB9bZUwtsQrJsC1vP28KrvbX0V2c5KkA
k5IMcrejW2f0OI1qz2pjigZBrfWQKVMM7nyQhVazqxoCJUUi5wtusyfoX0LfdkFQ
HmHxMoiLLHC/PmVbRMXnmsUOKhSVflnUP9EMUzTudFDECCk+naC7/R47VBoqgE0r
ixGwpHpvfwfOWTsn1IXfk6Lgx016r1RuIj9kCMRZvGa4yD76bajgLTZz4Tu4L77S
dgOgYnhG0Cpq2YXhPMqWPWRKmugHmNVE7G+xzlyT97rK3lQJY6auqthjaNpvhHVU
vTnGcy9yugUSBQ2mdq9M8rKkcPhlVyQfXqaGgRUsUsVgAD4kIjABODwaIf05KoyK
gZs4HOxbMeabQb9paelNfAzw8mY/yJeceKdyVP5wzewNxrInMyWT0AcUmP5AqQQk
r1yYw0iZfR+kXj1cbl2MFnkyaFr2qvNbiWuvZI1q7/UsJRYAc57st6i8UHf2D2PB
Ap5/WLrQ2kvYo7z1WPktuxFC+Xr/qKmXWE5aq/nZslmC3O2D75V4N6Cdj1bRp4Dt
lnjdAIrBPx+7l6uusEpTLY9E3oAyIokuSwPVALaqbe22LU01MsJzn864dSW75Cjp
5zXW/DEsfd62hBpYeDXRBK6WpX1Gq7M+rSVHUDAwlU+yTP23QMgTMuQeHQtp5gLn
m7yKl0Ji9IBNkXjxjd8/tJrahbYfhDGzNkh4GJZcNF0c15nkBeNUcdOHE3bbKTCe
qzgJkZGYWVd44ZdGuJ4/RYEQIKMne6HWBBOiUr2YD6ZwOfrszdcgKNH7ChqzyqZY
hcoNRpe0z9y4XaIW8+qQQerGgUjrTs7ZGgmJS2fXY8EGG1X34fOMBR8/i2nJVQyf
6/QcuS+bGs70rQyjQVR0XGVVHI0d6lCmrRkLKcMQHUoaCPIfBhDivPAPb8LeIX8D
HhJ3+in+PoRNzRFYF699sjFU0WvFyCKNJksAzPLEWIJ41j9OPexmHbCL8iV5GHeu
zfwZwRsYsLQSBPNkstmWkXgN4gA8jASJaYIi7vabdrZI10PaheloMM3kVVoZKcFL
acgpxbxy2IXMzlo7oXaQbupAaJQYBxGDx0JXHDsZOSLkmXrymFLBjBooCU7oz7q5
W996oaO2Mz3kihpvsJBQ/eWFRkUT+X5GLvtyU29041iQqE7l4H1/Yh7Nri06IsBB
5A0XfhFdRQZtKixihgzOYRyFkGa844KiCgm54x/UsX+x7gNTfqJnkxiAxxNfYxhh
xy6wKW68ENJwDPvcjSqZXqXF203vV2vX79HLxmCHTpV0VOJ8TXrUcyvXrvP9dbFv
f5WFCw46A9azg0HvnNSZ/WbQuhPajV8uQVh2JOpEDOysZzN+kdLSPsZeq4d7+15y
uPcvTjSTn2ehmuYEFeKg8RiOmO1vATvk2FGW+rAtlvgaMyG4/bcCy6FCslr4+GVY
RDa757l0ThKlb6QCHZ/cW3KSg2/5+aaQ/xV4YCf36ikluII6NpIGwLL7AKZlBKaw
zaX0TmIADmAwIaLASHQCVMiEQE4ViH6m2VkycQUwDWXFoVZLVOPfbd1czpC/54Z6
NFpIpXiptGdg/tljGOh/phTgnVm+ZGzU6B3BPaqzvQn/Pqhg5MXjLn3Q6E+JEWIh
XXYerSx9PHYf+HanlT5E4QuqJ2d/dU5WWnMwQCvBCMIcl9Az4qG4BdyFfhb5d1Ud
QQADmDv8Qjh4b2K9b5V9usCEaRtUdmNT2E+rGIE8+wmwDCtQQc2qBTOqAjFv4hOq
1bWTjHFHr622E0DPD/7rUJ0FTHArO0vfs7Gek71EPjWGxfbnyyVPVrOZEO2o/ygl
8/OcktHaSYHHOOuVYHek+EORyNMBJPUgOl8SDqoki9/fCpU/wmQZNL6v8pkFRSor
LQ6hgjYgVeAJhVc+b5ELYagTYKaTrITEee0FrOhyd0kXZk1eZZRn/MgikgXmZgnS
iz2yabOYJY4gxvrpobQSHUUqAdSpsbgi5VF2+exfrINVP40nGOOv04q+svqIhSEE
d+oehOLW9TiYbbYt0Scab03+0AYv6kUtUlrq2bkpMLBWdSe3SyXWWlLQWbopTr2M
ihujy67pEr2Ywdgqlq9Ee9F4MOyPzehBRoall6IMZrdztHccJ7u7rYj0fuxoQgid
V4XBlGQEXSAgbMfVgnh7pv1P+0QUzoGXZbT1xhoRoRcrQBgdqigTxsMWeMuD+A3Z
EQrtNVA7sWiSPOF0L2fBeF8nefd3Qtt4QnFwBn0uChx5VSCgErIjGWhlOKF+3hWA
vSRgQCdQ9JSHyRAGl70zWddO6qoItUl/jwVHf/9DzJShniXi/RHdODhAMhtsl9IP
qSR2pVEeT7YHMiIpSf1whMhbJNO/UEBOXjolXHHhAoLtEhcu4aVje6dkWwwzrj9M
sormiAo36rbq5/skrdmudRy/BagPqRb6OyvjZ6nVG9ZpwhskkZMqH0OIkGA2wDBc
PLWjyfA9YXfsFzjoQW6qu/XpVuvj+ad5RtSHvcr/eeimUR1dxAi06iFQH+h5/Ty6
EKqf/9LJfdhl8Ln71kVhthSIhblQEvs0I1p8oD4zl6WBtFGUDolooM53iQ6BODrk
177d0lJhoDlFz3WddMtdPq3WtKg1jrWWKGI8n4pxDQeYCejEEi4AFqyAcYyMJrSu
ISG0xBSnlJRkESOhXbPaoH9h8wAkKsi7AKoXjCdaJdIATqRcCbPSNVLMLYqWsqQv
tU2wubzuiUQMxFx+2u6uKdTbvZ9RoHO/9yJ2IXEJqHVTiMbpD5lECAWnj+xwbyY7
5mXpytsBkri87cv6yUKE8hHm96e15a/rP+SogbPARFLeWcvgAlno0sgQH2WnVI/W
NOJcFZn8qKqgJa3Mt3gBMQzFnQFqg6llTN+bdJROmKACFruuKmYfJId+Zalsrs5V
Wn4MiW7IujESBu81mbwFlmNSbHB7rdrPkIg45lzz6iifj2B9ODpqdyysDgbFcKmL
fK4wneuzvm1wTbWLa9PlvnntIfzQ2eRbzMshW6DEQSPAExy0MkGLPg8V1uSb0bQc
7H55wCGiLTT8YPEj+VZLXqS07S906b6pTQ1WsszmZTvEE0bkCIBJbqL3AdPzddkq
G6FpZU1BQx+wib3XIFIFVB0x8t/xOydGYi3XUhj06Sd2JIjTDUtxsqZ9+vp2la7S
ndnqDPR4lF01MTC3e9fkd6aYMoC2526HuPXUNJp8lmslWux4Xesm/fRr00tDgTfe
6zWjgpmuMGbBlwjSa04JyvQodWKiUHLywjkDbqGLQVl17nknNkKX9rp+lELMNyWM
hQecFwcDoyFzgR2Z1sFhqLoFQxndduIoqnGM8OQyeo8Do+OxIfpgGBbPEuMfgPXk
Sz0UFSXQVtZOJWJPXvacuYPKG7MKjk8+HHH8DQmpLgogg6/MGugzXeXflaojxT9E
BDYPf2wMg+kql6Rcfas/vwPQ0WElvldESSVVipOnEv/LqME8jg5H4SVGRDI8hKTR
WSJEc3qLR2FbfrNdDyhi7WYQothr3rKUBxd+t32vZvbPwJfjb6pVMC+I1R0fCVzw
Tr/LtbntVBaorr382E8UEHtwXC627SX/cnATyAoygv22Rf+qHzRlVbB5E0SM4prz
6D3wLqEyjRAr6mb6yN4idhMN1HPfQz4TQ+uUBUpgBwvSpWtswk9Se8NWCSM0vTeK
oIosg771yShFA1hgiq1CKImTOv3XdsH2bJYTaYdB0ZtxmprhACV7WI13SS8Jeg2+
BgJIiRJSFFkTz77wlt9KwQkidOeJw42tbu9e3NBs01AA48qu91ctBvZ7NUsyO4Vz
2uVTyO81gMB+HA0ztQrAZVyLwaXJWagrBsJwCBj7pKqtj8Xr1DKWux0eapTBA/fH
hpEmbZ4hA2hzN8e/U5AS4IHrsaI83j88TyWhkk/1ZZp/RaBiENBKCKlYINyeWKdW
AK2DD+xfLIQCdWxGIpaeu8ZhM7WskIai5rexFeEW7Wc1SW/i3R/ciS6NJq20KeDL
c4oMd26yJ8NXqA3xHKsXqYIfbmbUGmNrEcSib/CR7qnQZpIyaecSs71nR0WRG2Ia
dRFyQ2dPeQbpaoiDQtooqUA0W77zZUGSLKlZfD38+L8OLvmJIYpafZ8mYTRWrs9V
phm801XQZ7tfNwiqn7fANkkPj6f3UATKMjBf0FNd8OHdbaF17lvQVjByPixZ9kG4
WNMkgFv0gOHa2by71qgvrtUbR2qOPylcLF7CT0Tut2VZ8AKf8YbIeJoSaQ5JH4WH
sTHQpf6GyYvUlPvZVq4WmNxISwNeDQHTWpE2HDlkkquZBrCXo1T8uNIfd26bDaUZ
cPjHGf0EHOAx8lzsn8PSsIWppXV3JcWhQSXm+XxPNevFCG5Yzx0zPCQ7twUHRAMc
2D2+LPrBD3Xzzsxl7O7HjqlEXLUrtPw6HP/ZUU8pBulhMDPLMele/lnVJRSewGWv
5r1Vs1Y7SeTvnxFtZBru4S1Mfj3DVoFK3zo2g7SY7eoFqAo+QYvFo/r5/gj+Mix/
Xd45mnB//M5mT7WrTuUjQhm89KbkcBc/nFPKnaVxGAAT3/7T5+/ggvOpgjeldXEw
q3X1koLh6P6YSj3aqY6aYR4cY/sGRFxDQBm7rQUaI2qW0hod6GG9IR471J0fPd3l
lrCgZgX3jYQDpGrgflPIFNbiiUtRVBPwLE8QmS/y9RTaqFsef/yGNkTd6ZF+uEhL
bDfn5ol/GJUHcvE2VPl+4PmEg+tkC/KJAAlSWiMMiM4uuOo7ZsICouIj49FqrvJL
RCTiGHbTXzBuSgaCxoalc5NJyrjPfjpEEMFtucqId3hP8UEYTHoFPqs7FikA3v/r
4Kh7t7yZLYKwl9dsUlqsBQbL2S22Z7gpjq64y3NigjbDNkZm3wz1toEC3Le7dHte
KU2NH6JvAiDY4YYji3kFoMdvnnmRwMH8/7pKXKN35w/CmUvHmPTwro28sOQQ881P
6nYDxBAJuadDTol7R3X9z5OVmWap4WKaEuG90hOr9IrmJy55kbBukCy815HHFOhm
I4JiJjRl2ojB3puQ05TDSlEGP/+gcZSvwk02kS+wTfmciN5QaWDaTT/xmSn+wcDt
SqnPv/4LlsWQiSGN4OPpvAOgRLfU88JMTWf9nK6UVjBHSfSyvPAsrNA5dFVSDp6O
hkxz3BNpPWiIGwdL9+gQF5zlxagIj8SmzA72b9cBLQUXsPGswMkEIxXk7qJGj2up
+DV5ieuKsNe0JkXJDkqm6SLAr/ovKlgMrCFXPw18QCpgYUk0+pcBdS2OnL3X6SnO
XS2Z8N05MKLHU0roaOTcVwgkrJ6GU41zfrAj7L2PHWZoUQbiC3ubbypEJIrPKlwU
FSrJlbk8zBEivP2N6KcoicB48OH1IKXry9b4ajVY89PhER1db3d/hFLPQTdpJf+S
IHA/+gO3t1ph627fEEpKJP4Xe3BjYKBSISgexLPIEw8b7jPYGblt1kQuAIi20zWO
lKZx9/MM4PC81trCZ3rOwk2vjUkXFKigwkIaFw0DeMUiHPpqnpYGDOTkIdRsXNOI
W/Xy++2419i49j43SVM7ODMRBCh376s08WmQKi0Le3fRqP/uTOO+didfTOAHrSFw
zHwRFgMh+6F3Th7cvxOhNp+vTxX2SxOp34jWA0nhpAQU1ctZNkYQUvrdDdhTWTwN
Dm7PmXmsNuBGiBXrp35ETNza8Jw8lasv6HpinEQ+rvKeh3gFqxUSoawN8ShlklHi
iOewIaBjyuY0xO36qjvGjPh908tvwoHSptnao8IVkV5EJyHAra/5wHEjzIHpFIAj
Xu69lJE5cdlNaHq72DIdidexIMeqKA66hlI8qygV2mbX1JUEVBatb9lrzbmWfvBn
yb3MhuLCaoDlYsCFtajzCRSxUG6jhHK/Cgc5b6CPOVerGU3gZhL8R6/rhM+vIt1+
aAHj5SHkrhT5wuFnVhxYbDjVUjAuQ5ca7i9KoUWkf4vaUNnIf5JEyVaRV79AXcD8
h7tL1+jPFkK0B10Ja9ymXde954rJxQ/Mxq+d6K0qmOUtGDuK/LLnNTvb3encfvfn
0y6WW0CS/rS+61fYf9DOGK+LxwjLuvob8kwGJeMiA7sRUDpLJt2ovfRK2Ykz6N8Q
uMCi813rg0P3ZcZyjOqFara+IaHziw8gZ9/POgLx2eNGx0lWtcfvxjDx0kqfXY4K
vk3ZR13Tpx/FCFCEPHBFs5+VEDFIp9fqVgBPXnSJiHsreH3wmPv+2Rr23e1pqzDg
uXMzNb+R6U32x5ZSukJpg2ewtG1P4CYIwuDY2u0BUt4maT+paRGGct23ALZQXSps
7kTadq+VI45bsStCcYHM7ipjDdy6QnqvSYyApjIwlggAGlX5HeIu0yhsuK/LTJvW
Zj/3tsoaJbgObLyEpceBSclI6VRUacQTQsitel/VNTMgQjXoxvkAhvpVvFStekeH
9oV3fCbsNvqURjyHr4/gB4lt2WtjbWzve15a3+/BvE55MabF59FPiLSZisiORXVt
xZjP6P27oLSFA7upFhdpQiM8QT9HTqR4sktvsQKDfE1Ru1dbchwu3gyaaCfB5o7a
Kkle1G7+nxxgSevJ2IpYlnHKYQIBCrTIwBUcQR84OHYDEEDQHQASSUi+v6oZHIGk
BG7Vyp/hUv2Xne/GWzPtItHVWBwxVbUMUFjkUa1NeggkYAKXnfIe67sriDz3ao+e
9x7DaCHWLgI7X01LuaTT1VuqdLGU6z9YLg5eI6fBX6TpmngJbB0vfkSsmGCfCRQv
+4jP3UN6qMSFroeAlgKHHFqZlU5iw9hUJRIA6c1JE1NfMcCWPW0dSuMG+94lh7sk
D2Hf1Y/Wy0sWmnBH997qoBwAURM9Q0moHhp9ouS1F/N8r6vBuzQqfYp9EJ+gVpXA
fisWeDpHSOGp2clmeNhCle3L1fLCZLJ6+Isz8eo14sgTGhZbqftlkcGFfZsWorRX
ekF0QXOu8M8uwioOWrZhNxBMTGN1kMygEIDgxQFTl2UFlq1AKSzPLTceWQmVbKjB
3b9io7o4OYu+7rRw97xgRHsuHyL8jUtkNZ0ZX0dTbOJXQgq9LwFlOPzPWrshpNBn
JOKnQvb1iC+n5nCCJiQKw+oz/PR6Lu1FHvaeagHr5+mb3YZxfX38bkTSE4N9xou6
VlZawrlZQhzJ+/mRF8IcZXRMoizFBEaQu0dBxFRIYIQPKogspp783iiEaoYIiGNN
JLV14zFHvnPonIYuBcwZY9xKKGRNCmLAzL8iEzY6MqckPY7+Zuiklj9N7Bna+dB0
PJf5NXm396QWfzaX6h2uC6u37LZTxpAyyQdSJqlFtS2J8PKDETg2LU4FHJLB//Kn
vzpKPPrj3mrE6Ip/tpgUN8iWpL/VCLZofbs+TZ5PEWovJsaG005FBY2EC8v9q5PS
i8bdGcgQasJj7SCfhiuM2XhKjsU6HjeTWTFiY4acU2OlsbSDqY/S36fIPPmlwNlM
wKX8eCjYGfvyJ000S1YGaiuqJcZnYkr5yyV8guj2ebm6IXBEeroVbKGD8JmpxqGQ
7ldtKNdKaaWps5Bao1XBdfLofV1FHqZzYRATyDXPUgzVhhWs3cFQWyMC9INvcLaB
0y2AMNQWKkkZ6u6rxl19tO0l3HxwKNqmUI9oO/Rk8kaOoLO5LIifnnw5Q2jDfu7m
3s5w9ZPzBgqQ/btiE2+ZbbmObcJaJekR1m3t6lVQ7pBh7b1wBi/9wRMfmq22WmoG
o+4p2TP/QU5kLn2iNBV6ttsAg5vTfBIl5jAcJixTkneHefNIzmszKfL3peNId300
MKKceoAaJqFH9cbVkxDzLQ7X6lkAn6tMJWhhyb9DdQE0G6hQy3qwaxydG5xra8hN
L0RXNCDYkB5txfH7lbVin+A9RV3xK/Jn9cdz/rrNKZ73fSc+M4Eye/FSdsodk+kc
MYYBx2zbAzmzGdogBzgtH0dMJMGPBtixxB+U0vw0mFRsKkKNGBCWTeFdMMBy5Lih
W4ihTgeMtIgVdM1WwGGv4sjVNOKBfQqbJmoQq0mNRaMnyDSV5gif/b7oeGlOSEEJ
krDL1EK+iE0R56dPunHHU0Lr4WxT/oD1C45QLVTyvWQynJlYqG/eUIUo72E8YOH9
1mqJGqfQEmmStQ1BtSiNm7Q8aXZNzgLxw6Ls0Mr9sNjSZVGht5iFGBwwZi+zoliu
nyZfjR4+Kpx0BOPVLVwJCe0bgCIaEr+SCGzUiCw7s2R5bC4IJ9gC958sC4b+ABFL
c/8Bkv2TEfMAPjNuKbzU2VYH3MsfvYo5VmyOHT0EyVBO2gNAuF0i754E3mhRKcfM
YyevrxkNOQKI4q+LA6vjFy/SP8yNEjIoR2NRqtE8KXLoIgQ8GUsPpzz3azUgUspz
EAfPaUQ39sY+wxCkzDZtS9aqqe6jHk9lLBnPu4Sy3r96sUka7DmSaOhe7n10Bfeu
vU9rTB0OjiVKkK08srYDnUe8LcUegKZ3a+cqpMGjQz1kLsznkhpxwteBhAyOhowP
Qa+Di5rafl5jkCWuxghK/mt0M8bUpL9vC+9v9by6GjRAuDIlYEVfcXRdBSYZbC0z
PzUm8PVhpiJ06nLF9+nBFeu4p3K5w8Oel0phZNIuLgKfhc/RfnQ8IOG0r3WcZvlD
IzpQOrGRun1fEsWKoFTotqVRLEytAPzXnMUjQtGIrsJuq8lw7NHCuJlGr0RECkBX
bpEjW80+Zzw4Ux/3cK4IOi3dkWQMoDyJdjGSAyXIDMqINYCmkrX5TbZrujdfKKcJ
uuRd75x9lNxuxqPATD2/VaClf77HRZfhdAFSqQyjnUBzyRv/oOrbuxdCN0v5evkt
yRBKd7dXp145DzaJ21o0M+JI/93HMh6bQX44VCdhgaqfJ4slyYxma0MuCsmB7jEy
Ncy6hAzP/LkqsoFX/oNA+lFMGT5fB+ACtJCT+rZywpIsokXDjjo/Hp/KhA4hcxgc
XuHGHHZDMrgPTA+TSDxRKYHAXTxGaAYgr7LXbzwsHrRTQo8OcEbgGlQ+s9HxIOYl
b23ha4D5aXll/pkX3s0NnowLD3pHS05NtIUylvkiR3HCHIE8fPROlk/mlhZJk8LJ
wnfB6kwJuV/ZWJde9JP84oN/OShT1kMZZ6+c2IgO0uQ0kTd/GRHgkYuNRqnZiO0B
wFUYKycjtVTmF1CRTEMmFqMa6rV2lkScjkV7tmiTNwFuH7jqDJNOe+4Gz1ehlKwQ
TsU7PXxAZiieskrObvxo2qTK4QGsSJsuhWQzxIc039gf9g/F4X++Mtic/cKuHUzf
PuwoMGs4J2dzBZOhYaQuRYx03jUP9pXIFTIcuQecupDT+Dvr2yy682cLZEGHmA3H
MfjJlk2FNKk+BOi2/wjaZJRdclOgb2lil27VfQsDTezdPrIZN5Ccq3f44SoN75ne
id4Fn4b00CsGmdVGr2QUQWeavIl5/cDGfyxe4ugfIGAi70euEKBnCO4/CNj4U7/i
S5pX+aiHf8mUdPZVSZIPxcXCQG+msjeKq1CWoz3OyWA/kossB6o2hWuH2X3mfoyL
230i4jTiY4mlIh+3cCFV6WVKtLgI0BD7qL8Cb3SGdLOEz1LGI34TK3nNfEaRuPd1
hQjK9GahxP4fAZAUrEDyFrJ45l6jHwQU+g0VhcCwTI69GkIZbKd2NBWyMTqRO1xH
28UKzVzA0wywHvJBaq1BD8QnfAxxHyDt7ycbt/A0abYNl8FTiCEEJMfsJEtTqc1g
onHsFsf35mQk4OYm71wXhpiuYL/uCa1zpL9f5T3HwlFl7ODKN8wQbDyBPDF/Dxsk
AQmds/5cdefYv3IeR6X8B8G/BU3NSSWUG1/gtNQNBkh3ITiQcESu8ssDP/ramQbW
4PvVrjaEym6EyxVyMdLCzTn4pgGJrN8M3OCTIf60jM32dChLsBRWFEAG5PQTOpQq
lDVDNvsJEhrmcFfz9xNsJvPeIsDjpuBFNsNKOO3PCYClxE5KWYImcH9mvjITusKW
HG+hNNq8A3yw/EOaG7P30A7+CoHzp/ZkYTuNEP7lnwBHrXMBv8eRorot7dbdWC0Z
r2G0adpTTZbQjEHCUq0q+WnxmPQtHAM8Kv6AxRwFms1CTW2mcuylU1TANZ5rwnZX
VxXl/4x1avIfIkmFqJyc5WhFZBIk8MQ94yJ+MN8/NQ2n+PcSY0LqD2A1tVotOUhz
356FxSXBi95APj6jxsv9fHvjRUFksUNseQRw194s6B/ZCN2ujGoWdXIsg8h80H3v
9DLsed8uuoAlEfGRHVaSGOfuiv+6WUrIyU6iQXuGPMtmjpHgbT250fMzFGjfR3U4
Kz8s0pXR85LM/6UzNU3uUBKGXBMdm4rbQYZvvocBRbWq8s9GR5codnYrpLSIrF5R
mEyNT7WPQ6T+eymHQBIhvpuZw25NhuRheCUX7Tz3DEJBiG78Qr5Z54mQUQgtS5iI
W8zdoMA+ly/uTJcGOZH+BGDIi/qH5zggPgC+JVnWdqv1zXNK+rnUtmlA7AbJdfKk
AeVrYCcPdqoIJgwaWC1q+gWzk+bSHPDwG+GrV5NyeFlOuU5luyk1XcPBNXplxHYR
3Smaa3/cjtS/vSEx229bp0F9SBQZJFkLQ8+fCtOCsMs8ex89kj+0DhxzJQojBHbY
FoVqoq6Q90QADFBs3e1qOUuQ0l1ncHxaSg1mWPQLWTD44Bh5ZD7/OPC8v6vTNrSu
ih977L3w2xHv0O2sOxS3FqAAD0NQQ4ZTGAvbDeA8vu0zfXJm/VdrTHYFDAogB3QW
P423JtzczKxmUmtocuFjjYuUf3gasLjhvGYDCow5K9kn5Ca1nKYv7aaDz7r/b05S
heoEiWmd8gBvWGTtXVSl3V/flFjwxES+VtLNScdJ54MhACdWanou62jSb0VyQCEl
viQPdvJLR3NnkIBZOxchNBVQKo4WIR9250aaku8so5wxDTHy6Wly0VBk48YByRd2
xESNWVN7Q0psNt0qtqZq0CiA1tL0uZeMEdxFjrdK5CauXqiXS9Y8zLYsybqm91MP
2sh0lEaALFssg6z9TU/KbRJ5Xm0N9TMomh1kEak+Xisz5uG0D9ptx1uxUG0dvBlp
vxJHRFwFF04uz24Ag6SRYrcViVWSZgolYlvxs+tuCbOAelFn/5MuTqh9c8rYohyJ
4ke1hAcLYqFQNW/Z5UxGuCOOuWTjm/35YgHx0AXXYlG3/zaVbZwJlRUtEcL2Ptte
GtFkR3jpKpFWzDqa/XRaQgEILRAGVrBZSnQQ47oTqfkDMxN81H2LtaCY0fX5fd/+
fmRueJ9vPl/QM/tuu477GmACVJgjb1ZFKMfh/tGDcwgbo1Qyb4+8HqZQ0NOuE0ec
Zb4HHeqkTydZsWw1emKVaUQ94hLchDSY/yQJTYKRb1D9jH5d6kGs0pUh2gyHnTgV
rxr5UQnmorHmkTNnosfbf6M0v8hXaVU0TmS6K6KG4FqaEZaEH+UDwz9KidZlu8Yf
PhK77p1PInnLDwOJNoFUe54KvJ2DfpPXot4uH6MQDH3FKhtASbBx9XHUv7FQlWmr
SWLmhGIWeNqA1wRyxUazaX2FQ2LlE7/cbLOJaZltFxqYEvh0WfYqfEyCOiVYPHwf
nTexppnVyTGdq/pvrxWCjG9i31qCLi65nj/3eNISUyRdv8i3lf+klT8k/jvMK+wy
xRbcgIkA26YYyYbxpL0kTHd/8VFtq3eENdsG3nSwphKOwal450FbUB11bn4coNup
YXSB0uucj4S8D7s0+nZeP1eMDLwl2GmP5tLr3kGOhvQ6rTrVumBudC4uVwnjaBry
sCyuRk20fc53nDZtFp+/4fk7KMIYMmtPW63y9ZHCw62e5qGRz5yh7FGpPBYWHk4h
tdEcvbpjEeIBFP2y2946NlR0m2lmrH4VKBYmI+PtlogwH7OqadSBW5DJvrQgBJV8
2WK7VfQu5rMxlI5uEia4jGxIOpyrkR4iZDTDreoUf4P83K815mZBfWFwOrvaZ9+U
NnCyILmP91PVGBVSKoRc/Lu3Iz1rZKZ2eiu64I+W5N09M3x+PtE42VZx+2e//p+A
+slvxSyLcuFwjK7XgvfPnQYIoQhUHl+bzVrnCnLTdPlDdSowlusjAW/3Px4o/ZXS
e86l1+qyrpntz6nn+bPU0TATK5XUmT/h88oqwqF6ek2Djh422mM4XTKDEn7ekmUM
tzB+5wuJm+THOoQw5WQuWS069BSgOV2XoXJKRW4jQLTLaC89bsrbgDBvnnBVHBxX
0PXcmk3lLYFB3lywdrtbRqyRAISODPscL3EZCJ6j78USUnAdZh67fmPcDkNQjMRw
2ojG+lqO9I6Gq+EIvdd3atgdvWR1FCCtT3hhMx4ET/6xU2fyijHl1OGpsL2BI3QD
Iy5CSkJ4PXfGps4uKpu+M3osSlCtwnRkP9lWJJvtlw+EIBrjTWv6FEM0gZXe+6Sd
HrdLnUZRWr0GZXw5kIDvv3e4jE7vWikYO4OyNw6cNntjrTf2IIHCp8YQEWxzDEoM
um1Ntjl3SMK5fts52CUZrX7Oftz8Cuunt9yw1TKr4A4P2xO/JVAI+JDEIfh6ABs3
BviiTujEjXrCAHMu8h57wiamDH30Fxd7CZkfV2CNt17kzByfJ3DLS8n0b5Ji0HQ6
cChMKSUuFQ//Q0tHQorTx8h0WjxcxwzZg0w3Gv/g212vX4wSMPrH0jm2z3x35OMz
dUuyT3VbHx29cPq02WDOYk8Xof4KV4NoQSqeclk0rH0f3V6sUB1UDBVrHaJMz5dU
PY9tbkvgOTBJSVo6xNoNYsXEzZlvPbBtadY4E5r0GHKg8CJ+W4gPKsc+9/IqeATb
zOa3HYcOJKu8aFiG5XEE/XVR8IjZAn5+jLAOwWxwrucKW3XINwRTm+Iy+B/IWjfq
K4kWmpi7L87NNd3Jrx8gQgVohlJfD3UNMWg9243d60GbTEjBHDiRG3FfXa7DF6N4
RkFr8JKAAUzDmQMMDL5sXqDRbVa7EunmgKtUpJ4kpHkvRggbBA5l2sk5WlIb28EZ
SlVr2Zm1ldIC3F5JKy2vOJANnlFuf7n/4m0H3u+HPvtAB26JwzrLOEIIjlZLj19/
OFERIvtjuG7uJxJH7uoR19YiKNSgxWvICNfAxXfu3XuYv41Ww07dB5fd19Xhv0Pn
23oeBGX5cmRbkycJOZDn8wSBOkQTlU4zFeyFFlqScN4MVo+bK8yAypeW+F4iL9LM
rwpvuyd6bgPwoB2y0ql45Xh4J+w+ZPP+pdZRlzUFyRMc/DMKJXNdxSkxPkpo/82G
xCrsEWKYg8zPYOMaYOK4NgD50/Y8R+0PKg/Lf7/KkZ3dUDgt2SwMd7zh0B/wBkDa
9z723L5ZHWnsD9B+GPFk6uDC2sBmryKRyTtBH+M5VaUhe50Gv668OPi5ZqI36PBd
Vqbvt29qF4JaUhFnKya0X81KrwnvTDksv6xNVJTzOqnYV+iM7nZWH/BH3V34g0He
6shajpdDhAB2BcofRB/31gBptoJnwyLcCXIRO932OJZsU27NRbfCRW6aFhaZ24Dq
CZLfJ6WtjW+o7sBAZN7moGY/w0h1+0TogdczNgAhVfq4WfUSh75NA5mO6qxpzgqw
MsPpvgcdauPIO/uEdCPUvYHYsmWsbN2psjAyW2hetuAEc6EtxmckaXOIR9g9AYyB
9/wo3wdDXh/nkaqVm+4s/rW6bAsIzFzF633DTrGx3w/1eal3VwrbJKi+JjdBlLUL
v9/U7ULhc/hXOKJv1TJzqOw3YhfnaUlud8WH68fQGAAIVWKP7XBq7vWs3+iD2d3j
lRTDnwihtovpDHFvCvHOe+FYTp1QX3zfcB4/g+EwWqDKLAHTgtf0nZDyDqwxj9sk
3D7xdm5oSWQA8fhxW50GOOWaXcViPj6B2h6CdDk0Ufdg1Xx3gerXjo88RqyS2THt
MXAJsRq3NpEfkXwnJssj8P9/3MNiyUfDYphDFqhGVyixoj4FgfIRGn/+DubUwAAr
JU2G0xD4MhtCwxOpaN9WjCCakfuoq+xJB+p2pTNmFAy7YKi+XKW7m06w2tw79JWZ
VMmwSMlZl1M+Vo8vR0fTduk1h6FpubunqgA9B8oWQprKRoHmyTr954Dj7UNpkQBb
RT++C1l1aczfMWx8/4JPsJsQta5Iq61vzKPitDcUwNRMRt0Ose32XhtUN+I3bQq+
TuvKcS+EKgLS4h+anK1/nH4LB6rF9iKL6sXVJSdBfUGd5NtijfaHqRVObIpjFfvN
EgzyT4dtg9J7Qv1pvZcUzFjVUUcDi2vzM8BHF9WzLi2MrfKXJQnme10lHtYZWDTy
kbPUW76MZf7neoJ3dN1wOGGnImW3UxGdWOPUKP8MDPX7LsEOIBhpBTkzzZ0Utr6J
puKQO148jiXQeLNXykRcRbju9EfIm1L75S761shBDoC9LFVGcCQhDWGVW5AOE5Cd
V5lrP4eSQNM/oclN6VzIJ5CsYZax4nK5Bt4i0XzTOOPb6bCNhfi+7jIXH31f4O7a
sJ99mGzVX5PZuZIw3f7fWVxMt2FgHBjzj0sO7d6tzEAxX1bs2p3398g6pa3V/SB+
Wy02cFQfp1PP9LC0yxRinU1Qn53Po6erg99i/UY88m+b6gW4jLnRIMH2QNWK0dso
hTcaZoggM7qWST+7S4J5rjO5LjzuYshqMkEXcYcQc+DMhGEq6P8nemxQ9iy5YHQY
D31sQrAzAXaz9ORc3zRFqFGST+XvItHajb1VpD3uJGW7htUdg68XbI0+26wliljR
Qy+Pbgoq+nvQCd8syxgkSo/PCI1ZdUjvV8rsIkrtaDbUsgzTcgkjegx3wi3IQscx
HyDDBKJMJJ866ai4Ox7SGEiO09P0k/6GtRfOwXy/zmRhUKQpQrS7I1bSfrsbrCUf
zM0LL3UnwMH3h+ps3/JVSAg3Pqeqk18RUevdPVigJA+rWz2RRY1nbkXvRwWEswIP
h2FIBUHYMb8HQY78SwWE1SwwypbAW0gLffFgQC4fHQfZDwke4408wwyk+ODJrIOT
y3fY1g8BmkaQHxPUvVxdsTQ+6F/Lz+qFFW8hOANZ2QHzdkiXDvJ5yUabpH6GvkUw
XJXpx5mDY8qh5R28A/9sWjF4qEUyAy/L+oQ3x+pphl89ANRDcMtInAWsjhVBi3My
5iwkyLwFoBQSrIjMBGJv4a2VvqwBL7eRvCzQe5v14Lmn10yLEERRRjaz2DW2+zYu
K+bj9PjI8ICIRRmPM0NZHzDMbmS9nbH767+hZx20CzGe6Xr2cdsxf1gi8/kkwWin
q7vzFoUki8l0xP6x5PAb05+Cmw7COHe2gXGpZIrWzwrXLDnOz5oXqNsjoNJUquiB
xg/qRF/Qk8DUX0mw73V2di2U034bw8eVths/zRxExnSQfkMDdmDr6gS/zwiczHNX
p/vps0cyBMyKjnq0iWVRwKkM9vgJAvXrl0bX+18luvHvLRXFQ9Ft5JZnhiTtMwob
Lp/O0fYrw1TiGS0Y/Lok5ruMtGACAo6qRfaHK5khh9c+gIORDgdMsrPHRYTvz6Tm
41Wxe9Tg6RE2ro8ZGtG5Pe1gHSh6x08bkBuUtk71KQ6SDVitPYK/c2v4WViqfYy9
ZFowJxRoxJyfntyPGE/NwKZx6iVkdkAe1yOrtAkVkbhZwZIj7e8C+PYnwjtdJumh
0hJ/JfzsDEphXW7lloTInWAz5+0ZM9w18b9u/mmYCgH7excl2PT1Wr9afsT51zyW
VQcuZX/+DbR6np1RcB+wdzMj0pFIBaEO1+K06+kcZshd7Bt/v9TMduBUbVoObI+f
k47K7qXBdjHLxtktOnR/ncxju9htBDQxHSBXTLs/dzQHDHgmKUi3g39ej2pn0UtK
AwN6rC2orPaIkngb6e3IZOebK+viIEIyikEkOZ3BQpT4cM0/3uAVmJkAtKF/uXZK
sRwGRqkU3YV20+4Fs5twQHOz1u0yKtQxrfQP4AoRg7iUMlVY8dq7/NX51FwyYTLm
WFvbG/BcwpgTepoDfCQ02T3/B+pgUt694gNARKKFNT8+UYFWMluZ7wHH8Z9lbaYs
P26Lik/op6pK6Ufg+nFeOC5L2n/AcpEHvnqeS8UJBpyUGYGSOI8WyPXFjfYIZB5m
IV9Swe/oTfXRpuFWTKKj7uDgeQRk8dSTUFZxsxAvn+q7m04A+3VL73kKuKc16/q6
m8HEbnk2Psc2JxHLtwWcBVMOMopKmehwMOjxv8iguLEpk32FZIcMdbVhtL63a7dA
tw2aBCtQCGVbGzIw6yDdmZHrwVSy0B42ZN6kM6WIiqy7AHpte66xxm+Ioi+lUZB7
pWeM8wl+Hr5RH4qCEKZLDJqwx7a9JbV2v+k/sD1ZXBajXWVDmdp9w+rW4oqbrO9U
5qQZ4LZshaMelnlATZxRke2VU0XV5vsECG6PhDnqpMLiHeEXIA1KG5FAfoL+7K0X
51pCB7j9CYnoUf3bj0/GZ/ABLSE8kjdoiBT1+FKHRphZDP0Mjfm9JdvCIwNeNX/3
22YKimyesvKL4sgIbLLSDJ/SvEo1f+cYlfc/iw4I7wHW4sFNPu6muF93ByyeNoo0
n8010psnfLSwXqbi2jXOB2qWrlcrMzHlJKrIp8DotN/XR0mW6Z5LzEjg08l8jXLm
45EiMNupnd7DXNMqr0ByJ8rQasaLxWVjtYI+peJGDYe0ktAtUYUFt6NWSVru4O7T
aT08sjeWbDIlurdBXH4SPiyvJJuQKihMZIfBEfGRK3/f6IW9h+kPEXMEAJoJlPFS
O5VNGLDRtbHnPnrhFSmWHThYAfDr/8UnvlnfISUjHSJ04ItLhRQ6Fwe/VrfzMwnS
1KilKaghvo6By/k4k5LDmuEStBI1v+KWY62fy49nFv6AhKqS0tdfXsfgL83sgJ9G
wjTVy+Ryf+otCGm42Njvn4Y7UdxBn3+7ukG3E854fMiRqmtQGj1RL8ZSnqGLk9Y1
uYkFXgw5WFfOMnP78DA1/9JHonmbBoreTGJTXIHskX0wiEUidO2thKDtvMdtYBOO
ZlVK++gN+JDfG3BI0RKw9IHcBl3rIlV94nHCW/zGJSJk4J4Zv5WZxYLLTcv3VjpG
rFcQIHOvUwdKpKjuGmYse1mvV7JBpGrPcLHLOKFVXbPrTRNcccLos2Nfd4vNhpn2
Zxm5Tf8zLlW/4R4Pi5MrN+Xf3ylwknWvKjwpF//dSBcbqPvnOwn10uYH6fhoyXvK
WVTHXzAk4bJ4yrABd+X0hGDuX83nrRphlMeBbgFMNOmbYn054eH82Jl9ftkyrzZq
cG+89KUzGX61YGFO1e0YOsEO/Ftr4Qv8WWoD8yafl0eloZL/VwFTyGHSuBlfVCX1
nk57aX0SHKVJunW6cj0nqoN4pNZ0mKj13AlJO12tyG70ZAgawGXiFs9Q5oDrEVB2
0oivFAiEdsqQDktodJVRAYdrE9aNylwHDd2/v4vEPf3i0+3zsoHVor0AtY/nx7FT
FIutgQbmasEwaUgZ4bX5YLNiVsJJrhSPlpZSFC/EzlRO1z4y0jNo+r/QLKnQxoxN
7tleMBSGtE6Q4ofBE6yo9lsk5NmjuMOH3bu8+Fn+mU3u/DwB/UtjmgP/HOWAQ7Ce
2K15TIFLv2CXNEWKZNYbRhlJ0ukAI0ohMuGxSPDF/F1O7E/ECA7jhHqrZLAxSalt
Ln6gJJWM1MKyCk5O0X9NoovcP2ASMf1Gsu61A8a+2q50bcWrat/zKJeCet7mMtVM
sfsID7x8/UCYmfAgdGdV5BAGYR7mOMp6pydjIo9NCHYxabAn7ekK03fcEB1t/x5Y
HJhGji7tTznfZG4YdN8/yD5nZcpaXq21zhqSKL6B5f0EGStRuxtbKsyqt9VWEO7f
DZwRurByrHeielmLpcaq5qUZxMo4LrdUZAviWsxOJGG3TPZgSzV91omLgrh+a5U8
l9epy3lwKSScNwma6VZMaKUNlpA8DIKRSj+tWuUoMIxAQ3rxDO3zwNvcJHQqz/+5
8YdxfdGRVaPSVSkYyHqvPDaZENSrs1syQa7FefqwHw9i94wnCCmTBX3ixKR+84wG
zDlqJiEckQ2QjhsffHgIDJGYO8vpYm/bUtJxgKX7RuZe+s8LuP+DJTap5+6mphz8
qzoSXGXxWGXzx3uNdfwnKQzRsuqMVNMJNinIS0wp0ZNiKvWmep6yI4Tf413Aa5Ea
DBzdRk51K2ql0k/rj44XJ725lBuYKWocj5W+MHR5de7Kh6iCtyWQP98ZeDuDVPbA
QF7B1IGc2Zkn5RMBa4KrQ73NRlNlmA6uQq0tJ0H5E3CTR3Psk2E6CJlgEoHnlAng
C9cM0nN7kA05sYy8txmGKeoz/Jhe/3i/UhjY0MrUuq7bwQHhBcYMoxfLAtGeJg+x
Dryh3N+zc5cMt9t3qJuo+B7heLJMtiHcQq+Z1sIPJFcEgPZpfteRnnWgs9FylxkL
0USR/KkaQ6NYaR1NFIp3M6qfEBY0OfpR1FYbUaeWlyj8oFdeP1uotO2ZK3HeVFmZ
vdPAjJXv3TkeDVPQAxAPEEnbdbbpVIfWfUFZZ/QQrcx/jXTZC6EJZwp1HioN31qy
p1HEV/6i+b6zCmdq82rJjZ3sxGutoU4I7xD7eYfB3ztLT3xiasjmJKUbZ1Kmmj8t
owp94n5ON06ZxX24bLm9ebWYzXkKHdqkUlqrLbOiSJXRoYVTp+sN+Ja1OoLRur4Z
W0dIcWbhUAgzazgQorNr6G4i9t2qbcnAXJ7N33H502DCeMIyR2KIKZdnY2iF/FnJ
e7n4UA6C7TCHH+0AhluD8ddYQJtFwhPmR4VWXQpPvz+2ygZ9ww3k8aWweZ0rrIeA
xb8FMTygj9MxWrsA+lE8fBSFlm9paY877fXTTlJWSacql+peZ9jcLp3ybbQJOZy9
pG14oc+UTgaXoCeVSTtQscxLRabg1Ac+yjBNDR2Y63ntwRyff4MIZoddjczkKISW
gImdKtyhO9DXcKBWlSzacvlbErLI8FSHPp41cBk/usDd25zHc2eyu/pNzWOiW3F7
8rgJfqBQPfOjYD9Xo/m1vUYZhM2hU42YXSg01FUe0CUf0DWpRDGr11pNCfPJIzBi
sQ+MdtS43lrRle1Vr1N/NnNaZy/BWwv4BhAobn1L/QkecPhrrbTEcU0VoZPUbkXV
XcMnO2H/cuQowVYfpvEmxpvaNQODQ3rbyuQvnHu0QiS5V205whv7C+8Mxq749K69
b0CvMlLfo5UbMFwnBafaTFM/3XCTA2H0IoIpOWK4TCv/a5Ub4gRSXLeDNPieRNBY
qBwmrefbAK6pnDo3Lf8KAG6pxvccNEvUqwcE/SbHG6IHOzPVNLj4qGdZAdP+q3fB
xKN2ca1juFeIdcHUOGZVZ6eveqk0+MO+q3jbazljoS+wMDc7unHYe+okFAEPc1vH
Y2WmY+WPhgYvssVwbu+iHjxaaDhYFKDyDja+VxpOvuY0UBddzpKXctADj3vowK/Y
hiDohrt6iJCLfdI32693qlgHU0Hgp2CEd/qOjFtoZyepX8b9x0tXsH4wZ0BNhLbj
2kU/GQpEZZfe1sk49jy63qLpY+nWUSsA69OULzkuduvDormhtVFPU9P78GFZ4pXV
whFWxcxa4z75HwRl9cB6m1/O9fgzHHfiR6oXcLV2bDzESYB6/SDdWUI8aElp2U0+
6hzivvkaWe6tDOn5YXFr3Aa8ONzC7PT6YHGCTrb6EyHOIh0OuwgCstAxiNnrmTmJ
bFGfghtGiO9jdZJjPQ4ikG1SbDQn4mqh6X4pLjUmZMhl/6q+ZjzDjm4ZKFWn+hZb
r3nO+dhf3Vnc+szs92MiZFrZdsGhxv9iTogFqfA+o+sfKWLcut4y2QqavrrcG6rK
0MraQN9Ohdg2WgHOZ0DHGfUp3y2erOaj+NCpTmMQQeuxTPkITe8fLM9J8ep01VPo
r8BTPBcFNBHqVjcyncQm51AueVifMOwHxmUKda4zh+BiR8NsS6H5+7diTYFHyYxH
8rBKDGp4oVa4DEHubUzKqhLcAKIjiF9Zgp5KxfZDMwFZHWP2/aXKqSEE5UBE4nXV
4eTXIyeJKAxLNgRrwT334Oa8yN9rDUvL18CXZ06b3QSlebdXivnzT/ZyV8mi0wA/
2/iT8x1soeILnKNuYKU/H6yFpPK+L1d3FTLaKtGWBI/kwQboHth/MF1Ft0q+Sop8
u42KfrZV1G9YIgG3TSRMvSBjsN6XD2hf6fgP1SQ+Yj4MiVH999fNM6U7LPcW1xmW
l8omIaLj2nfA7VSY37GxDhndSIiYCSgqu27mvinlgBVkTQ7bmRpqHoSRrgi/6l7T
IdrNP+ZMAvkklsY/yz2iGYXonC4DCmDs48UpkOV5DeBN5nQpUWIW/YQAbdTOu31t
izdhYfPZW0GdPOJuF85VebKE08IyMmCsYYUEc5ImJwaoR6vEwXlgbz8SYg6LxyrX
SkmxDw7DHWgocIhsNISVGPLsDxLOn0mP1Ldhwr3RboXgbJAIf9Yc3KHOJUB3l57j
5ytmAquC7deC+cbIpfX7c7rq3uDkG8yDH5BMpGGZLGdXSvl1+DRBLnOmu1sBErd6
mVDKgH/jPpN2RuyfbRWQuyD2iFF9XCNqfT7fsnvNp8QJ0OKrC2uwl6ARGW8XcJtE
6DG+c4M2u3yturozEvTJEdY+alk3ZmDjwcL1ef/I31/+i87IlOmRU/nWDVm3sL9P
wapS6cTE4lNu99WTye+irbFB98ekVBqWR5/1AsJp7WZ3IMp5A+WzEw5KIp1tk0qR
BBBy8PEoCn4LhlM0+eH5wJKSjqqEfIx+uYahT3jrjr472n9v+mRt5KMSa9bQj+hI
I4QCUInSkPFeTHgPleiqYdFo5RKkOk8u2k3P0zCRTq8wu/V1qlRpNfEGC64lWasx
k+3yG4mxanNDY4th/i7ZXY5FnWnrPPV5tKeQz5UskFgZopv0MfXzmCENaCbRXBtm
4ZOg7oqcUbtTtvzZAiGIR3XbQyyojz8s64Uu+mmTxuk+LZ3+HPwASjSSy1DQzWS2
aAWj24WLcN8jpIY4BrEvsGRIJmZFI8yKgdPc6FquOSpFG+zXpr3PPfs/wBkTFmr+
xPtwXUsVgYIHXZ0x4FDvflyxdyhEDGSERq4/uVoTNN0u9+/xL/DKt/+fZYVjn4zt
DQY3uv0g6pDaCHGFyFJgH3PnWDlkhOeIXa+IhM/qcfWxJ5ZLAuQjCVdeArRoTZK5
ynfBk6yrXG0GlZBNo0IyEnkqVqa3mW9XOoCLrbm78zvLf380SUhOilSR1Z30r1YP
Y0SyZwQZUbSN69vcI416aEjKLB1wqSxvBB0tswQKhonKIJUyPkYN3hYhrRBLjEC7
MrHhJESZP4XNWERCDhGNAr/CReNVeE8Td7HXt++lQoiAmRweNB4jn3PdevQkj4el
b0ifDkcbdl+rrvI3AZFRBchY1J/AE9PAwrCMF2Jgf3rqAVpUjFAuG6P5sQ7uH7Ll
Bs3i2KWsFulNe3QTRIrivaV4HCIx1MpY+l7cJ0vql8m5iZz6tBMyzjxjOBNyJ/Uf
A88haJ1kRQXKGGS4OySVPGBEG4DnhwWcSShjojrElY1RX4pQvqTDkwCGHs3fCNXR
hCeSkY3Y4AL8vhg1n1nQFAAmS021SV0jN8QW4Q45+D10vHII3HHKxnjWmg6fQ0z9
NU4cfE+E/T4TXZUJzXeP3pFJ1KvLIBxUcmKNls3xYLrZ4QCKzyDSIQoZS+7060yz
8qp1oKmRo/nGO0B8B0H/Z0SgYMYSc1Ig41bK2jk/+kpFmyQQysk4Ru7/udCaD5Xx
MKAvGZWwmX2r9OoQv/u0QJkdh7ZMy1OY76VvEhze9hhC0nd3D7YCDakQPjFyuiby
G5eyCcmu0vdRnz/PK0De24pLwmUYJ/HSfGlMYPW/gmSsLsD8+2vpdfLKIxhiaqwY
ONsel2NgEjFEuVQSXxjyw7/b7e+wwJeHCquFw1nxV9M/lXcSALYTF9cMNLJUe3uN
oEKEwMMqoIFsrsE72VcdJISv79BuhEvH+oN8puwK/HtoJ3jEHidPiQ64vflRP87Z
to3yGUs+3uM3YQBAA/uKuAkD1mWlpV1/UMels6bS84uY4KQezOCFXo5iX4cRt1Nf
lt+j54BYXd3HXonC1Jq8hTFll9GH+2vbP6rqmzbuBFna3auw6LkUlHXnLmodz+ky
eBmxkQu2wirABv6lMgkpWSgvrj3A16GargHmd8/y3xoKyJsyrVMSE7pCyK8EEAjo
vx0pMxob3+1L24ay1p4QZ5xeuiDb1lztTKVhYvzjHzzenILjtmdYRSMcd8PMkJwS
5ZdKFDXUtf6l9PvkbEOxExh7j5Onwnzfc/o7+oo8A5c9bX0ubNOQ/IgzWMNFqMah
blNBvC3uOwWRbIpo0qWWJndNeTUi1bMqmTzlaNVIEE/HqfoJeEW+Pco33R0TI/7P
3KXzm5QX+1h8IE0fo5jfV0Wxlfuust+YD0tFBDVj1ME8sGNe2ElHxc7BQBPpEBI/
cTjcQ0vW/HhrX9j+WVz6GExLPlfEg0r0rNlrzy8HIMPzuNpEELxeMR1ZpdThTIT5
6DwPcMWZY3c8XbjhsI7Fuh3dPdC33NLpRmIl582bMX6Z5diqyhuo3+lRZayYsJxF
9LEAHBQBeR2kOQ2Mdr9vpqjJ1ol4avGEZbSHBXcO0KHqKHBw+3i8XYqbf9/yN8sq
OsPLMW9lrk6qKy75U5CSMpjzFcPVm85srEPhPBksA4ANQ6SrCnyHkdziyPHZv6Ia
j8tb60GHT02ToKUihQrMQ1Of/J9lWjDYXH+Q0gpJRYYQCSGhtqPujm5PyHzVoG7d
HfsZrXUxuKfXlxegyIJBHbYIb0Dn4RezkwwRvHWjZErtHnkC/BRWdvIK7lDpTIsA
tNhNO8tlglE/dzi53km3TnoMtSfd6ySUNZTJlXdq3pGaY1chGwkNkITEVORNdgSf
I/dUUIwTPj5wZIiUFSTY+L1T3WLhYWXd+lP7+FnN7EzrtyrfnLCkDIrQ+5RMLhND
7WflvnILBpeI+be3b64+kCH9OffWTi5maE2goPC/sJAabOfTuwOCsLvwlBtkA6d/
qEzdG1lMBin+vzQijgn3YLMGi7p7Uy5gscheG+DC9/l7ZACD++17O+oSlVvGkFdZ
unWYt8kok0SPDc0n/gqCXiimGRAFBC1lc6jV9P/Me14xGved9cFyJ5GZ6Ow7aXh8
AcD4WGghHSFs0f96y75LLVPvFrUm3z2yU79pHGwNd45q1jKuXt0nDSvMBmCT/j2r
P1mJe5XLk1+jOR3nho5vlAkOQd1tdsdFIHRPZ6NkB4/cUMh0+hfktRwAKidUyOsR
TIQ4M1asIPHQpEx1oorh27RZQiG11rVhcniBs/VpWMr+ZRmhAF+xuQIkYJUvPuLM
SZznh3U0PUSZ016yS5Rfg15+n8FkAYpr841DbPHzUkCLuHJflQxutuVjIkTKIrFL
Kyqylaa59HtuinqhTEhJYANdrKbLLmidFfzn0cKAcMh61aBiKTBSwtqLyTzry5Zk
0/lNgVrBbmdFgKbzIf1zsur7q+5HQTcGjr4YaEwfB9UgROipXKSMQsJ0+hnHttTW
SA8Bhaq06uuSqcFoQAJonNU/J9jwBA2SjUr3/JFG/uRH+m+zDmPF+zjcAVZZX8jK
OHMsEzg1en3XFlxOxeSpOCyhWPFESYPD7DIKrZBXJ/kGejZunhv9K6k/V9AgDUXt
oEIn7glys0QhFakaRGs8OrKSP0uvRIXaDhEBd8vxoxuXi+Py+UOczxnM5nztovDf
pw38/B43P78KaqNt4FdX1ySFF3nwPo4/KO2ub+xnAhUqMUL9bB0fcJi8ox4t32n+
4DjUkj1sRZeFKFqbU3Fe85ymx4abLma8PFe5a6p7u4+vwizp6u7OEiu8C9WqWMwk
Nxa2Yocu7Jdb7vQWtWOFTdBgHR7GsBNaEluPfRAG8bzK7DO96D8weAsKxAkhGH8l
qDyQc69p8/u1ZQzpj236VZlSfHGF2qGQgkleHRtYd7Do5XRS5zRjze4GyfIB0KOC
A76P3Ol9O/iZvRA5qnsc4txvWwxYedU9dGUN9A+eJOi4tu+h2pdQFWRLZIorQ2XA
NnS5vSxBBUmzGFq9DOWxQZqiALUAabr73iF9YirkcGFcWCCexF+3/uymt06SVtf0
EJevPsWLmq47095SJVwtMhf4S6DeYSZMKKwRyfnLU+v0CUO7jo0q0tB6zgNyFHEZ
v7Jel++T6PZt2aRgw2RjMFbmxcfWrGhVENoTmPW5GJCJc0FKQz5aBSfLgA3Y3P1x
N9WEOuwPhk44wG3/RL+vY6RQTPeg1IB7+6Wxpb2Kq3a3KVh+eayyEapZBFAv9/ax
9oxhE4Pr7WoFpdSv7/wmmU1zG+d9cuWO3BN9fTZjezpCBHDDr9gqogMoN+m9tz+A
XZPSz/YniWg7hrqxJPdhZ+1bqsV24w42wFGV/OZNM0FVfT865cuVC8xOQPCt7DNw
6p5DTA5jd0oEWKziNZ9bpzR7gk9/0vOEP+DQogSWRziyxKn/hPxsT5kU/8nhyH8s
p8aTYEcbneRmKujonwic+XF5pAKHNC/Mj0cD4gqFHlpOhAW9itperuFEploxgtDq
7/lVzRRwZ7XAcnU4+OJYG+hB5LJpWrifptHIMjHEl+cd/30RBKWMcZb7NrXI5dnp
PxXbk2IVUK5bK8+9N1rEd3lY4ADucIyb1GZgHNDnao15u9nbBaLNsdoStA9m8VpU
1HGMR+6SSOAcqrq3zfaJC8QHej+m0XCvqnU8dKAMiA6trV0ojErsGweJaxQW5oAe
gNK638BkQiSF4iEkx7Y2H6LhltJEVrGQcZRnKcJPyFpU3lSisqbtzXmtuhXz7js1
nORsYrwbiVKXVuxIT5iKzWY2WOSGYHuUiHhOU004uoRxU03d2CHrLWr4owxKakW1
/A+6eVu+v9ncezxqS0LVZVunjKN+pok4C5zCLhlnlKMbrXqttyT9sHs+eVPYpSVA
Guow3A+ue0S4FgwlpZWLpwC0ZaqlsU3RuGcZp4OytcOkbg0xevtw8ThnOBC6+6qR
rWZvaVDSiwfvXJZLLNsc5N6dWUNJqacWQFsXQ+Dn2C4ZHd4y2fHrCrOu/9zCiIRb
dgRpaTP3BUiKX9gp4KRBi8er6MZJFFx6ILeViQPLvm6NliBuIcPMT/28G/fTf+ut
sXiPfpKz4ci7Zk1IHz/PL4b74GSC95qrtV8Sc4DlDCJKmh6eGKeM5YK0hM+8mNzb
6GAEKz7ld0UQsZLJ/LizYwA+uszZuvgdbAXFEQRvwwO/7p5A2S1AzfupYA+bY1RW
CDJPZS99gxAIRI69cYb6cBBlRPawitmZ0AWs87P6mCm3GqPWhreC6d6qvZ0QjIB3
CBDwZX9uIFL9Dva+mklmZ+AawEJofd7356ZYGQKe4Vcmlm2lR/JGURX/YphOPjhu
VG8KOTqCLAU+uBBw6C8A8zhMhWfRDNtJAds5lgGFGiCU0UtHEIP8XYA6PH9sWgZ3
ZapDPgGTZZBO+oaApq3ktyfqO0s6mMNDS0ZAzKUmv2s1F0RN2pgxv5YB0VpS/OeO
yoyTPOIuPfFtu1aZ2/jCMtdccxVCRGAe6tcohtT5JAENnw71MvZIW8xwBB0+4fgG
orkpNrAy9F/t6m241RkgIQRY770ecuJXVtFw6TE3w+YsmiG5J771F0AF+jFdxPB1
UcPoRm7UkxIQQHdxeAkW8890d/ZTmAe2VDEjpK4G4aHcNzA26MGV4Btq2ggrhHvF
DnmMXOGjphUUMZhava6GdTTfDfD4CZmzO1TDfibNK0hxtFgIIXu0Be5/2DpvuzwQ
2m8xWxeCOWkGUoBvnmxXi3up+l8hGJYHS0TuPBWXzA3P7pj37Z209tzrkHJjsSpw
lBUokLFDjfOBSrPcfPBqrsVLGVJJCgzsgZ8jWHXafhI/GdY20evL5etY8aEXRpmh
qSayk96som0vhXH7lb9AO2QhyydbFnn8Ey2a7oYF1DKomXYbwlK7pN3lCy3poWxj
fw1lWJaRjszDEOT7GDZy+tcKOxerKYT2KAP2AhBT8n/4+plpi429hC1lPwwUh82d
yz3LjzAxDq/xd/GYYTGJ7rV7qCGmlf4jLxE3MN+50GhDzG1CNQvxW6OgYjx8De7M
EdfLN0b6bhK2OMZhB3eOCs3DzhFN64+VhIav4/zEqJKUzjyaDHBeMzITFfHZwRwq
aM+jUVWQrw1hPs1X5Tqs2cgyQotV1UXQs27j2ngpCMFCt+Fsp/dWbS+uLQXoUpsB
f9V9H3s76zGeixOK+UFjQe8bqAz2rhQuBfS7+nG+FcmJCl1PvXDCO90cFGSp6S/h
IrSJ7N+d+fPo9Qkk+L8iALvAFHzdbgN5XjKSyRO1lEEO5dg76A3EN90Ko2MSowaP
GwtfrrhO9oXao+Tc7rn02uXYkykAc1jVoY+YPEoAw/uYxu0hOYJIkO6vZl1PV0xa
HQS0wLUogogWxTT7f4gWczgUT2kWx52z9aCRL9gzjc/kAPtKpUY9gmX4CsNW5QfD
7Kxk2z8KQ5lMlpqmNIXnbs6yoLzQ8j4ZB7PnrXFaa2kzCa8PnY1iI/LMEM1jAPSY
KbG+8NdwG9Vwvd0SJLGw0Xc4cEyGvIcjB1SvqRRocVXKioxriYyYNen1nm74TDsP
3VHHo1dYEuIEdgCuo47ZQtBF89OXab1GV4YjSRQsmqRrit+X37BFRQ7Y4BEe6Pj+
5dlXj9ZeM+QEBwN1wAB4lAc3w1aV/X4Xzbo9DsVUj6fLUnc5vqEByCOWLS1KHkiQ
nOoLpxVoFpMbi6VF7w2BR7q9R+Fx0VYQKYTQoxs5pP3Nmm4EB3N9jmL8O+x0Fybi
uDKVhLVk6FDkzOrziT0CtiQ9cn9DFWzp4EPgzDC+pZ7+OfyOxJdCjhuQJrugM4It
8NOQt6Cnu7YHCMYCe5zH06uwO2+QNw9kXMRdKwViNkUo6nXDTseyku9if4+X3vVM
+eJmLrg9Bk1H3Arq5EA1ArI3pjyXFasNN+AaWJw09ghJ+bDIWMJopsAQCvrwn5s3
eqmUsUA8z2UsEngwT+x00EfCILgV37dJyGjJZO66OL+b1nXfiusP4fHRIAk8rZGJ
PwT0FFsVe72/+3oRE/PUPVS065qMzcVxVjXsDAOCuLRl/4jsJPZgvDwl6WoHJeXS
+E/qgCdPcyY9bnZHJFMT0gPjtMPLvOXgKBC2hDIt4jf772W/z5YyoP9H0yEUzZ2g
tQn+/tLxweTTIaK27z0ZzGIfvu4gOq6kz+JR/7pon5h1NvTwk4QhX1AxpcNWFJO6
bUcMXPCuAQ076m/uSQSbKVRaEAo0HLC7bV7zFd+YRXFazW82GyN8vT0xQrn1OCoe
wuLxuiRPPOAA2d4z/jtxOgpzjVQ823g4Z0lrcDcmfmMhNfaOnck0CjQMtLjNgkTs
mtVOOVrcDHa5irxXzBZc394+2cXgepPrkUbHGk+S2KI42GLgL8l6nf9ylLlmb8Db
f14yZTum37yfC3+HUMO+D028e88YJR3xfUbpkmNhu8G+WC8NNYMwzwoEu4kuBhdi
jB2hYZWm/eEGBLl6teKi0Lf1vq/wLf4c9yNTEEer6z9i9IGjSMg/hef3r8hkfiTf
LJ8GJx3JXm+bYxl/V8NRkksYPc5UABwvUnV9sTFp4VnWKKOHD4SEpC3g/xbYi6HZ
py4xDEim83Uj4EGC6Ilia6Tz46WKiWo06TjGn3EtIPYn/v49UCiKLdFkyhjsnhjg
GZpykIgY1FM9OwT8BqOc908ru0Xx2MS8/rdES0fo5rjZd+JKwFpgwpM2EQjYSlyE
/3T4uzhqQs30qJWgeC3hqJKLYnZooFTDc3okle/Gn4VffGHZvRsXAQohr/AWM9Uo
EnpU4bQPGtWbgkAR6wZRjHB933dWpFG2QTsMmWrE5aO/hag1OkHd6dSmVGbgutjv
6TnxHFE8H67qLVbBvP+NOvjP1H99tloVYs/RLv22eCpd6y3hpHT8koDS+5PtWZwN
4400Rnf5Shj/cGa0Wj4mbtXFkHruijLL3B9sr90OI2X3JUKUHC2emtNLA6EX/xyB
3Vyz5pTkB7OG6Voyf2iayDL0U0qoA+3VWlGDaCwupyP9dhyVA4bFHL4IDeoYxc4F
2GDiAPNE/6B0o5LnduwOpcYzKSBCsh5jaGcuLCNhsdeM89I7kbSg4VqFjZrvSbPU
fOziObXIfEG6wQsnvOwvjNkJDlXNLu5E2V8ueqOycCAGkQAZuVgARvRU/nXyK5Ye
J7mXBA76BYaK22fnRc01YTtWTG2RdUGcfhTLEfsWZygFpddGNC2UEp0F4Q4UmtUz
dNhjJ5Jc4DnIPHZUJXu8dR7djmMW59t5y5W9HaODg9LvRbcIGm48WQhH++yQmpZs
1I5mvC2vl1NlUnw4IXH1FQzqeiZ6APPG8pX9MgiYLd8MIVxdbEuFguI8x5xafTDt
7DH3F6fbs2hKhMvN0DVwPPM5/V5vxkzuE8YW/9lFhar4p1EOJnM5C7rc7PWYPnyb
l+8k/zuvQxQYgW9nHQ2cndZotK2QPCKCIFGI1qU8LrXaUfsGOu6NhD0i68rs30uf
reGi7py12P0lVAC1cdBPuSQnQGiLtBPHjTZyfG5jJrXppnOyQO91NG2qJ7N2+KDz
N5se4fbcrbdxoofGY+tCQNXK66LgRaUYGAokfPB9cCAVDVsbmDJDi8HaBio2sjb+
DZefMPEeHz1DZ4dBZz3ottLIUZjrKjeviu+nr76uh9/DtdyEKiQGJgvGymRzD8ts
BbcVY07ZqOPcMCVelWIkg6AgjNpH8i4jlmvxzGPfE+Fk9wG352Km4fk6j+th7o6U
7bEMSzsXVGO9D7gU+4DskZgNIMRpwZcgRaDIeIwumurSA79+ipCqfO8oImQMu+BD
sicGz52akxBGp5fBPIWiN8MXRE5EyN4xuRcc+gWbKXlQWleGSuIBNdXrJAPFrRuX
cKH0FpwXLZVoT9FqDJPhoK7GFWIizO6bD5oq4E6Gzstpk5CTm3wjmPEL823zDaYX
43quVF/+62+9+TyGXwGn0uCy3jDCtKCTF3/YgQXWSiJn9BP9el1kh09psJwBvHJg
KTGb5OKd1o6QmXnSZ2lit132/HXgq5aSMltgFjZ5HSVupNIDNVdWNT0Y038AvQN5
HQYm7BvoaQRUoa4VVdWPK5YMIP5UevblHDFHWZO0yNqzpnEWwwHEm6+Am79xaFD/
tJr5LX22uRwragwQ8ffnlDSFMpesPlasgv4HaNzKwOsB/ir5QBiLFyEQOeWs5R6I
QA2Y6pHWsAtp0st+wo1J9vMhoxaKIMyA8LxvIomUcUUPlyV8WUT74wlOSXnho8XZ
REDUTg+7EEqCrE88ygORM5QCWGQwJ7eO0sXAOriX/ziJ91PE0nYwIwL+P8OgGaOo
mu8XKchs/tOi/G53nqpbBmssDzsSG/CrhG/K9Bn9fzw+LCgZZn0Xk4lyCbEfhYSk
5gkGpYqwEk6pVOGkagzklhOX4mU28BOXQiZNTQUWhM7E4mfsuML5tgbcKBz8g9m1
f30LHsQGRpw71Spcy0dJ6ugor7yYZheuUU/9hb11t2USmRkang112+fHWfNQ/cKa
gWCQv6MZncNNe3dJzog/0RNGImYWFel2iVPC7hRxNbTJCbXfzumbNf1Og99L1FQn
Jeo0nCG6cpR9ibEwMvtkJIIojKjbIpqDV8QLXUFb0uxznB11vh9VdCaUksjuE+ux
n1dkOIB9aLVV1tbUcWqHFKLqBo20i9c46vEpxi8u+a+eWGpUOqtOzgHIehBQpfwz
hlh2KQMa3U91yPyBpH7GSJrOwN8ShHbCozCfU+Ck9jd+Milq1dfNXWyGz5Ri/ee1
KPv4tepvNoWDZhpGmZrO4QWYY9U6ZhnlFf9zYBZ9SH+AnHMk/U3yWzcnA6s1jGtC
w3vlyh0QIm01SG3JSqXMeKTqHLK/cZXi1IUNFUkPAxH0ju3ZrJzrNESrvYpcizPY
IdnJo0521RdF2AxvBVjZvfHJbTWFbSHSobOIyEJIWGA1SacJltjgJ5pA8TvvM8qG
BlNbakBOYB3IM9CRSAI7uCsUCXs8mcfWsE9oqgnbSdaRTDPV9WwJgv7iT0+qsBBx
8KYxLrRmhoocC+Bjk3qk+SSV89uDkEPyCScTKYnVdJ3BOZcHblp2CHWaan7tccWQ
kF3UmoxmCXnncZBhjKxVlZNxj/SUPzPwT7QyvNSzJ2Z9l2nzqjkbPsCGOnOcbqj7
FzDSR0uTv4wv1hz5/iNS5bIVPoHGRTvRjgrnw8zI+IMW/rgJdEP0ZiQvZTyEGC5G
fIoAeNbXHWT9MrtAQw3sF7WfRriiiSlmA4ubLtc7gOtKbIyRnj+QHVkn0Bo0fqcZ
ULBKNVbSPj882gjV4MGxeDpAMBRDOsYYY3bWyl+Y0cYsVXt/FaakiiaREo1xiwvM
jNlQ52XXsnEPw5QY/uGMBm2z2vaOah4/REg+xFP7nvX7txRM+y6OijWxObVd/F1V
Of5I2eYIQC3un84vLDNHqrPfi9s+ane0X1X/Fvmwq7vN8ln4EeDMSOIikIBk46ha
+ktu/kmdh8VB2iyI/jtDDG76V9h6MIX6HPxqN97L0XsOT2An4E+OL8HIlSDwZd8M
fiimOc31em7pbZQg74OD40pp9Q3suPjuVww+M1ppZ/cuOPZlBzLStnihLMH6vILy
/IKOJuhzLkirodH02Mk/0SAXkYyJmE1xZeCFl0PaCfFvYkXJlRMeCt2iBevBHwqi
73AciQELbnXvdwhDh0XGx7/XBlfwME3PwsDakhJRgtctLRFlJMPQXEz6rwL+ZXY4
e8/jsJn4i0u7PEivisSd0WGz3HuUG0d4LNmDOPbNDqSGjQVNiHURk1PCqOVjEkgV
UvfPircaH/eQQDZ5dSr9ROOHrS0X1P8GDh9J6wT2r4+aqHXeYQbwG2l40pW0x037
Iz/9c1HpZOoZSogam8IAwgTmS1qbmh3PbuTPKgHOcsTiCzAoa9PT0xmpCnVi7Vy/
boHWSZzOx6n0urFYT8tBjSXiaX7Z3422jtIRGLWE4tFjN99e1wke4aDmiLOw+3S5
tDmmnRoH1pJ3qXx5VB0zUVxBlVwWz6maBEHUDBYydX7zvd9/Z5G6Zul/WrZx4dGp
FaaKBagGEd8BuNds0acL39iNSs0v2qvWxVQi9GDix7iI3ilkF+hasEZ0ggE5ql37
wbF0LnHOoBWmmVS4FEkauotUC2rFArn/hWTbLgbZhon1qUE1rQh3D/5ZQJAaD+o8
rqHWCZxMMXM7KNkMYB2O587Qu4IIe/qkaR/iUEmuyRXFUzKMYjlIPDcXE7/OZx4F
LhzYISK04l3SgO6KI1d8bQE1jy6rM0tJVn506FeCM84PeMvEp0qBWxYfO+7S+6pp
77oS5AyqfzjgKY4iNPUVPw9dRixcbZNQg0Bvltb8SfWXFhH2X32NIOQiUzfn3Gsm
CAJxdk9ocptDeIROiIyA/1Cd3nfrxsIGmaTdZ/cvwIT+dMSQZqcaBrPIpJGThp4u
YSZBMzToAFVIsJhgH3lQGOCb9L/gn/sM8DQ0yftgq3yiE7+5QBu80V2Tjz/2wwbO
sIdy+xUH5ChK7T1AQxTgeTaispTdoB1/n8dR2Sw5HkBQ5LiOVjKsE2G9kI2TAj9A
9wB1Q5DXbvD76brYxFQWCwqJYBGa7jlb4j3mofBQG/uSunFaI1RYK0fTR4yI7xP4
psPYj+i+2mezXVqLcMdRYN98VplodvgV+0y9tr3meqF3n/MWNwzF0GClwyJMk2P7
5L18p+rqrHQkkcmzm5RlwroZVJ8nLI8Aohr301jLWvI01RDH/W5+5FAZLY3T0XJQ
n9haGUDm3uN9ieZ1IemKcsdS7XbYL2IDIUnZknmLe8yZa9RSLbQxJplzwRS2FhP+
SyRuTG8JePfmOF01fXl8mClgCLsV95awSHjqULtHJM8uyuI3GlUPal+p9UHklDQE
pqTMRiMU9R+f+6SZztkIfdfLVmhQ3INmgBjlhtc9Y79WUlaDzFAKSJ7fscKgobjH
zGsBY7Wi6vQuKuMiWWS6kDtK7zLZl1z4ZamFHLf5o5JQzd+b6NCstbWkHPlLhJDB
YAFc4xPpTu8rie6ww4lJBZ9iA335tprktf8jUOPK4xYYDcySREksg4oKLjIanpcS
mhwIg8SGacnxhfLSukoV6axA+C1RwGaeahRS4EPCt6SZzVqb3dDplW6sn7Ae+gw5
GfyoFIhaRgPINnOqcohaTQVLju6CBYbJog0mvQ8+XF5nvnUI1YekBhtHvs6CY0vh
YWd9SsNrMTptEEp7EDNrAyuIyk5hSFjpcQSnIAK8MtFzkJwxd1jHAyTlgFw9CFGJ
O8wYeHDIF1cCUp/ZYZNtA8ovCAiSZsskSdJL0d7w4kBdWXAL7qBdIsXxSq6bxqAs
Y0A4dvKfWrVmIuRg53w29MWsyYMhr16TQwWTldQZ1bZWyu1Ql95ucHl/jNdT4qbU
ZwQMTzBKMKbxWjQu8Sh1QmaqJqhfe7q3R/IRoFWXAtZHI5gFt+XQ3sl/weWhgPdi
kNmIkwqUOySV6WDk3R4cHhQbS3zF6iwEtpfYWJDadbCiEJmtUF6YdZSeocV2bRM4
avJQt8FwFpBHMj3eH/HjJQ==
//pragma protect end_data_block
//pragma protect digest_block
jLuaOHhMriUywHvvccBcRNY6qkQ=
//pragma protect end_digest_block
//pragma protect end_protected
